VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder
  CLASS BLOCK ;
  FOREIGN decoder ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 75.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.460 14.490 26.660 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 100.060 14.490 102.260 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 175.660 14.490 177.860 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 251.260 14.490 253.460 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 326.860 14.490 329.060 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 402.460 14.490 404.660 56.920 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 478.060 14.490 480.260 56.920 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 5.540 33.820 494.140 36.020 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.260 14.900 20.460 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 93.860 14.900 96.060 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 169.460 14.900 171.660 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 245.060 14.900 247.260 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 320.660 14.900 322.860 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 396.260 14.900 398.460 57.330 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 471.860 14.900 474.060 57.330 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT 5.540 27.620 494.140 29.820 ;
    END
  END VPWR
  PIN ena_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 74.600 31.400 75.000 ;
    END
  END ena_i
  PIN input_ni[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 74.600 86.120 75.000 ;
    END
  END input_ni[0]
  PIN input_ni[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 140.440 74.600 140.840 75.000 ;
    END
  END input_ni[1]
  PIN input_ni[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 195.160 74.600 195.560 75.000 ;
    END
  END input_ni[2]
  PIN input_ni[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 249.880 74.600 250.280 75.000 ;
    END
  END input_ni[3]
  PIN input_ni[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 304.600 74.600 305.000 75.000 ;
    END
  END input_ni[4]
  PIN input_ni[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.320 74.600 359.720 75.000 ;
    END
  END input_ni[5]
  PIN input_ni[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 414.040 74.600 414.440 75.000 ;
    END
  END input_ni[6]
  PIN input_ni[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 468.760 74.600 469.160 75.000 ;
    END
  END input_ni[7]
  PIN output_no[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 4.120 0.000 4.520 0.400 ;
    END
  END output_no[0]
  PIN output_no[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 196.120 0.000 196.520 0.400 ;
    END
  END output_no[100]
  PIN output_no[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 198.040 0.000 198.440 0.400 ;
    END
  END output_no[101]
  PIN output_no[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 199.960 0.000 200.360 0.400 ;
    END
  END output_no[102]
  PIN output_no[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 201.880 0.000 202.280 0.400 ;
    END
  END output_no[103]
  PIN output_no[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 203.800 0.000 204.200 0.400 ;
    END
  END output_no[104]
  PIN output_no[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 205.720 0.000 206.120 0.400 ;
    END
  END output_no[105]
  PIN output_no[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 207.640 0.000 208.040 0.400 ;
    END
  END output_no[106]
  PIN output_no[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 209.560 0.000 209.960 0.400 ;
    END
  END output_no[107]
  PIN output_no[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 211.480 0.000 211.880 0.400 ;
    END
  END output_no[108]
  PIN output_no[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 213.400 0.000 213.800 0.400 ;
    END
  END output_no[109]
  PIN output_no[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END output_no[10]
  PIN output_no[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 215.320 0.000 215.720 0.400 ;
    END
  END output_no[110]
  PIN output_no[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 217.240 0.000 217.640 0.400 ;
    END
  END output_no[111]
  PIN output_no[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 219.160 0.000 219.560 0.400 ;
    END
  END output_no[112]
  PIN output_no[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 221.080 0.000 221.480 0.400 ;
    END
  END output_no[113]
  PIN output_no[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 223.000 0.000 223.400 0.400 ;
    END
  END output_no[114]
  PIN output_no[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 224.920 0.000 225.320 0.400 ;
    END
  END output_no[115]
  PIN output_no[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 226.840 0.000 227.240 0.400 ;
    END
  END output_no[116]
  PIN output_no[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 228.760 0.000 229.160 0.400 ;
    END
  END output_no[117]
  PIN output_no[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 230.680 0.000 231.080 0.400 ;
    END
  END output_no[118]
  PIN output_no[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 232.600 0.000 233.000 0.400 ;
    END
  END output_no[119]
  PIN output_no[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END output_no[11]
  PIN output_no[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 234.520 0.000 234.920 0.400 ;
    END
  END output_no[120]
  PIN output_no[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 236.440 0.000 236.840 0.400 ;
    END
  END output_no[121]
  PIN output_no[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 238.360 0.000 238.760 0.400 ;
    END
  END output_no[122]
  PIN output_no[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 240.280 0.000 240.680 0.400 ;
    END
  END output_no[123]
  PIN output_no[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 242.200 0.000 242.600 0.400 ;
    END
  END output_no[124]
  PIN output_no[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 244.120 0.000 244.520 0.400 ;
    END
  END output_no[125]
  PIN output_no[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 246.040 0.000 246.440 0.400 ;
    END
  END output_no[126]
  PIN output_no[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 247.960 0.000 248.360 0.400 ;
    END
  END output_no[127]
  PIN output_no[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 249.880 0.000 250.280 0.400 ;
    END
  END output_no[128]
  PIN output_no[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 251.800 0.000 252.200 0.400 ;
    END
  END output_no[129]
  PIN output_no[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END output_no[12]
  PIN output_no[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 253.720 0.000 254.120 0.400 ;
    END
  END output_no[130]
  PIN output_no[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 255.640 0.000 256.040 0.400 ;
    END
  END output_no[131]
  PIN output_no[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 257.560 0.000 257.960 0.400 ;
    END
  END output_no[132]
  PIN output_no[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 259.480 0.000 259.880 0.400 ;
    END
  END output_no[133]
  PIN output_no[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 261.400 0.000 261.800 0.400 ;
    END
  END output_no[134]
  PIN output_no[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 263.320 0.000 263.720 0.400 ;
    END
  END output_no[135]
  PIN output_no[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 265.240 0.000 265.640 0.400 ;
    END
  END output_no[136]
  PIN output_no[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 267.160 0.000 267.560 0.400 ;
    END
  END output_no[137]
  PIN output_no[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 269.080 0.000 269.480 0.400 ;
    END
  END output_no[138]
  PIN output_no[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 271.000 0.000 271.400 0.400 ;
    END
  END output_no[139]
  PIN output_no[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END output_no[13]
  PIN output_no[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 272.920 0.000 273.320 0.400 ;
    END
  END output_no[140]
  PIN output_no[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 274.840 0.000 275.240 0.400 ;
    END
  END output_no[141]
  PIN output_no[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 276.760 0.000 277.160 0.400 ;
    END
  END output_no[142]
  PIN output_no[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 278.680 0.000 279.080 0.400 ;
    END
  END output_no[143]
  PIN output_no[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 280.600 0.000 281.000 0.400 ;
    END
  END output_no[144]
  PIN output_no[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 282.520 0.000 282.920 0.400 ;
    END
  END output_no[145]
  PIN output_no[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 284.440 0.000 284.840 0.400 ;
    END
  END output_no[146]
  PIN output_no[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 286.360 0.000 286.760 0.400 ;
    END
  END output_no[147]
  PIN output_no[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 288.280 0.000 288.680 0.400 ;
    END
  END output_no[148]
  PIN output_no[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 290.200 0.000 290.600 0.400 ;
    END
  END output_no[149]
  PIN output_no[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END output_no[14]
  PIN output_no[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 292.120 0.000 292.520 0.400 ;
    END
  END output_no[150]
  PIN output_no[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 294.040 0.000 294.440 0.400 ;
    END
  END output_no[151]
  PIN output_no[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 295.960 0.000 296.360 0.400 ;
    END
  END output_no[152]
  PIN output_no[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 297.880 0.000 298.280 0.400 ;
    END
  END output_no[153]
  PIN output_no[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 299.800 0.000 300.200 0.400 ;
    END
  END output_no[154]
  PIN output_no[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 301.720 0.000 302.120 0.400 ;
    END
  END output_no[155]
  PIN output_no[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 303.640 0.000 304.040 0.400 ;
    END
  END output_no[156]
  PIN output_no[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 305.560 0.000 305.960 0.400 ;
    END
  END output_no[157]
  PIN output_no[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 307.480 0.000 307.880 0.400 ;
    END
  END output_no[158]
  PIN output_no[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 309.400 0.000 309.800 0.400 ;
    END
  END output_no[159]
  PIN output_no[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END output_no[15]
  PIN output_no[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 311.320 0.000 311.720 0.400 ;
    END
  END output_no[160]
  PIN output_no[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 313.240 0.000 313.640 0.400 ;
    END
  END output_no[161]
  PIN output_no[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 315.160 0.000 315.560 0.400 ;
    END
  END output_no[162]
  PIN output_no[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 317.080 0.000 317.480 0.400 ;
    END
  END output_no[163]
  PIN output_no[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 319.000 0.000 319.400 0.400 ;
    END
  END output_no[164]
  PIN output_no[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 320.920 0.000 321.320 0.400 ;
    END
  END output_no[165]
  PIN output_no[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 322.840 0.000 323.240 0.400 ;
    END
  END output_no[166]
  PIN output_no[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 324.760 0.000 325.160 0.400 ;
    END
  END output_no[167]
  PIN output_no[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 326.680 0.000 327.080 0.400 ;
    END
  END output_no[168]
  PIN output_no[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 328.600 0.000 329.000 0.400 ;
    END
  END output_no[169]
  PIN output_no[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END output_no[16]
  PIN output_no[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 330.520 0.000 330.920 0.400 ;
    END
  END output_no[170]
  PIN output_no[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 332.440 0.000 332.840 0.400 ;
    END
  END output_no[171]
  PIN output_no[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 334.360 0.000 334.760 0.400 ;
    END
  END output_no[172]
  PIN output_no[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 336.280 0.000 336.680 0.400 ;
    END
  END output_no[173]
  PIN output_no[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 338.200 0.000 338.600 0.400 ;
    END
  END output_no[174]
  PIN output_no[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 340.120 0.000 340.520 0.400 ;
    END
  END output_no[175]
  PIN output_no[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 342.040 0.000 342.440 0.400 ;
    END
  END output_no[176]
  PIN output_no[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 343.960 0.000 344.360 0.400 ;
    END
  END output_no[177]
  PIN output_no[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 345.880 0.000 346.280 0.400 ;
    END
  END output_no[178]
  PIN output_no[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 347.800 0.000 348.200 0.400 ;
    END
  END output_no[179]
  PIN output_no[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END output_no[17]
  PIN output_no[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 349.720 0.000 350.120 0.400 ;
    END
  END output_no[180]
  PIN output_no[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 351.640 0.000 352.040 0.400 ;
    END
  END output_no[181]
  PIN output_no[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 353.560 0.000 353.960 0.400 ;
    END
  END output_no[182]
  PIN output_no[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 355.480 0.000 355.880 0.400 ;
    END
  END output_no[183]
  PIN output_no[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 357.400 0.000 357.800 0.400 ;
    END
  END output_no[184]
  PIN output_no[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 359.320 0.000 359.720 0.400 ;
    END
  END output_no[185]
  PIN output_no[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 361.240 0.000 361.640 0.400 ;
    END
  END output_no[186]
  PIN output_no[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 363.160 0.000 363.560 0.400 ;
    END
  END output_no[187]
  PIN output_no[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 365.080 0.000 365.480 0.400 ;
    END
  END output_no[188]
  PIN output_no[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 367.000 0.000 367.400 0.400 ;
    END
  END output_no[189]
  PIN output_no[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END output_no[18]
  PIN output_no[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 368.920 0.000 369.320 0.400 ;
    END
  END output_no[190]
  PIN output_no[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 370.840 0.000 371.240 0.400 ;
    END
  END output_no[191]
  PIN output_no[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 372.760 0.000 373.160 0.400 ;
    END
  END output_no[192]
  PIN output_no[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 374.680 0.000 375.080 0.400 ;
    END
  END output_no[193]
  PIN output_no[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 376.600 0.000 377.000 0.400 ;
    END
  END output_no[194]
  PIN output_no[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 378.520 0.000 378.920 0.400 ;
    END
  END output_no[195]
  PIN output_no[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 380.440 0.000 380.840 0.400 ;
    END
  END output_no[196]
  PIN output_no[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 382.360 0.000 382.760 0.400 ;
    END
  END output_no[197]
  PIN output_no[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 384.280 0.000 384.680 0.400 ;
    END
  END output_no[198]
  PIN output_no[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 386.200 0.000 386.600 0.400 ;
    END
  END output_no[199]
  PIN output_no[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END output_no[19]
  PIN output_no[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 6.040 0.000 6.440 0.400 ;
    END
  END output_no[1]
  PIN output_no[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 388.120 0.000 388.520 0.400 ;
    END
  END output_no[200]
  PIN output_no[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 390.040 0.000 390.440 0.400 ;
    END
  END output_no[201]
  PIN output_no[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 391.960 0.000 392.360 0.400 ;
    END
  END output_no[202]
  PIN output_no[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 393.880 0.000 394.280 0.400 ;
    END
  END output_no[203]
  PIN output_no[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 395.800 0.000 396.200 0.400 ;
    END
  END output_no[204]
  PIN output_no[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 397.720 0.000 398.120 0.400 ;
    END
  END output_no[205]
  PIN output_no[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 399.640 0.000 400.040 0.400 ;
    END
  END output_no[206]
  PIN output_no[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 401.560 0.000 401.960 0.400 ;
    END
  END output_no[207]
  PIN output_no[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 403.480 0.000 403.880 0.400 ;
    END
  END output_no[208]
  PIN output_no[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 405.400 0.000 405.800 0.400 ;
    END
  END output_no[209]
  PIN output_no[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END output_no[20]
  PIN output_no[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 407.320 0.000 407.720 0.400 ;
    END
  END output_no[210]
  PIN output_no[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 409.240 0.000 409.640 0.400 ;
    END
  END output_no[211]
  PIN output_no[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 411.160 0.000 411.560 0.400 ;
    END
  END output_no[212]
  PIN output_no[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 413.080 0.000 413.480 0.400 ;
    END
  END output_no[213]
  PIN output_no[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 415.000 0.000 415.400 0.400 ;
    END
  END output_no[214]
  PIN output_no[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 416.920 0.000 417.320 0.400 ;
    END
  END output_no[215]
  PIN output_no[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 418.840 0.000 419.240 0.400 ;
    END
  END output_no[216]
  PIN output_no[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 420.760 0.000 421.160 0.400 ;
    END
  END output_no[217]
  PIN output_no[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 422.680 0.000 423.080 0.400 ;
    END
  END output_no[218]
  PIN output_no[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 424.600 0.000 425.000 0.400 ;
    END
  END output_no[219]
  PIN output_no[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END output_no[21]
  PIN output_no[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 426.520 0.000 426.920 0.400 ;
    END
  END output_no[220]
  PIN output_no[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 428.440 0.000 428.840 0.400 ;
    END
  END output_no[221]
  PIN output_no[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 430.360 0.000 430.760 0.400 ;
    END
  END output_no[222]
  PIN output_no[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 432.280 0.000 432.680 0.400 ;
    END
  END output_no[223]
  PIN output_no[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 434.200 0.000 434.600 0.400 ;
    END
  END output_no[224]
  PIN output_no[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 436.120 0.000 436.520 0.400 ;
    END
  END output_no[225]
  PIN output_no[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 438.040 0.000 438.440 0.400 ;
    END
  END output_no[226]
  PIN output_no[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 439.960 0.000 440.360 0.400 ;
    END
  END output_no[227]
  PIN output_no[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 441.880 0.000 442.280 0.400 ;
    END
  END output_no[228]
  PIN output_no[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 443.800 0.000 444.200 0.400 ;
    END
  END output_no[229]
  PIN output_no[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END output_no[22]
  PIN output_no[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 445.720 0.000 446.120 0.400 ;
    END
  END output_no[230]
  PIN output_no[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 447.640 0.000 448.040 0.400 ;
    END
  END output_no[231]
  PIN output_no[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 449.560 0.000 449.960 0.400 ;
    END
  END output_no[232]
  PIN output_no[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 451.480 0.000 451.880 0.400 ;
    END
  END output_no[233]
  PIN output_no[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 453.400 0.000 453.800 0.400 ;
    END
  END output_no[234]
  PIN output_no[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 455.320 0.000 455.720 0.400 ;
    END
  END output_no[235]
  PIN output_no[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 457.240 0.000 457.640 0.400 ;
    END
  END output_no[236]
  PIN output_no[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 459.160 0.000 459.560 0.400 ;
    END
  END output_no[237]
  PIN output_no[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 461.080 0.000 461.480 0.400 ;
    END
  END output_no[238]
  PIN output_no[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 463.000 0.000 463.400 0.400 ;
    END
  END output_no[239]
  PIN output_no[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END output_no[23]
  PIN output_no[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 464.920 0.000 465.320 0.400 ;
    END
  END output_no[240]
  PIN output_no[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 466.840 0.000 467.240 0.400 ;
    END
  END output_no[241]
  PIN output_no[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 468.760 0.000 469.160 0.400 ;
    END
  END output_no[242]
  PIN output_no[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 470.680 0.000 471.080 0.400 ;
    END
  END output_no[243]
  PIN output_no[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 472.600 0.000 473.000 0.400 ;
    END
  END output_no[244]
  PIN output_no[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 474.520 0.000 474.920 0.400 ;
    END
  END output_no[245]
  PIN output_no[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 476.440 0.000 476.840 0.400 ;
    END
  END output_no[246]
  PIN output_no[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 478.360 0.000 478.760 0.400 ;
    END
  END output_no[247]
  PIN output_no[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 480.280 0.000 480.680 0.400 ;
    END
  END output_no[248]
  PIN output_no[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 482.200 0.000 482.600 0.400 ;
    END
  END output_no[249]
  PIN output_no[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END output_no[24]
  PIN output_no[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 484.120 0.000 484.520 0.400 ;
    END
  END output_no[250]
  PIN output_no[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 486.040 0.000 486.440 0.400 ;
    END
  END output_no[251]
  PIN output_no[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 487.960 0.000 488.360 0.400 ;
    END
  END output_no[252]
  PIN output_no[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 489.880 0.000 490.280 0.400 ;
    END
  END output_no[253]
  PIN output_no[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 491.800 0.000 492.200 0.400 ;
    END
  END output_no[254]
  PIN output_no[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 493.720 0.000 494.120 0.400 ;
    END
  END output_no[255]
  PIN output_no[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END output_no[25]
  PIN output_no[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END output_no[26]
  PIN output_no[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END output_no[27]
  PIN output_no[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END output_no[28]
  PIN output_no[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END output_no[29]
  PIN output_no[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 7.960 0.000 8.360 0.400 ;
    END
  END output_no[2]
  PIN output_no[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END output_no[30]
  PIN output_no[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END output_no[31]
  PIN output_no[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END output_no[32]
  PIN output_no[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END output_no[33]
  PIN output_no[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END output_no[34]
  PIN output_no[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END output_no[35]
  PIN output_no[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END output_no[36]
  PIN output_no[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END output_no[37]
  PIN output_no[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END output_no[38]
  PIN output_no[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END output_no[39]
  PIN output_no[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 9.880 0.000 10.280 0.400 ;
    END
  END output_no[3]
  PIN output_no[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END output_no[40]
  PIN output_no[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END output_no[41]
  PIN output_no[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END output_no[42]
  PIN output_no[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END output_no[43]
  PIN output_no[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END output_no[44]
  PIN output_no[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END output_no[45]
  PIN output_no[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END output_no[46]
  PIN output_no[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END output_no[47]
  PIN output_no[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END output_no[48]
  PIN output_no[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 98.200 0.000 98.600 0.400 ;
    END
  END output_no[49]
  PIN output_no[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 11.800 0.000 12.200 0.400 ;
    END
  END output_no[4]
  PIN output_no[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 100.120 0.000 100.520 0.400 ;
    END
  END output_no[50]
  PIN output_no[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 102.040 0.000 102.440 0.400 ;
    END
  END output_no[51]
  PIN output_no[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 103.960 0.000 104.360 0.400 ;
    END
  END output_no[52]
  PIN output_no[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 105.880 0.000 106.280 0.400 ;
    END
  END output_no[53]
  PIN output_no[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 107.800 0.000 108.200 0.400 ;
    END
  END output_no[54]
  PIN output_no[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 109.720 0.000 110.120 0.400 ;
    END
  END output_no[55]
  PIN output_no[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 111.640 0.000 112.040 0.400 ;
    END
  END output_no[56]
  PIN output_no[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 113.560 0.000 113.960 0.400 ;
    END
  END output_no[57]
  PIN output_no[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 115.480 0.000 115.880 0.400 ;
    END
  END output_no[58]
  PIN output_no[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 117.400 0.000 117.800 0.400 ;
    END
  END output_no[59]
  PIN output_no[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END output_no[5]
  PIN output_no[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 119.320 0.000 119.720 0.400 ;
    END
  END output_no[60]
  PIN output_no[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 121.240 0.000 121.640 0.400 ;
    END
  END output_no[61]
  PIN output_no[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 123.160 0.000 123.560 0.400 ;
    END
  END output_no[62]
  PIN output_no[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 125.080 0.000 125.480 0.400 ;
    END
  END output_no[63]
  PIN output_no[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.000 0.000 127.400 0.400 ;
    END
  END output_no[64]
  PIN output_no[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 128.920 0.000 129.320 0.400 ;
    END
  END output_no[65]
  PIN output_no[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 130.840 0.000 131.240 0.400 ;
    END
  END output_no[66]
  PIN output_no[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 132.760 0.000 133.160 0.400 ;
    END
  END output_no[67]
  PIN output_no[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 134.680 0.000 135.080 0.400 ;
    END
  END output_no[68]
  PIN output_no[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 136.600 0.000 137.000 0.400 ;
    END
  END output_no[69]
  PIN output_no[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END output_no[6]
  PIN output_no[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 138.520 0.000 138.920 0.400 ;
    END
  END output_no[70]
  PIN output_no[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 140.440 0.000 140.840 0.400 ;
    END
  END output_no[71]
  PIN output_no[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.360 0.000 142.760 0.400 ;
    END
  END output_no[72]
  PIN output_no[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.280 0.000 144.680 0.400 ;
    END
  END output_no[73]
  PIN output_no[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.200 0.000 146.600 0.400 ;
    END
  END output_no[74]
  PIN output_no[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 0.000 148.520 0.400 ;
    END
  END output_no[75]
  PIN output_no[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 150.040 0.000 150.440 0.400 ;
    END
  END output_no[76]
  PIN output_no[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.960 0.000 152.360 0.400 ;
    END
  END output_no[77]
  PIN output_no[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.880 0.000 154.280 0.400 ;
    END
  END output_no[78]
  PIN output_no[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.800 0.000 156.200 0.400 ;
    END
  END output_no[79]
  PIN output_no[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END output_no[7]
  PIN output_no[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.720 0.000 158.120 0.400 ;
    END
  END output_no[80]
  PIN output_no[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 159.640 0.000 160.040 0.400 ;
    END
  END output_no[81]
  PIN output_no[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 0.000 161.960 0.400 ;
    END
  END output_no[82]
  PIN output_no[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 163.480 0.000 163.880 0.400 ;
    END
  END output_no[83]
  PIN output_no[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 165.400 0.000 165.800 0.400 ;
    END
  END output_no[84]
  PIN output_no[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 167.320 0.000 167.720 0.400 ;
    END
  END output_no[85]
  PIN output_no[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 169.240 0.000 169.640 0.400 ;
    END
  END output_no[86]
  PIN output_no[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 171.160 0.000 171.560 0.400 ;
    END
  END output_no[87]
  PIN output_no[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 173.080 0.000 173.480 0.400 ;
    END
  END output_no[88]
  PIN output_no[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 175.000 0.000 175.400 0.400 ;
    END
  END output_no[89]
  PIN output_no[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END output_no[8]
  PIN output_no[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 176.920 0.000 177.320 0.400 ;
    END
  END output_no[90]
  PIN output_no[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 178.840 0.000 179.240 0.400 ;
    END
  END output_no[91]
  PIN output_no[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 180.760 0.000 181.160 0.400 ;
    END
  END output_no[92]
  PIN output_no[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 182.680 0.000 183.080 0.400 ;
    END
  END output_no[93]
  PIN output_no[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 184.600 0.000 185.000 0.400 ;
    END
  END output_no[94]
  PIN output_no[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 186.520 0.000 186.920 0.400 ;
    END
  END output_no[95]
  PIN output_no[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 188.440 0.000 188.840 0.400 ;
    END
  END output_no[96]
  PIN output_no[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 190.360 0.000 190.760 0.400 ;
    END
  END output_no[97]
  PIN output_no[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 192.280 0.000 192.680 0.400 ;
    END
  END output_no[98]
  PIN output_no[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 194.200 0.000 194.600 0.400 ;
    END
  END output_no[99]
  PIN output_no[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END output_no[9]
  PIN output_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 5.080 0.000 5.480 0.400 ;
    END
  END output_o[0]
  PIN output_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 197.080 0.000 197.480 0.400 ;
    END
  END output_o[100]
  PIN output_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 199.000 0.000 199.400 0.400 ;
    END
  END output_o[101]
  PIN output_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 200.920 0.000 201.320 0.400 ;
    END
  END output_o[102]
  PIN output_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 202.840 0.000 203.240 0.400 ;
    END
  END output_o[103]
  PIN output_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 204.760 0.000 205.160 0.400 ;
    END
  END output_o[104]
  PIN output_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 206.680 0.000 207.080 0.400 ;
    END
  END output_o[105]
  PIN output_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 208.600 0.000 209.000 0.400 ;
    END
  END output_o[106]
  PIN output_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 210.520 0.000 210.920 0.400 ;
    END
  END output_o[107]
  PIN output_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 212.440 0.000 212.840 0.400 ;
    END
  END output_o[108]
  PIN output_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 214.360 0.000 214.760 0.400 ;
    END
  END output_o[109]
  PIN output_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 24.280 0.000 24.680 0.400 ;
    END
  END output_o[10]
  PIN output_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 216.280 0.000 216.680 0.400 ;
    END
  END output_o[110]
  PIN output_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 218.200 0.000 218.600 0.400 ;
    END
  END output_o[111]
  PIN output_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 220.120 0.000 220.520 0.400 ;
    END
  END output_o[112]
  PIN output_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 222.040 0.000 222.440 0.400 ;
    END
  END output_o[113]
  PIN output_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 223.960 0.000 224.360 0.400 ;
    END
  END output_o[114]
  PIN output_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 225.880 0.000 226.280 0.400 ;
    END
  END output_o[115]
  PIN output_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 227.800 0.000 228.200 0.400 ;
    END
  END output_o[116]
  PIN output_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 229.720 0.000 230.120 0.400 ;
    END
  END output_o[117]
  PIN output_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 231.640 0.000 232.040 0.400 ;
    END
  END output_o[118]
  PIN output_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 233.560 0.000 233.960 0.400 ;
    END
  END output_o[119]
  PIN output_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 0.000 26.600 0.400 ;
    END
  END output_o[11]
  PIN output_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 235.480 0.000 235.880 0.400 ;
    END
  END output_o[120]
  PIN output_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 237.400 0.000 237.800 0.400 ;
    END
  END output_o[121]
  PIN output_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 239.320 0.000 239.720 0.400 ;
    END
  END output_o[122]
  PIN output_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 241.240 0.000 241.640 0.400 ;
    END
  END output_o[123]
  PIN output_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 243.160 0.000 243.560 0.400 ;
    END
  END output_o[124]
  PIN output_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 245.080 0.000 245.480 0.400 ;
    END
  END output_o[125]
  PIN output_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 247.000 0.000 247.400 0.400 ;
    END
  END output_o[126]
  PIN output_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 248.920 0.000 249.320 0.400 ;
    END
  END output_o[127]
  PIN output_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 250.840 0.000 251.240 0.400 ;
    END
  END output_o[128]
  PIN output_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 252.760 0.000 253.160 0.400 ;
    END
  END output_o[129]
  PIN output_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 0.000 28.520 0.400 ;
    END
  END output_o[12]
  PIN output_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 254.680 0.000 255.080 0.400 ;
    END
  END output_o[130]
  PIN output_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 256.600 0.000 257.000 0.400 ;
    END
  END output_o[131]
  PIN output_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 258.520 0.000 258.920 0.400 ;
    END
  END output_o[132]
  PIN output_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 260.440 0.000 260.840 0.400 ;
    END
  END output_o[133]
  PIN output_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 262.360 0.000 262.760 0.400 ;
    END
  END output_o[134]
  PIN output_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 264.280 0.000 264.680 0.400 ;
    END
  END output_o[135]
  PIN output_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 266.200 0.000 266.600 0.400 ;
    END
  END output_o[136]
  PIN output_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 268.120 0.000 268.520 0.400 ;
    END
  END output_o[137]
  PIN output_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 270.040 0.000 270.440 0.400 ;
    END
  END output_o[138]
  PIN output_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 271.960 0.000 272.360 0.400 ;
    END
  END output_o[139]
  PIN output_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.040 0.000 30.440 0.400 ;
    END
  END output_o[13]
  PIN output_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 273.880 0.000 274.280 0.400 ;
    END
  END output_o[140]
  PIN output_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 0.000 276.200 0.400 ;
    END
  END output_o[141]
  PIN output_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 277.720 0.000 278.120 0.400 ;
    END
  END output_o[142]
  PIN output_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 279.640 0.000 280.040 0.400 ;
    END
  END output_o[143]
  PIN output_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 281.560 0.000 281.960 0.400 ;
    END
  END output_o[144]
  PIN output_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 283.480 0.000 283.880 0.400 ;
    END
  END output_o[145]
  PIN output_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 285.400 0.000 285.800 0.400 ;
    END
  END output_o[146]
  PIN output_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 287.320 0.000 287.720 0.400 ;
    END
  END output_o[147]
  PIN output_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 289.240 0.000 289.640 0.400 ;
    END
  END output_o[148]
  PIN output_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 291.160 0.000 291.560 0.400 ;
    END
  END output_o[149]
  PIN output_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 0.000 32.360 0.400 ;
    END
  END output_o[14]
  PIN output_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 293.080 0.000 293.480 0.400 ;
    END
  END output_o[150]
  PIN output_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 295.000 0.000 295.400 0.400 ;
    END
  END output_o[151]
  PIN output_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 296.920 0.000 297.320 0.400 ;
    END
  END output_o[152]
  PIN output_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 298.840 0.000 299.240 0.400 ;
    END
  END output_o[153]
  PIN output_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 300.760 0.000 301.160 0.400 ;
    END
  END output_o[154]
  PIN output_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 302.680 0.000 303.080 0.400 ;
    END
  END output_o[155]
  PIN output_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 304.600 0.000 305.000 0.400 ;
    END
  END output_o[156]
  PIN output_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 306.520 0.000 306.920 0.400 ;
    END
  END output_o[157]
  PIN output_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 308.440 0.000 308.840 0.400 ;
    END
  END output_o[158]
  PIN output_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 310.360 0.000 310.760 0.400 ;
    END
  END output_o[159]
  PIN output_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 0.000 34.280 0.400 ;
    END
  END output_o[15]
  PIN output_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 312.280 0.000 312.680 0.400 ;
    END
  END output_o[160]
  PIN output_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 314.200 0.000 314.600 0.400 ;
    END
  END output_o[161]
  PIN output_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 316.120 0.000 316.520 0.400 ;
    END
  END output_o[162]
  PIN output_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 318.040 0.000 318.440 0.400 ;
    END
  END output_o[163]
  PIN output_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 319.960 0.000 320.360 0.400 ;
    END
  END output_o[164]
  PIN output_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 321.880 0.000 322.280 0.400 ;
    END
  END output_o[165]
  PIN output_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 323.800 0.000 324.200 0.400 ;
    END
  END output_o[166]
  PIN output_o[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 325.720 0.000 326.120 0.400 ;
    END
  END output_o[167]
  PIN output_o[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 327.640 0.000 328.040 0.400 ;
    END
  END output_o[168]
  PIN output_o[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 329.560 0.000 329.960 0.400 ;
    END
  END output_o[169]
  PIN output_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 0.000 36.200 0.400 ;
    END
  END output_o[16]
  PIN output_o[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 331.480 0.000 331.880 0.400 ;
    END
  END output_o[170]
  PIN output_o[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 333.400 0.000 333.800 0.400 ;
    END
  END output_o[171]
  PIN output_o[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 335.320 0.000 335.720 0.400 ;
    END
  END output_o[172]
  PIN output_o[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 337.240 0.000 337.640 0.400 ;
    END
  END output_o[173]
  PIN output_o[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 339.160 0.000 339.560 0.400 ;
    END
  END output_o[174]
  PIN output_o[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 341.080 0.000 341.480 0.400 ;
    END
  END output_o[175]
  PIN output_o[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 343.000 0.000 343.400 0.400 ;
    END
  END output_o[176]
  PIN output_o[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 344.920 0.000 345.320 0.400 ;
    END
  END output_o[177]
  PIN output_o[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 346.840 0.000 347.240 0.400 ;
    END
  END output_o[178]
  PIN output_o[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 348.760 0.000 349.160 0.400 ;
    END
  END output_o[179]
  PIN output_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END output_o[17]
  PIN output_o[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 350.680 0.000 351.080 0.400 ;
    END
  END output_o[180]
  PIN output_o[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 352.600 0.000 353.000 0.400 ;
    END
  END output_o[181]
  PIN output_o[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 354.520 0.000 354.920 0.400 ;
    END
  END output_o[182]
  PIN output_o[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 356.440 0.000 356.840 0.400 ;
    END
  END output_o[183]
  PIN output_o[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 358.360 0.000 358.760 0.400 ;
    END
  END output_o[184]
  PIN output_o[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 360.280 0.000 360.680 0.400 ;
    END
  END output_o[185]
  PIN output_o[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 362.200 0.000 362.600 0.400 ;
    END
  END output_o[186]
  PIN output_o[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 364.120 0.000 364.520 0.400 ;
    END
  END output_o[187]
  PIN output_o[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 366.040 0.000 366.440 0.400 ;
    END
  END output_o[188]
  PIN output_o[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 367.960 0.000 368.360 0.400 ;
    END
  END output_o[189]
  PIN output_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END output_o[18]
  PIN output_o[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 369.880 0.000 370.280 0.400 ;
    END
  END output_o[190]
  PIN output_o[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 371.800 0.000 372.200 0.400 ;
    END
  END output_o[191]
  PIN output_o[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 373.720 0.000 374.120 0.400 ;
    END
  END output_o[192]
  PIN output_o[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 375.640 0.000 376.040 0.400 ;
    END
  END output_o[193]
  PIN output_o[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 377.560 0.000 377.960 0.400 ;
    END
  END output_o[194]
  PIN output_o[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 379.480 0.000 379.880 0.400 ;
    END
  END output_o[195]
  PIN output_o[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 381.400 0.000 381.800 0.400 ;
    END
  END output_o[196]
  PIN output_o[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 383.320 0.000 383.720 0.400 ;
    END
  END output_o[197]
  PIN output_o[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 385.240 0.000 385.640 0.400 ;
    END
  END output_o[198]
  PIN output_o[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 387.160 0.000 387.560 0.400 ;
    END
  END output_o[199]
  PIN output_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END output_o[19]
  PIN output_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 7.000 0.000 7.400 0.400 ;
    END
  END output_o[1]
  PIN output_o[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 389.080 0.000 389.480 0.400 ;
    END
  END output_o[200]
  PIN output_o[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 391.000 0.000 391.400 0.400 ;
    END
  END output_o[201]
  PIN output_o[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 392.920 0.000 393.320 0.400 ;
    END
  END output_o[202]
  PIN output_o[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 394.840 0.000 395.240 0.400 ;
    END
  END output_o[203]
  PIN output_o[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 396.760 0.000 397.160 0.400 ;
    END
  END output_o[204]
  PIN output_o[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 398.680 0.000 399.080 0.400 ;
    END
  END output_o[205]
  PIN output_o[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 400.600 0.000 401.000 0.400 ;
    END
  END output_o[206]
  PIN output_o[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 402.520 0.000 402.920 0.400 ;
    END
  END output_o[207]
  PIN output_o[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 404.440 0.000 404.840 0.400 ;
    END
  END output_o[208]
  PIN output_o[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 406.360 0.000 406.760 0.400 ;
    END
  END output_o[209]
  PIN output_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END output_o[20]
  PIN output_o[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 408.280 0.000 408.680 0.400 ;
    END
  END output_o[210]
  PIN output_o[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 410.200 0.000 410.600 0.400 ;
    END
  END output_o[211]
  PIN output_o[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 412.120 0.000 412.520 0.400 ;
    END
  END output_o[212]
  PIN output_o[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 414.040 0.000 414.440 0.400 ;
    END
  END output_o[213]
  PIN output_o[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 415.960 0.000 416.360 0.400 ;
    END
  END output_o[214]
  PIN output_o[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 417.880 0.000 418.280 0.400 ;
    END
  END output_o[215]
  PIN output_o[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 419.800 0.000 420.200 0.400 ;
    END
  END output_o[216]
  PIN output_o[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 421.720 0.000 422.120 0.400 ;
    END
  END output_o[217]
  PIN output_o[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 423.640 0.000 424.040 0.400 ;
    END
  END output_o[218]
  PIN output_o[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 425.560 0.000 425.960 0.400 ;
    END
  END output_o[219]
  PIN output_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END output_o[21]
  PIN output_o[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 427.480 0.000 427.880 0.400 ;
    END
  END output_o[220]
  PIN output_o[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 429.400 0.000 429.800 0.400 ;
    END
  END output_o[221]
  PIN output_o[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 431.320 0.000 431.720 0.400 ;
    END
  END output_o[222]
  PIN output_o[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 433.240 0.000 433.640 0.400 ;
    END
  END output_o[223]
  PIN output_o[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 435.160 0.000 435.560 0.400 ;
    END
  END output_o[224]
  PIN output_o[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 437.080 0.000 437.480 0.400 ;
    END
  END output_o[225]
  PIN output_o[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 439.000 0.000 439.400 0.400 ;
    END
  END output_o[226]
  PIN output_o[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 440.920 0.000 441.320 0.400 ;
    END
  END output_o[227]
  PIN output_o[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 442.840 0.000 443.240 0.400 ;
    END
  END output_o[228]
  PIN output_o[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 444.760 0.000 445.160 0.400 ;
    END
  END output_o[229]
  PIN output_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.720 0.400 ;
    END
  END output_o[22]
  PIN output_o[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 446.680 0.000 447.080 0.400 ;
    END
  END output_o[230]
  PIN output_o[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 448.600 0.000 449.000 0.400 ;
    END
  END output_o[231]
  PIN output_o[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 450.520 0.000 450.920 0.400 ;
    END
  END output_o[232]
  PIN output_o[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 452.440 0.000 452.840 0.400 ;
    END
  END output_o[233]
  PIN output_o[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 454.360 0.000 454.760 0.400 ;
    END
  END output_o[234]
  PIN output_o[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 456.280 0.000 456.680 0.400 ;
    END
  END output_o[235]
  PIN output_o[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 458.200 0.000 458.600 0.400 ;
    END
  END output_o[236]
  PIN output_o[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 460.120 0.000 460.520 0.400 ;
    END
  END output_o[237]
  PIN output_o[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 462.040 0.000 462.440 0.400 ;
    END
  END output_o[238]
  PIN output_o[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 463.960 0.000 464.360 0.400 ;
    END
  END output_o[239]
  PIN output_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END output_o[23]
  PIN output_o[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 465.880 0.000 466.280 0.400 ;
    END
  END output_o[240]
  PIN output_o[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 467.800 0.000 468.200 0.400 ;
    END
  END output_o[241]
  PIN output_o[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 469.720 0.000 470.120 0.400 ;
    END
  END output_o[242]
  PIN output_o[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 471.640 0.000 472.040 0.400 ;
    END
  END output_o[243]
  PIN output_o[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 473.560 0.000 473.960 0.400 ;
    END
  END output_o[244]
  PIN output_o[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 475.480 0.000 475.880 0.400 ;
    END
  END output_o[245]
  PIN output_o[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 477.400 0.000 477.800 0.400 ;
    END
  END output_o[246]
  PIN output_o[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 479.320 0.000 479.720 0.400 ;
    END
  END output_o[247]
  PIN output_o[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 481.240 0.000 481.640 0.400 ;
    END
  END output_o[248]
  PIN output_o[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 483.160 0.000 483.560 0.400 ;
    END
  END output_o[249]
  PIN output_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END output_o[24]
  PIN output_o[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 485.080 0.000 485.480 0.400 ;
    END
  END output_o[250]
  PIN output_o[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 487.000 0.000 487.400 0.400 ;
    END
  END output_o[251]
  PIN output_o[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 488.920 0.000 489.320 0.400 ;
    END
  END output_o[252]
  PIN output_o[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 490.840 0.000 491.240 0.400 ;
    END
  END output_o[253]
  PIN output_o[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 492.760 0.000 493.160 0.400 ;
    END
  END output_o[254]
  PIN output_o[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 494.680 0.000 495.080 0.400 ;
    END
  END output_o[255]
  PIN output_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 0.000 53.480 0.400 ;
    END
  END output_o[25]
  PIN output_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END output_o[26]
  PIN output_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END output_o[27]
  PIN output_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END output_o[28]
  PIN output_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END output_o[29]
  PIN output_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 8.920 0.000 9.320 0.400 ;
    END
  END output_o[2]
  PIN output_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END output_o[30]
  PIN output_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END output_o[31]
  PIN output_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END output_o[32]
  PIN output_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END output_o[33]
  PIN output_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END output_o[34]
  PIN output_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END output_o[35]
  PIN output_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END output_o[36]
  PIN output_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END output_o[37]
  PIN output_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END output_o[38]
  PIN output_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END output_o[39]
  PIN output_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.840 0.000 11.240 0.400 ;
    END
  END output_o[3]
  PIN output_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END output_o[40]
  PIN output_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END output_o[41]
  PIN output_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END output_o[42]
  PIN output_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END output_o[43]
  PIN output_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END output_o[44]
  PIN output_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END output_o[45]
  PIN output_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END output_o[46]
  PIN output_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END output_o[47]
  PIN output_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END output_o[48]
  PIN output_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 99.160 0.000 99.560 0.400 ;
    END
  END output_o[49]
  PIN output_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 0.000 13.160 0.400 ;
    END
  END output_o[4]
  PIN output_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 0.000 101.480 0.400 ;
    END
  END output_o[50]
  PIN output_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 103.000 0.000 103.400 0.400 ;
    END
  END output_o[51]
  PIN output_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 104.920 0.000 105.320 0.400 ;
    END
  END output_o[52]
  PIN output_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 106.840 0.000 107.240 0.400 ;
    END
  END output_o[53]
  PIN output_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 108.760 0.000 109.160 0.400 ;
    END
  END output_o[54]
  PIN output_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 110.680 0.000 111.080 0.400 ;
    END
  END output_o[55]
  PIN output_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 112.600 0.000 113.000 0.400 ;
    END
  END output_o[56]
  PIN output_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 114.520 0.000 114.920 0.400 ;
    END
  END output_o[57]
  PIN output_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 116.440 0.000 116.840 0.400 ;
    END
  END output_o[58]
  PIN output_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 118.360 0.000 118.760 0.400 ;
    END
  END output_o[59]
  PIN output_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 0.000 15.080 0.400 ;
    END
  END output_o[5]
  PIN output_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 120.280 0.000 120.680 0.400 ;
    END
  END output_o[60]
  PIN output_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 122.200 0.000 122.600 0.400 ;
    END
  END output_o[61]
  PIN output_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 124.120 0.000 124.520 0.400 ;
    END
  END output_o[62]
  PIN output_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.040 0.000 126.440 0.400 ;
    END
  END output_o[63]
  PIN output_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.960 0.000 128.360 0.400 ;
    END
  END output_o[64]
  PIN output_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 129.880 0.000 130.280 0.400 ;
    END
  END output_o[65]
  PIN output_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 131.800 0.000 132.200 0.400 ;
    END
  END output_o[66]
  PIN output_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.720 0.000 134.120 0.400 ;
    END
  END output_o[67]
  PIN output_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 135.640 0.000 136.040 0.400 ;
    END
  END output_o[68]
  PIN output_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.560 0.000 137.960 0.400 ;
    END
  END output_o[69]
  PIN output_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.600 0.000 17.000 0.400 ;
    END
  END output_o[6]
  PIN output_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.480 0.000 139.880 0.400 ;
    END
  END output_o[70]
  PIN output_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.400 0.000 141.800 0.400 ;
    END
  END output_o[71]
  PIN output_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 143.320 0.000 143.720 0.400 ;
    END
  END output_o[72]
  PIN output_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 145.240 0.000 145.640 0.400 ;
    END
  END output_o[73]
  PIN output_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 147.160 0.000 147.560 0.400 ;
    END
  END output_o[74]
  PIN output_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 149.080 0.000 149.480 0.400 ;
    END
  END output_o[75]
  PIN output_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.000 0.000 151.400 0.400 ;
    END
  END output_o[76]
  PIN output_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 152.920 0.000 153.320 0.400 ;
    END
  END output_o[77]
  PIN output_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 0.000 155.240 0.400 ;
    END
  END output_o[78]
  PIN output_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 156.760 0.000 157.160 0.400 ;
    END
  END output_o[79]
  PIN output_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 18.520 0.000 18.920 0.400 ;
    END
  END output_o[7]
  PIN output_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 158.680 0.000 159.080 0.400 ;
    END
  END output_o[80]
  PIN output_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 160.600 0.000 161.000 0.400 ;
    END
  END output_o[81]
  PIN output_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.520 0.000 162.920 0.400 ;
    END
  END output_o[82]
  PIN output_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.440 0.000 164.840 0.400 ;
    END
  END output_o[83]
  PIN output_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.360 0.000 166.760 0.400 ;
    END
  END output_o[84]
  PIN output_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 168.280 0.000 168.680 0.400 ;
    END
  END output_o[85]
  PIN output_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 170.200 0.000 170.600 0.400 ;
    END
  END output_o[86]
  PIN output_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 172.120 0.000 172.520 0.400 ;
    END
  END output_o[87]
  PIN output_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 174.040 0.000 174.440 0.400 ;
    END
  END output_o[88]
  PIN output_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 175.960 0.000 176.360 0.400 ;
    END
  END output_o[89]
  PIN output_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END output_o[8]
  PIN output_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 177.880 0.000 178.280 0.400 ;
    END
  END output_o[90]
  PIN output_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 179.800 0.000 180.200 0.400 ;
    END
  END output_o[91]
  PIN output_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 181.720 0.000 182.120 0.400 ;
    END
  END output_o[92]
  PIN output_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 183.640 0.000 184.040 0.400 ;
    END
  END output_o[93]
  PIN output_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 185.560 0.000 185.960 0.400 ;
    END
  END output_o[94]
  PIN output_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 187.480 0.000 187.880 0.400 ;
    END
  END output_o[95]
  PIN output_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 189.400 0.000 189.800 0.400 ;
    END
  END output_o[96]
  PIN output_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 191.320 0.000 191.720 0.400 ;
    END
  END output_o[97]
  PIN output_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 193.240 0.000 193.640 0.400 ;
    END
  END output_o[98]
  PIN output_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 195.160 0.000 195.560 0.400 ;
    END
  END output_o[99]
  PIN output_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 22.360 0.000 22.760 0.400 ;
    END
  END output_o[9]
  OBS
      LAYER GatPoly ;
        RECT 5.760 14.970 493.920 56.850 ;
      LAYER Metal1 ;
        RECT 5.760 14.900 493.920 56.920 ;
      LAYER Metal2 ;
        RECT 4.220 74.390 30.790 74.600 ;
        RECT 31.610 74.390 85.510 74.600 ;
        RECT 86.330 74.390 140.230 74.600 ;
        RECT 141.050 74.390 194.950 74.600 ;
        RECT 195.770 74.390 249.670 74.600 ;
        RECT 250.490 74.390 304.390 74.600 ;
        RECT 305.210 74.390 359.110 74.600 ;
        RECT 359.930 74.390 413.830 74.600 ;
        RECT 414.650 74.390 468.550 74.600 ;
        RECT 469.370 74.390 494.985 74.600 ;
        RECT 4.220 0.610 494.985 74.390 ;
        RECT 4.730 0.320 4.870 0.610 ;
        RECT 5.690 0.320 5.830 0.610 ;
        RECT 6.650 0.320 6.790 0.610 ;
        RECT 7.610 0.320 7.750 0.610 ;
        RECT 8.570 0.320 8.710 0.610 ;
        RECT 9.530 0.320 9.670 0.610 ;
        RECT 10.490 0.320 10.630 0.610 ;
        RECT 11.450 0.320 11.590 0.610 ;
        RECT 12.410 0.320 12.550 0.610 ;
        RECT 13.370 0.320 13.510 0.610 ;
        RECT 14.330 0.320 14.470 0.610 ;
        RECT 15.290 0.320 15.430 0.610 ;
        RECT 16.250 0.320 16.390 0.610 ;
        RECT 17.210 0.320 17.350 0.610 ;
        RECT 18.170 0.320 18.310 0.610 ;
        RECT 19.130 0.320 19.270 0.610 ;
        RECT 20.090 0.320 20.230 0.610 ;
        RECT 21.050 0.320 21.190 0.610 ;
        RECT 22.010 0.320 22.150 0.610 ;
        RECT 22.970 0.320 23.110 0.610 ;
        RECT 23.930 0.320 24.070 0.610 ;
        RECT 24.890 0.320 25.030 0.610 ;
        RECT 25.850 0.320 25.990 0.610 ;
        RECT 26.810 0.320 26.950 0.610 ;
        RECT 27.770 0.320 27.910 0.610 ;
        RECT 28.730 0.320 28.870 0.610 ;
        RECT 29.690 0.320 29.830 0.610 ;
        RECT 30.650 0.320 30.790 0.610 ;
        RECT 31.610 0.320 31.750 0.610 ;
        RECT 32.570 0.320 32.710 0.610 ;
        RECT 33.530 0.320 33.670 0.610 ;
        RECT 34.490 0.320 34.630 0.610 ;
        RECT 35.450 0.320 35.590 0.610 ;
        RECT 36.410 0.320 36.550 0.610 ;
        RECT 37.370 0.320 37.510 0.610 ;
        RECT 38.330 0.320 38.470 0.610 ;
        RECT 39.290 0.320 39.430 0.610 ;
        RECT 40.250 0.320 40.390 0.610 ;
        RECT 41.210 0.320 41.350 0.610 ;
        RECT 42.170 0.320 42.310 0.610 ;
        RECT 43.130 0.320 43.270 0.610 ;
        RECT 44.090 0.320 44.230 0.610 ;
        RECT 45.050 0.320 45.190 0.610 ;
        RECT 46.010 0.320 46.150 0.610 ;
        RECT 46.970 0.320 47.110 0.610 ;
        RECT 47.930 0.320 48.070 0.610 ;
        RECT 48.890 0.320 49.030 0.610 ;
        RECT 49.850 0.320 49.990 0.610 ;
        RECT 50.810 0.320 50.950 0.610 ;
        RECT 51.770 0.320 51.910 0.610 ;
        RECT 52.730 0.320 52.870 0.610 ;
        RECT 53.690 0.320 53.830 0.610 ;
        RECT 54.650 0.320 54.790 0.610 ;
        RECT 55.610 0.320 55.750 0.610 ;
        RECT 56.570 0.320 56.710 0.610 ;
        RECT 57.530 0.320 57.670 0.610 ;
        RECT 58.490 0.320 58.630 0.610 ;
        RECT 59.450 0.320 59.590 0.610 ;
        RECT 60.410 0.320 60.550 0.610 ;
        RECT 61.370 0.320 61.510 0.610 ;
        RECT 62.330 0.320 62.470 0.610 ;
        RECT 63.290 0.320 63.430 0.610 ;
        RECT 64.250 0.320 64.390 0.610 ;
        RECT 65.210 0.320 65.350 0.610 ;
        RECT 66.170 0.320 66.310 0.610 ;
        RECT 67.130 0.320 67.270 0.610 ;
        RECT 68.090 0.320 68.230 0.610 ;
        RECT 69.050 0.320 69.190 0.610 ;
        RECT 70.010 0.320 70.150 0.610 ;
        RECT 70.970 0.320 71.110 0.610 ;
        RECT 71.930 0.320 72.070 0.610 ;
        RECT 72.890 0.320 73.030 0.610 ;
        RECT 73.850 0.320 73.990 0.610 ;
        RECT 74.810 0.320 74.950 0.610 ;
        RECT 75.770 0.320 75.910 0.610 ;
        RECT 76.730 0.320 76.870 0.610 ;
        RECT 77.690 0.320 77.830 0.610 ;
        RECT 78.650 0.320 78.790 0.610 ;
        RECT 79.610 0.320 79.750 0.610 ;
        RECT 80.570 0.320 80.710 0.610 ;
        RECT 81.530 0.320 81.670 0.610 ;
        RECT 82.490 0.320 82.630 0.610 ;
        RECT 83.450 0.320 83.590 0.610 ;
        RECT 84.410 0.320 84.550 0.610 ;
        RECT 85.370 0.320 85.510 0.610 ;
        RECT 86.330 0.320 86.470 0.610 ;
        RECT 87.290 0.320 87.430 0.610 ;
        RECT 88.250 0.320 88.390 0.610 ;
        RECT 89.210 0.320 89.350 0.610 ;
        RECT 90.170 0.320 90.310 0.610 ;
        RECT 91.130 0.320 91.270 0.610 ;
        RECT 92.090 0.320 92.230 0.610 ;
        RECT 93.050 0.320 93.190 0.610 ;
        RECT 94.010 0.320 94.150 0.610 ;
        RECT 94.970 0.320 95.110 0.610 ;
        RECT 95.930 0.320 96.070 0.610 ;
        RECT 96.890 0.320 97.030 0.610 ;
        RECT 97.850 0.320 97.990 0.610 ;
        RECT 98.810 0.320 98.950 0.610 ;
        RECT 99.770 0.320 99.910 0.610 ;
        RECT 100.730 0.320 100.870 0.610 ;
        RECT 101.690 0.320 101.830 0.610 ;
        RECT 102.650 0.320 102.790 0.610 ;
        RECT 103.610 0.320 103.750 0.610 ;
        RECT 104.570 0.320 104.710 0.610 ;
        RECT 105.530 0.320 105.670 0.610 ;
        RECT 106.490 0.320 106.630 0.610 ;
        RECT 107.450 0.320 107.590 0.610 ;
        RECT 108.410 0.320 108.550 0.610 ;
        RECT 109.370 0.320 109.510 0.610 ;
        RECT 110.330 0.320 110.470 0.610 ;
        RECT 111.290 0.320 111.430 0.610 ;
        RECT 112.250 0.320 112.390 0.610 ;
        RECT 113.210 0.320 113.350 0.610 ;
        RECT 114.170 0.320 114.310 0.610 ;
        RECT 115.130 0.320 115.270 0.610 ;
        RECT 116.090 0.320 116.230 0.610 ;
        RECT 117.050 0.320 117.190 0.610 ;
        RECT 118.010 0.320 118.150 0.610 ;
        RECT 118.970 0.320 119.110 0.610 ;
        RECT 119.930 0.320 120.070 0.610 ;
        RECT 120.890 0.320 121.030 0.610 ;
        RECT 121.850 0.320 121.990 0.610 ;
        RECT 122.810 0.320 122.950 0.610 ;
        RECT 123.770 0.320 123.910 0.610 ;
        RECT 124.730 0.320 124.870 0.610 ;
        RECT 125.690 0.320 125.830 0.610 ;
        RECT 126.650 0.320 126.790 0.610 ;
        RECT 127.610 0.320 127.750 0.610 ;
        RECT 128.570 0.320 128.710 0.610 ;
        RECT 129.530 0.320 129.670 0.610 ;
        RECT 130.490 0.320 130.630 0.610 ;
        RECT 131.450 0.320 131.590 0.610 ;
        RECT 132.410 0.320 132.550 0.610 ;
        RECT 133.370 0.320 133.510 0.610 ;
        RECT 134.330 0.320 134.470 0.610 ;
        RECT 135.290 0.320 135.430 0.610 ;
        RECT 136.250 0.320 136.390 0.610 ;
        RECT 137.210 0.320 137.350 0.610 ;
        RECT 138.170 0.320 138.310 0.610 ;
        RECT 139.130 0.320 139.270 0.610 ;
        RECT 140.090 0.320 140.230 0.610 ;
        RECT 141.050 0.320 141.190 0.610 ;
        RECT 142.010 0.320 142.150 0.610 ;
        RECT 142.970 0.320 143.110 0.610 ;
        RECT 143.930 0.320 144.070 0.610 ;
        RECT 144.890 0.320 145.030 0.610 ;
        RECT 145.850 0.320 145.990 0.610 ;
        RECT 146.810 0.320 146.950 0.610 ;
        RECT 147.770 0.320 147.910 0.610 ;
        RECT 148.730 0.320 148.870 0.610 ;
        RECT 149.690 0.320 149.830 0.610 ;
        RECT 150.650 0.320 150.790 0.610 ;
        RECT 151.610 0.320 151.750 0.610 ;
        RECT 152.570 0.320 152.710 0.610 ;
        RECT 153.530 0.320 153.670 0.610 ;
        RECT 154.490 0.320 154.630 0.610 ;
        RECT 155.450 0.320 155.590 0.610 ;
        RECT 156.410 0.320 156.550 0.610 ;
        RECT 157.370 0.320 157.510 0.610 ;
        RECT 158.330 0.320 158.470 0.610 ;
        RECT 159.290 0.320 159.430 0.610 ;
        RECT 160.250 0.320 160.390 0.610 ;
        RECT 161.210 0.320 161.350 0.610 ;
        RECT 162.170 0.320 162.310 0.610 ;
        RECT 163.130 0.320 163.270 0.610 ;
        RECT 164.090 0.320 164.230 0.610 ;
        RECT 165.050 0.320 165.190 0.610 ;
        RECT 166.010 0.320 166.150 0.610 ;
        RECT 166.970 0.320 167.110 0.610 ;
        RECT 167.930 0.320 168.070 0.610 ;
        RECT 168.890 0.320 169.030 0.610 ;
        RECT 169.850 0.320 169.990 0.610 ;
        RECT 170.810 0.320 170.950 0.610 ;
        RECT 171.770 0.320 171.910 0.610 ;
        RECT 172.730 0.320 172.870 0.610 ;
        RECT 173.690 0.320 173.830 0.610 ;
        RECT 174.650 0.320 174.790 0.610 ;
        RECT 175.610 0.320 175.750 0.610 ;
        RECT 176.570 0.320 176.710 0.610 ;
        RECT 177.530 0.320 177.670 0.610 ;
        RECT 178.490 0.320 178.630 0.610 ;
        RECT 179.450 0.320 179.590 0.610 ;
        RECT 180.410 0.320 180.550 0.610 ;
        RECT 181.370 0.320 181.510 0.610 ;
        RECT 182.330 0.320 182.470 0.610 ;
        RECT 183.290 0.320 183.430 0.610 ;
        RECT 184.250 0.320 184.390 0.610 ;
        RECT 185.210 0.320 185.350 0.610 ;
        RECT 186.170 0.320 186.310 0.610 ;
        RECT 187.130 0.320 187.270 0.610 ;
        RECT 188.090 0.320 188.230 0.610 ;
        RECT 189.050 0.320 189.190 0.610 ;
        RECT 190.010 0.320 190.150 0.610 ;
        RECT 190.970 0.320 191.110 0.610 ;
        RECT 191.930 0.320 192.070 0.610 ;
        RECT 192.890 0.320 193.030 0.610 ;
        RECT 193.850 0.320 193.990 0.610 ;
        RECT 194.810 0.320 194.950 0.610 ;
        RECT 195.770 0.320 195.910 0.610 ;
        RECT 196.730 0.320 196.870 0.610 ;
        RECT 197.690 0.320 197.830 0.610 ;
        RECT 198.650 0.320 198.790 0.610 ;
        RECT 199.610 0.320 199.750 0.610 ;
        RECT 200.570 0.320 200.710 0.610 ;
        RECT 201.530 0.320 201.670 0.610 ;
        RECT 202.490 0.320 202.630 0.610 ;
        RECT 203.450 0.320 203.590 0.610 ;
        RECT 204.410 0.320 204.550 0.610 ;
        RECT 205.370 0.320 205.510 0.610 ;
        RECT 206.330 0.320 206.470 0.610 ;
        RECT 207.290 0.320 207.430 0.610 ;
        RECT 208.250 0.320 208.390 0.610 ;
        RECT 209.210 0.320 209.350 0.610 ;
        RECT 210.170 0.320 210.310 0.610 ;
        RECT 211.130 0.320 211.270 0.610 ;
        RECT 212.090 0.320 212.230 0.610 ;
        RECT 213.050 0.320 213.190 0.610 ;
        RECT 214.010 0.320 214.150 0.610 ;
        RECT 214.970 0.320 215.110 0.610 ;
        RECT 215.930 0.320 216.070 0.610 ;
        RECT 216.890 0.320 217.030 0.610 ;
        RECT 217.850 0.320 217.990 0.610 ;
        RECT 218.810 0.320 218.950 0.610 ;
        RECT 219.770 0.320 219.910 0.610 ;
        RECT 220.730 0.320 220.870 0.610 ;
        RECT 221.690 0.320 221.830 0.610 ;
        RECT 222.650 0.320 222.790 0.610 ;
        RECT 223.610 0.320 223.750 0.610 ;
        RECT 224.570 0.320 224.710 0.610 ;
        RECT 225.530 0.320 225.670 0.610 ;
        RECT 226.490 0.320 226.630 0.610 ;
        RECT 227.450 0.320 227.590 0.610 ;
        RECT 228.410 0.320 228.550 0.610 ;
        RECT 229.370 0.320 229.510 0.610 ;
        RECT 230.330 0.320 230.470 0.610 ;
        RECT 231.290 0.320 231.430 0.610 ;
        RECT 232.250 0.320 232.390 0.610 ;
        RECT 233.210 0.320 233.350 0.610 ;
        RECT 234.170 0.320 234.310 0.610 ;
        RECT 235.130 0.320 235.270 0.610 ;
        RECT 236.090 0.320 236.230 0.610 ;
        RECT 237.050 0.320 237.190 0.610 ;
        RECT 238.010 0.320 238.150 0.610 ;
        RECT 238.970 0.320 239.110 0.610 ;
        RECT 239.930 0.320 240.070 0.610 ;
        RECT 240.890 0.320 241.030 0.610 ;
        RECT 241.850 0.320 241.990 0.610 ;
        RECT 242.810 0.320 242.950 0.610 ;
        RECT 243.770 0.320 243.910 0.610 ;
        RECT 244.730 0.320 244.870 0.610 ;
        RECT 245.690 0.320 245.830 0.610 ;
        RECT 246.650 0.320 246.790 0.610 ;
        RECT 247.610 0.320 247.750 0.610 ;
        RECT 248.570 0.320 248.710 0.610 ;
        RECT 249.530 0.320 249.670 0.610 ;
        RECT 250.490 0.320 250.630 0.610 ;
        RECT 251.450 0.320 251.590 0.610 ;
        RECT 252.410 0.320 252.550 0.610 ;
        RECT 253.370 0.320 253.510 0.610 ;
        RECT 254.330 0.320 254.470 0.610 ;
        RECT 255.290 0.320 255.430 0.610 ;
        RECT 256.250 0.320 256.390 0.610 ;
        RECT 257.210 0.320 257.350 0.610 ;
        RECT 258.170 0.320 258.310 0.610 ;
        RECT 259.130 0.320 259.270 0.610 ;
        RECT 260.090 0.320 260.230 0.610 ;
        RECT 261.050 0.320 261.190 0.610 ;
        RECT 262.010 0.320 262.150 0.610 ;
        RECT 262.970 0.320 263.110 0.610 ;
        RECT 263.930 0.320 264.070 0.610 ;
        RECT 264.890 0.320 265.030 0.610 ;
        RECT 265.850 0.320 265.990 0.610 ;
        RECT 266.810 0.320 266.950 0.610 ;
        RECT 267.770 0.320 267.910 0.610 ;
        RECT 268.730 0.320 268.870 0.610 ;
        RECT 269.690 0.320 269.830 0.610 ;
        RECT 270.650 0.320 270.790 0.610 ;
        RECT 271.610 0.320 271.750 0.610 ;
        RECT 272.570 0.320 272.710 0.610 ;
        RECT 273.530 0.320 273.670 0.610 ;
        RECT 274.490 0.320 274.630 0.610 ;
        RECT 275.450 0.320 275.590 0.610 ;
        RECT 276.410 0.320 276.550 0.610 ;
        RECT 277.370 0.320 277.510 0.610 ;
        RECT 278.330 0.320 278.470 0.610 ;
        RECT 279.290 0.320 279.430 0.610 ;
        RECT 280.250 0.320 280.390 0.610 ;
        RECT 281.210 0.320 281.350 0.610 ;
        RECT 282.170 0.320 282.310 0.610 ;
        RECT 283.130 0.320 283.270 0.610 ;
        RECT 284.090 0.320 284.230 0.610 ;
        RECT 285.050 0.320 285.190 0.610 ;
        RECT 286.010 0.320 286.150 0.610 ;
        RECT 286.970 0.320 287.110 0.610 ;
        RECT 287.930 0.320 288.070 0.610 ;
        RECT 288.890 0.320 289.030 0.610 ;
        RECT 289.850 0.320 289.990 0.610 ;
        RECT 290.810 0.320 290.950 0.610 ;
        RECT 291.770 0.320 291.910 0.610 ;
        RECT 292.730 0.320 292.870 0.610 ;
        RECT 293.690 0.320 293.830 0.610 ;
        RECT 294.650 0.320 294.790 0.610 ;
        RECT 295.610 0.320 295.750 0.610 ;
        RECT 296.570 0.320 296.710 0.610 ;
        RECT 297.530 0.320 297.670 0.610 ;
        RECT 298.490 0.320 298.630 0.610 ;
        RECT 299.450 0.320 299.590 0.610 ;
        RECT 300.410 0.320 300.550 0.610 ;
        RECT 301.370 0.320 301.510 0.610 ;
        RECT 302.330 0.320 302.470 0.610 ;
        RECT 303.290 0.320 303.430 0.610 ;
        RECT 304.250 0.320 304.390 0.610 ;
        RECT 305.210 0.320 305.350 0.610 ;
        RECT 306.170 0.320 306.310 0.610 ;
        RECT 307.130 0.320 307.270 0.610 ;
        RECT 308.090 0.320 308.230 0.610 ;
        RECT 309.050 0.320 309.190 0.610 ;
        RECT 310.010 0.320 310.150 0.610 ;
        RECT 310.970 0.320 311.110 0.610 ;
        RECT 311.930 0.320 312.070 0.610 ;
        RECT 312.890 0.320 313.030 0.610 ;
        RECT 313.850 0.320 313.990 0.610 ;
        RECT 314.810 0.320 314.950 0.610 ;
        RECT 315.770 0.320 315.910 0.610 ;
        RECT 316.730 0.320 316.870 0.610 ;
        RECT 317.690 0.320 317.830 0.610 ;
        RECT 318.650 0.320 318.790 0.610 ;
        RECT 319.610 0.320 319.750 0.610 ;
        RECT 320.570 0.320 320.710 0.610 ;
        RECT 321.530 0.320 321.670 0.610 ;
        RECT 322.490 0.320 322.630 0.610 ;
        RECT 323.450 0.320 323.590 0.610 ;
        RECT 324.410 0.320 324.550 0.610 ;
        RECT 325.370 0.320 325.510 0.610 ;
        RECT 326.330 0.320 326.470 0.610 ;
        RECT 327.290 0.320 327.430 0.610 ;
        RECT 328.250 0.320 328.390 0.610 ;
        RECT 329.210 0.320 329.350 0.610 ;
        RECT 330.170 0.320 330.310 0.610 ;
        RECT 331.130 0.320 331.270 0.610 ;
        RECT 332.090 0.320 332.230 0.610 ;
        RECT 333.050 0.320 333.190 0.610 ;
        RECT 334.010 0.320 334.150 0.610 ;
        RECT 334.970 0.320 335.110 0.610 ;
        RECT 335.930 0.320 336.070 0.610 ;
        RECT 336.890 0.320 337.030 0.610 ;
        RECT 337.850 0.320 337.990 0.610 ;
        RECT 338.810 0.320 338.950 0.610 ;
        RECT 339.770 0.320 339.910 0.610 ;
        RECT 340.730 0.320 340.870 0.610 ;
        RECT 341.690 0.320 341.830 0.610 ;
        RECT 342.650 0.320 342.790 0.610 ;
        RECT 343.610 0.320 343.750 0.610 ;
        RECT 344.570 0.320 344.710 0.610 ;
        RECT 345.530 0.320 345.670 0.610 ;
        RECT 346.490 0.320 346.630 0.610 ;
        RECT 347.450 0.320 347.590 0.610 ;
        RECT 348.410 0.320 348.550 0.610 ;
        RECT 349.370 0.320 349.510 0.610 ;
        RECT 350.330 0.320 350.470 0.610 ;
        RECT 351.290 0.320 351.430 0.610 ;
        RECT 352.250 0.320 352.390 0.610 ;
        RECT 353.210 0.320 353.350 0.610 ;
        RECT 354.170 0.320 354.310 0.610 ;
        RECT 355.130 0.320 355.270 0.610 ;
        RECT 356.090 0.320 356.230 0.610 ;
        RECT 357.050 0.320 357.190 0.610 ;
        RECT 358.010 0.320 358.150 0.610 ;
        RECT 358.970 0.320 359.110 0.610 ;
        RECT 359.930 0.320 360.070 0.610 ;
        RECT 360.890 0.320 361.030 0.610 ;
        RECT 361.850 0.320 361.990 0.610 ;
        RECT 362.810 0.320 362.950 0.610 ;
        RECT 363.770 0.320 363.910 0.610 ;
        RECT 364.730 0.320 364.870 0.610 ;
        RECT 365.690 0.320 365.830 0.610 ;
        RECT 366.650 0.320 366.790 0.610 ;
        RECT 367.610 0.320 367.750 0.610 ;
        RECT 368.570 0.320 368.710 0.610 ;
        RECT 369.530 0.320 369.670 0.610 ;
        RECT 370.490 0.320 370.630 0.610 ;
        RECT 371.450 0.320 371.590 0.610 ;
        RECT 372.410 0.320 372.550 0.610 ;
        RECT 373.370 0.320 373.510 0.610 ;
        RECT 374.330 0.320 374.470 0.610 ;
        RECT 375.290 0.320 375.430 0.610 ;
        RECT 376.250 0.320 376.390 0.610 ;
        RECT 377.210 0.320 377.350 0.610 ;
        RECT 378.170 0.320 378.310 0.610 ;
        RECT 379.130 0.320 379.270 0.610 ;
        RECT 380.090 0.320 380.230 0.610 ;
        RECT 381.050 0.320 381.190 0.610 ;
        RECT 382.010 0.320 382.150 0.610 ;
        RECT 382.970 0.320 383.110 0.610 ;
        RECT 383.930 0.320 384.070 0.610 ;
        RECT 384.890 0.320 385.030 0.610 ;
        RECT 385.850 0.320 385.990 0.610 ;
        RECT 386.810 0.320 386.950 0.610 ;
        RECT 387.770 0.320 387.910 0.610 ;
        RECT 388.730 0.320 388.870 0.610 ;
        RECT 389.690 0.320 389.830 0.610 ;
        RECT 390.650 0.320 390.790 0.610 ;
        RECT 391.610 0.320 391.750 0.610 ;
        RECT 392.570 0.320 392.710 0.610 ;
        RECT 393.530 0.320 393.670 0.610 ;
        RECT 394.490 0.320 394.630 0.610 ;
        RECT 395.450 0.320 395.590 0.610 ;
        RECT 396.410 0.320 396.550 0.610 ;
        RECT 397.370 0.320 397.510 0.610 ;
        RECT 398.330 0.320 398.470 0.610 ;
        RECT 399.290 0.320 399.430 0.610 ;
        RECT 400.250 0.320 400.390 0.610 ;
        RECT 401.210 0.320 401.350 0.610 ;
        RECT 402.170 0.320 402.310 0.610 ;
        RECT 403.130 0.320 403.270 0.610 ;
        RECT 404.090 0.320 404.230 0.610 ;
        RECT 405.050 0.320 405.190 0.610 ;
        RECT 406.010 0.320 406.150 0.610 ;
        RECT 406.970 0.320 407.110 0.610 ;
        RECT 407.930 0.320 408.070 0.610 ;
        RECT 408.890 0.320 409.030 0.610 ;
        RECT 409.850 0.320 409.990 0.610 ;
        RECT 410.810 0.320 410.950 0.610 ;
        RECT 411.770 0.320 411.910 0.610 ;
        RECT 412.730 0.320 412.870 0.610 ;
        RECT 413.690 0.320 413.830 0.610 ;
        RECT 414.650 0.320 414.790 0.610 ;
        RECT 415.610 0.320 415.750 0.610 ;
        RECT 416.570 0.320 416.710 0.610 ;
        RECT 417.530 0.320 417.670 0.610 ;
        RECT 418.490 0.320 418.630 0.610 ;
        RECT 419.450 0.320 419.590 0.610 ;
        RECT 420.410 0.320 420.550 0.610 ;
        RECT 421.370 0.320 421.510 0.610 ;
        RECT 422.330 0.320 422.470 0.610 ;
        RECT 423.290 0.320 423.430 0.610 ;
        RECT 424.250 0.320 424.390 0.610 ;
        RECT 425.210 0.320 425.350 0.610 ;
        RECT 426.170 0.320 426.310 0.610 ;
        RECT 427.130 0.320 427.270 0.610 ;
        RECT 428.090 0.320 428.230 0.610 ;
        RECT 429.050 0.320 429.190 0.610 ;
        RECT 430.010 0.320 430.150 0.610 ;
        RECT 430.970 0.320 431.110 0.610 ;
        RECT 431.930 0.320 432.070 0.610 ;
        RECT 432.890 0.320 433.030 0.610 ;
        RECT 433.850 0.320 433.990 0.610 ;
        RECT 434.810 0.320 434.950 0.610 ;
        RECT 435.770 0.320 435.910 0.610 ;
        RECT 436.730 0.320 436.870 0.610 ;
        RECT 437.690 0.320 437.830 0.610 ;
        RECT 438.650 0.320 438.790 0.610 ;
        RECT 439.610 0.320 439.750 0.610 ;
        RECT 440.570 0.320 440.710 0.610 ;
        RECT 441.530 0.320 441.670 0.610 ;
        RECT 442.490 0.320 442.630 0.610 ;
        RECT 443.450 0.320 443.590 0.610 ;
        RECT 444.410 0.320 444.550 0.610 ;
        RECT 445.370 0.320 445.510 0.610 ;
        RECT 446.330 0.320 446.470 0.610 ;
        RECT 447.290 0.320 447.430 0.610 ;
        RECT 448.250 0.320 448.390 0.610 ;
        RECT 449.210 0.320 449.350 0.610 ;
        RECT 450.170 0.320 450.310 0.610 ;
        RECT 451.130 0.320 451.270 0.610 ;
        RECT 452.090 0.320 452.230 0.610 ;
        RECT 453.050 0.320 453.190 0.610 ;
        RECT 454.010 0.320 454.150 0.610 ;
        RECT 454.970 0.320 455.110 0.610 ;
        RECT 455.930 0.320 456.070 0.610 ;
        RECT 456.890 0.320 457.030 0.610 ;
        RECT 457.850 0.320 457.990 0.610 ;
        RECT 458.810 0.320 458.950 0.610 ;
        RECT 459.770 0.320 459.910 0.610 ;
        RECT 460.730 0.320 460.870 0.610 ;
        RECT 461.690 0.320 461.830 0.610 ;
        RECT 462.650 0.320 462.790 0.610 ;
        RECT 463.610 0.320 463.750 0.610 ;
        RECT 464.570 0.320 464.710 0.610 ;
        RECT 465.530 0.320 465.670 0.610 ;
        RECT 466.490 0.320 466.630 0.610 ;
        RECT 467.450 0.320 467.590 0.610 ;
        RECT 468.410 0.320 468.550 0.610 ;
        RECT 469.370 0.320 469.510 0.610 ;
        RECT 470.330 0.320 470.470 0.610 ;
        RECT 471.290 0.320 471.430 0.610 ;
        RECT 472.250 0.320 472.390 0.610 ;
        RECT 473.210 0.320 473.350 0.610 ;
        RECT 474.170 0.320 474.310 0.610 ;
        RECT 475.130 0.320 475.270 0.610 ;
        RECT 476.090 0.320 476.230 0.610 ;
        RECT 477.050 0.320 477.190 0.610 ;
        RECT 478.010 0.320 478.150 0.610 ;
        RECT 478.970 0.320 479.110 0.610 ;
        RECT 479.930 0.320 480.070 0.610 ;
        RECT 480.890 0.320 481.030 0.610 ;
        RECT 481.850 0.320 481.990 0.610 ;
        RECT 482.810 0.320 482.950 0.610 ;
        RECT 483.770 0.320 483.910 0.610 ;
        RECT 484.730 0.320 484.870 0.610 ;
        RECT 485.690 0.320 485.830 0.610 ;
        RECT 486.650 0.320 486.790 0.610 ;
        RECT 487.610 0.320 487.750 0.610 ;
        RECT 488.570 0.320 488.710 0.610 ;
        RECT 489.530 0.320 489.670 0.610 ;
        RECT 490.490 0.320 490.630 0.610 ;
        RECT 491.450 0.320 491.590 0.610 ;
        RECT 492.410 0.320 492.550 0.610 ;
        RECT 493.370 0.320 493.510 0.610 ;
        RECT 494.330 0.320 494.470 0.610 ;
      LAYER Metal3 ;
        RECT 5.135 0.320 495.025 59.740 ;
      LAYER Metal4 ;
        RECT 6.135 0.695 490.665 56.845 ;
      LAYER Metal5 ;
        RECT 6.095 14.810 490.705 57.010 ;
      LAYER TopMetal1 ;
        RECT 7.530 16.400 16.620 23.080 ;
        RECT 22.100 16.400 22.820 23.080 ;
        RECT 28.300 16.400 92.220 23.080 ;
        RECT 97.700 16.400 98.420 23.080 ;
        RECT 103.900 16.400 166.750 23.080 ;
      LAYER TopMetal2 ;
        RECT 7.480 17.000 166.800 23.000 ;
  END
END decoder
END LIBRARY

