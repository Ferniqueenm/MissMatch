magic
tech ihp-sg13g2
magscale 1 2
timestamp 1752134018
<< metal1 >>
rect 1152 11360 98784 11384
rect 1152 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 33928 11360
rect 33968 11320 34010 11360
rect 34050 11320 34092 11360
rect 34132 11320 34174 11360
rect 34214 11320 34256 11360
rect 34296 11320 49048 11360
rect 49088 11320 49130 11360
rect 49170 11320 49212 11360
rect 49252 11320 49294 11360
rect 49334 11320 49376 11360
rect 49416 11320 64168 11360
rect 64208 11320 64250 11360
rect 64290 11320 64332 11360
rect 64372 11320 64414 11360
rect 64454 11320 64496 11360
rect 64536 11320 79288 11360
rect 79328 11320 79370 11360
rect 79410 11320 79452 11360
rect 79492 11320 79534 11360
rect 79574 11320 79616 11360
rect 79656 11320 94408 11360
rect 94448 11320 94490 11360
rect 94530 11320 94572 11360
rect 94612 11320 94654 11360
rect 94694 11320 94736 11360
rect 94776 11320 98784 11360
rect 1152 11296 98784 11320
rect 11883 11192 11925 11201
rect 11883 11152 11884 11192
rect 11924 11152 11925 11192
rect 11883 11143 11925 11152
rect 30891 11192 30933 11201
rect 30891 11152 30892 11192
rect 30932 11152 30933 11192
rect 30891 11143 30933 11152
rect 19563 11108 19605 11117
rect 19563 11068 19564 11108
rect 19604 11068 19605 11108
rect 19563 11059 19605 11068
rect 50083 11024 50141 11025
rect 50083 10984 50092 11024
rect 50132 10984 50141 11024
rect 50083 10983 50141 10984
rect 11787 10940 11829 10949
rect 11787 10900 11788 10940
rect 11828 10900 11829 10940
rect 11787 10891 11829 10900
rect 11971 10940 12029 10941
rect 11971 10900 11980 10940
rect 12020 10900 12029 10940
rect 11971 10899 12029 10900
rect 12163 10940 12221 10941
rect 12163 10900 12172 10940
rect 12212 10900 12221 10940
rect 12163 10899 12221 10900
rect 12363 10940 12405 10949
rect 12363 10900 12364 10940
rect 12404 10900 12405 10940
rect 12363 10891 12405 10900
rect 15627 10940 15669 10949
rect 15627 10900 15628 10940
rect 15668 10900 15669 10940
rect 15627 10891 15669 10900
rect 15811 10940 15869 10941
rect 15811 10900 15820 10940
rect 15860 10900 15869 10940
rect 15811 10899 15869 10900
rect 17251 10940 17309 10941
rect 17251 10900 17260 10940
rect 17300 10900 17309 10940
rect 17251 10899 17309 10900
rect 17443 10940 17501 10941
rect 17443 10900 17452 10940
rect 17492 10900 17501 10940
rect 17443 10899 17501 10900
rect 19467 10940 19509 10949
rect 19467 10900 19468 10940
rect 19508 10900 19509 10940
rect 19467 10891 19509 10900
rect 19651 10940 19709 10941
rect 19651 10900 19660 10940
rect 19700 10900 19709 10940
rect 19651 10899 19709 10900
rect 24171 10940 24213 10949
rect 24171 10900 24172 10940
rect 24212 10900 24213 10940
rect 24171 10891 24213 10900
rect 24355 10940 24413 10941
rect 24355 10900 24364 10940
rect 24404 10900 24413 10940
rect 24355 10899 24413 10900
rect 24555 10940 24597 10949
rect 24555 10900 24556 10940
rect 24596 10900 24597 10940
rect 24555 10891 24597 10900
rect 24739 10940 24797 10941
rect 24739 10900 24748 10940
rect 24788 10900 24797 10940
rect 24739 10899 24797 10900
rect 24939 10940 24981 10949
rect 24939 10900 24940 10940
rect 24980 10900 24981 10940
rect 24939 10891 24981 10900
rect 25123 10940 25181 10941
rect 25123 10900 25132 10940
rect 25172 10900 25181 10940
rect 25123 10899 25181 10900
rect 28195 10940 28253 10941
rect 28195 10900 28204 10940
rect 28244 10900 28253 10940
rect 28195 10899 28253 10900
rect 28387 10940 28445 10941
rect 28387 10900 28396 10940
rect 28436 10900 28445 10940
rect 28387 10899 28445 10900
rect 30795 10940 30837 10949
rect 30795 10900 30796 10940
rect 30836 10900 30837 10940
rect 30795 10891 30837 10900
rect 30979 10940 31037 10941
rect 30979 10900 30988 10940
rect 31028 10900 31037 10940
rect 30979 10899 31037 10900
rect 31179 10940 31221 10949
rect 31179 10900 31180 10940
rect 31220 10900 31221 10940
rect 31179 10891 31221 10900
rect 31363 10940 31421 10941
rect 31363 10900 31372 10940
rect 31412 10900 31421 10940
rect 31363 10899 31421 10900
rect 36459 10940 36501 10949
rect 36459 10900 36460 10940
rect 36500 10900 36501 10940
rect 36459 10891 36501 10900
rect 36643 10940 36701 10941
rect 36643 10900 36652 10940
rect 36692 10900 36701 10940
rect 36643 10899 36701 10900
rect 36843 10940 36885 10949
rect 36843 10900 36844 10940
rect 36884 10900 36885 10940
rect 36843 10891 36885 10900
rect 37027 10940 37085 10941
rect 37027 10900 37036 10940
rect 37076 10900 37085 10940
rect 37027 10899 37085 10900
rect 39139 10940 39197 10941
rect 39139 10900 39148 10940
rect 39188 10900 39197 10940
rect 39139 10899 39197 10900
rect 39331 10940 39389 10941
rect 39331 10900 39340 10940
rect 39380 10900 39389 10940
rect 39331 10899 39389 10900
rect 61027 10940 61085 10941
rect 61027 10900 61036 10940
rect 61076 10900 61085 10940
rect 61027 10899 61085 10900
rect 61219 10940 61277 10941
rect 61219 10900 61228 10940
rect 61268 10900 61277 10940
rect 61219 10899 61277 10900
rect 71971 10940 72029 10941
rect 71971 10900 71980 10940
rect 72020 10900 72029 10940
rect 71971 10899 72029 10900
rect 72163 10940 72221 10941
rect 72163 10900 72172 10940
rect 72212 10900 72221 10940
rect 72163 10899 72221 10900
rect 82915 10940 82973 10941
rect 82915 10900 82924 10940
rect 82964 10900 82973 10940
rect 82915 10899 82973 10900
rect 83107 10940 83165 10941
rect 83107 10900 83116 10940
rect 83156 10900 83165 10940
rect 83107 10899 83165 10900
rect 12267 10856 12309 10865
rect 12267 10816 12268 10856
rect 12308 10816 12309 10856
rect 12267 10807 12309 10816
rect 15723 10856 15765 10865
rect 15723 10816 15724 10856
rect 15764 10816 15765 10856
rect 15723 10807 15765 10816
rect 24267 10856 24309 10865
rect 24267 10816 24268 10856
rect 24308 10816 24309 10856
rect 24267 10807 24309 10816
rect 24651 10856 24693 10865
rect 24651 10816 24652 10856
rect 24692 10816 24693 10856
rect 24651 10807 24693 10816
rect 25035 10856 25077 10865
rect 25035 10816 25036 10856
rect 25076 10816 25077 10856
rect 25035 10807 25077 10816
rect 31275 10856 31317 10865
rect 31275 10816 31276 10856
rect 31316 10816 31317 10856
rect 31275 10807 31317 10816
rect 36555 10856 36597 10865
rect 36555 10816 36556 10856
rect 36596 10816 36597 10856
rect 36555 10807 36597 10816
rect 36939 10856 36981 10865
rect 36939 10816 36940 10856
rect 36980 10816 36981 10856
rect 36939 10807 36981 10816
rect 50283 10772 50325 10781
rect 50283 10732 50284 10772
rect 50324 10732 50325 10772
rect 50283 10723 50325 10732
rect 1152 10604 98784 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 65408 10604
rect 65448 10564 65490 10604
rect 65530 10564 65572 10604
rect 65612 10564 65654 10604
rect 65694 10564 65736 10604
rect 65776 10564 80528 10604
rect 80568 10564 80610 10604
rect 80650 10564 80692 10604
rect 80732 10564 80774 10604
rect 80814 10564 80856 10604
rect 80896 10564 95648 10604
rect 95688 10564 95730 10604
rect 95770 10564 95812 10604
rect 95852 10564 95894 10604
rect 95934 10564 95976 10604
rect 96016 10564 98784 10604
rect 1152 10540 98784 10564
rect 57675 10436 57717 10445
rect 57675 10396 57676 10436
rect 57716 10396 57717 10436
rect 57675 10387 57717 10396
rect 10923 10352 10965 10361
rect 10923 10312 10924 10352
rect 10964 10312 10965 10352
rect 10923 10303 10965 10312
rect 19083 10352 19125 10361
rect 19083 10312 19084 10352
rect 19124 10312 19125 10352
rect 19083 10303 19125 10312
rect 19851 10352 19893 10361
rect 19851 10312 19852 10352
rect 19892 10312 19893 10352
rect 19851 10303 19893 10312
rect 23883 10352 23925 10361
rect 23883 10312 23884 10352
rect 23924 10312 23925 10352
rect 23883 10303 23925 10312
rect 36075 10352 36117 10361
rect 36075 10312 36076 10352
rect 36116 10312 36117 10352
rect 36075 10303 36117 10312
rect 36459 10352 36501 10361
rect 36459 10312 36460 10352
rect 36500 10312 36501 10352
rect 36459 10303 36501 10312
rect 49411 10352 49469 10353
rect 49411 10312 49420 10352
rect 49460 10312 49469 10352
rect 49411 10311 49469 10312
rect 84075 10352 84117 10361
rect 84075 10312 84076 10352
rect 84116 10312 84117 10352
rect 84075 10303 84117 10312
rect 88299 10352 88341 10361
rect 88299 10312 88300 10352
rect 88340 10312 88341 10352
rect 88299 10303 88341 10312
rect 12355 10289 12413 10290
rect 10827 10268 10869 10277
rect 10827 10228 10828 10268
rect 10868 10228 10869 10268
rect 10827 10219 10869 10228
rect 11011 10268 11069 10269
rect 11011 10228 11020 10268
rect 11060 10228 11069 10268
rect 11011 10227 11069 10228
rect 11203 10268 11261 10269
rect 11203 10228 11212 10268
rect 11252 10228 11261 10268
rect 11203 10227 11261 10228
rect 11403 10268 11445 10277
rect 11403 10228 11404 10268
rect 11444 10228 11445 10268
rect 11403 10219 11445 10228
rect 11595 10268 11637 10277
rect 11595 10228 11596 10268
rect 11636 10228 11637 10268
rect 11595 10219 11637 10228
rect 11779 10268 11837 10269
rect 11779 10228 11788 10268
rect 11828 10228 11837 10268
rect 11779 10227 11837 10228
rect 11971 10268 12029 10269
rect 11971 10228 11980 10268
rect 12020 10228 12029 10268
rect 11971 10227 12029 10228
rect 12171 10268 12213 10277
rect 12171 10228 12172 10268
rect 12212 10228 12213 10268
rect 12355 10249 12364 10289
rect 12404 10249 12413 10289
rect 24355 10289 24413 10290
rect 12355 10248 12413 10249
rect 12555 10268 12597 10277
rect 12171 10219 12213 10228
rect 12555 10228 12556 10268
rect 12596 10228 12597 10268
rect 12555 10219 12597 10228
rect 12739 10268 12797 10269
rect 12739 10228 12748 10268
rect 12788 10228 12797 10268
rect 12739 10227 12797 10228
rect 12939 10268 12981 10277
rect 12939 10228 12940 10268
rect 12980 10228 12981 10268
rect 12939 10219 12981 10228
rect 14571 10268 14613 10277
rect 14571 10228 14572 10268
rect 14612 10228 14613 10268
rect 14571 10219 14613 10228
rect 14755 10268 14813 10269
rect 14755 10228 14764 10268
rect 14804 10228 14813 10268
rect 14755 10227 14813 10228
rect 14955 10268 14997 10277
rect 14955 10228 14956 10268
rect 14996 10228 14997 10268
rect 14955 10219 14997 10228
rect 15139 10268 15197 10269
rect 15139 10228 15148 10268
rect 15188 10228 15197 10268
rect 15139 10227 15197 10228
rect 15339 10268 15381 10277
rect 15339 10228 15340 10268
rect 15380 10228 15381 10268
rect 15339 10219 15381 10228
rect 15523 10268 15581 10269
rect 15523 10228 15532 10268
rect 15572 10228 15581 10268
rect 15523 10227 15581 10228
rect 15723 10268 15765 10277
rect 15723 10228 15724 10268
rect 15764 10228 15765 10268
rect 15723 10219 15765 10228
rect 15907 10268 15965 10269
rect 15907 10228 15916 10268
rect 15956 10228 15965 10268
rect 15907 10227 15965 10228
rect 16099 10268 16157 10269
rect 16099 10228 16108 10268
rect 16148 10228 16157 10268
rect 16099 10227 16157 10228
rect 16299 10268 16341 10277
rect 16299 10228 16300 10268
rect 16340 10228 16341 10268
rect 16299 10219 16341 10228
rect 18595 10268 18653 10269
rect 18595 10228 18604 10268
rect 18644 10228 18653 10268
rect 18595 10227 18653 10228
rect 18795 10268 18837 10277
rect 18795 10228 18796 10268
rect 18836 10228 18837 10268
rect 18795 10219 18837 10228
rect 18987 10268 19029 10277
rect 18987 10228 18988 10268
rect 19028 10228 19029 10268
rect 18987 10219 19029 10228
rect 19171 10268 19229 10269
rect 19171 10228 19180 10268
rect 19220 10228 19229 10268
rect 19171 10227 19229 10228
rect 19371 10268 19413 10277
rect 19371 10228 19372 10268
rect 19412 10228 19413 10268
rect 19371 10219 19413 10228
rect 19555 10268 19613 10269
rect 19555 10228 19564 10268
rect 19604 10228 19613 10268
rect 19555 10227 19613 10228
rect 19755 10268 19797 10277
rect 19755 10228 19756 10268
rect 19796 10228 19797 10268
rect 19755 10219 19797 10228
rect 19939 10268 19997 10269
rect 19939 10228 19948 10268
rect 19988 10228 19997 10268
rect 20323 10268 20381 10269
rect 19939 10227 19997 10228
rect 20130 10253 20172 10262
rect 20130 10213 20131 10253
rect 20171 10213 20172 10253
rect 20323 10228 20332 10268
rect 20372 10228 20381 10268
rect 20323 10227 20381 10228
rect 21675 10268 21717 10277
rect 21675 10228 21676 10268
rect 21716 10228 21717 10268
rect 21675 10219 21717 10228
rect 23779 10268 23837 10269
rect 23779 10228 23788 10268
rect 23828 10228 23837 10268
rect 23779 10227 23837 10228
rect 23979 10268 24021 10277
rect 23979 10228 23980 10268
rect 24020 10228 24021 10268
rect 23979 10219 24021 10228
rect 24171 10268 24213 10277
rect 24171 10228 24172 10268
rect 24212 10228 24213 10268
rect 24355 10249 24364 10289
rect 24404 10249 24413 10289
rect 31171 10289 31229 10290
rect 24355 10248 24413 10249
rect 24555 10268 24597 10277
rect 24171 10219 24213 10228
rect 24555 10228 24556 10268
rect 24596 10228 24597 10268
rect 24555 10219 24597 10228
rect 24739 10268 24797 10269
rect 24739 10228 24748 10268
rect 24788 10228 24797 10268
rect 24739 10227 24797 10228
rect 25419 10268 25461 10277
rect 25419 10228 25420 10268
rect 25460 10228 25461 10268
rect 25419 10219 25461 10228
rect 30219 10268 30261 10277
rect 30219 10228 30220 10268
rect 30260 10228 30261 10268
rect 30219 10219 30261 10228
rect 30403 10268 30461 10269
rect 30403 10228 30412 10268
rect 30452 10228 30461 10268
rect 30403 10227 30461 10228
rect 30603 10268 30645 10277
rect 30603 10228 30604 10268
rect 30644 10228 30645 10268
rect 30603 10219 30645 10228
rect 30787 10268 30845 10269
rect 30787 10228 30796 10268
rect 30836 10228 30845 10268
rect 30787 10227 30845 10228
rect 30987 10268 31029 10277
rect 30987 10228 30988 10268
rect 31028 10228 31029 10268
rect 31171 10249 31180 10289
rect 31220 10249 31229 10289
rect 31171 10248 31229 10249
rect 31371 10268 31413 10277
rect 30987 10219 31029 10228
rect 31371 10228 31372 10268
rect 31412 10228 31413 10268
rect 31371 10219 31413 10228
rect 31555 10268 31613 10269
rect 31555 10228 31564 10268
rect 31604 10228 31613 10268
rect 31555 10227 31613 10228
rect 32043 10268 32085 10277
rect 32043 10228 32044 10268
rect 32084 10228 32085 10268
rect 32043 10219 32085 10228
rect 35587 10268 35645 10269
rect 35587 10228 35596 10268
rect 35636 10228 35645 10268
rect 35587 10227 35645 10228
rect 35787 10268 35829 10277
rect 35787 10228 35788 10268
rect 35828 10228 35829 10268
rect 35787 10219 35829 10228
rect 35979 10268 36021 10277
rect 35979 10228 35980 10268
rect 36020 10228 36021 10268
rect 35979 10219 36021 10228
rect 36163 10268 36221 10269
rect 36163 10228 36172 10268
rect 36212 10228 36221 10268
rect 36163 10227 36221 10228
rect 36363 10268 36405 10277
rect 36363 10228 36364 10268
rect 36404 10228 36405 10268
rect 36363 10219 36405 10228
rect 36547 10268 36605 10269
rect 36547 10228 36556 10268
rect 36596 10228 36605 10268
rect 36547 10227 36605 10228
rect 36747 10268 36789 10277
rect 36747 10228 36748 10268
rect 36788 10228 36789 10268
rect 36747 10219 36789 10228
rect 36931 10268 36989 10269
rect 36931 10228 36940 10268
rect 36980 10228 36989 10268
rect 36931 10227 36989 10228
rect 37411 10268 37469 10269
rect 37411 10228 37420 10268
rect 37460 10228 37469 10268
rect 37411 10227 37469 10228
rect 37611 10268 37653 10277
rect 37611 10228 37612 10268
rect 37652 10228 37653 10268
rect 37611 10219 37653 10228
rect 37803 10268 37845 10277
rect 37803 10228 37804 10268
rect 37844 10228 37845 10268
rect 37803 10219 37845 10228
rect 37987 10268 38045 10269
rect 37987 10228 37996 10268
rect 38036 10228 38045 10268
rect 37987 10227 38045 10228
rect 38187 10268 38229 10277
rect 38187 10228 38188 10268
rect 38228 10228 38229 10268
rect 38187 10219 38229 10228
rect 38371 10268 38429 10269
rect 38371 10228 38380 10268
rect 38420 10228 38429 10268
rect 38371 10227 38429 10228
rect 38571 10268 38613 10277
rect 38571 10228 38572 10268
rect 38612 10228 38613 10268
rect 38571 10219 38613 10228
rect 38755 10268 38813 10269
rect 38755 10228 38764 10268
rect 38804 10228 38813 10268
rect 38755 10227 38813 10228
rect 38955 10268 38997 10277
rect 38955 10228 38956 10268
rect 38996 10228 38997 10268
rect 38955 10219 38997 10228
rect 39139 10268 39197 10269
rect 39139 10228 39148 10268
rect 39188 10228 39197 10268
rect 39139 10227 39197 10228
rect 40579 10268 40637 10269
rect 40579 10228 40588 10268
rect 40628 10228 40637 10268
rect 40579 10227 40637 10228
rect 41539 10268 41597 10269
rect 41539 10228 41548 10268
rect 41588 10228 41597 10268
rect 41539 10227 41597 10228
rect 41827 10268 41885 10269
rect 41827 10228 41836 10268
rect 41876 10228 41885 10268
rect 41827 10227 41885 10228
rect 42787 10268 42845 10269
rect 42787 10228 42796 10268
rect 42836 10228 42845 10268
rect 42787 10227 42845 10228
rect 50275 10268 50333 10269
rect 50275 10228 50284 10268
rect 50324 10228 50333 10268
rect 50275 10227 50333 10228
rect 52099 10268 52157 10269
rect 52099 10228 52108 10268
rect 52148 10228 52157 10268
rect 52099 10227 52157 10228
rect 53059 10268 53117 10269
rect 53059 10228 53068 10268
rect 53108 10228 53117 10268
rect 53059 10227 53117 10228
rect 57579 10268 57621 10277
rect 57579 10228 57580 10268
rect 57620 10228 57621 10268
rect 57579 10219 57621 10228
rect 57771 10268 57813 10277
rect 57771 10228 57772 10268
rect 57812 10228 57813 10268
rect 57771 10219 57813 10228
rect 58155 10268 58197 10277
rect 58155 10228 58156 10268
rect 58196 10228 58197 10268
rect 58155 10219 58197 10228
rect 58617 10268 58659 10277
rect 58617 10228 58618 10268
rect 58658 10228 58659 10268
rect 58617 10219 58659 10228
rect 58923 10268 58965 10277
rect 58923 10228 58924 10268
rect 58964 10228 58965 10268
rect 58923 10219 58965 10228
rect 59115 10268 59157 10277
rect 59115 10228 59116 10268
rect 59156 10228 59157 10268
rect 59115 10219 59157 10228
rect 59883 10268 59925 10277
rect 59883 10228 59884 10268
rect 59924 10228 59925 10268
rect 59883 10219 59925 10228
rect 60075 10268 60117 10277
rect 60075 10228 60076 10268
rect 60116 10228 60117 10268
rect 60075 10219 60117 10228
rect 60267 10268 60309 10277
rect 60267 10228 60268 10268
rect 60308 10228 60309 10268
rect 60267 10219 60309 10228
rect 60459 10268 60501 10277
rect 60459 10228 60460 10268
rect 60500 10228 60501 10268
rect 60459 10219 60501 10228
rect 68419 10268 68477 10269
rect 68419 10228 68428 10268
rect 68468 10228 68477 10268
rect 68419 10227 68477 10228
rect 69571 10268 69629 10269
rect 69571 10228 69580 10268
rect 69620 10228 69629 10268
rect 69571 10227 69629 10228
rect 69763 10268 69821 10269
rect 69763 10228 69772 10268
rect 69812 10228 69821 10268
rect 69763 10227 69821 10228
rect 71307 10268 71349 10277
rect 71307 10228 71308 10268
rect 71348 10228 71349 10268
rect 71307 10219 71349 10228
rect 71491 10268 71549 10269
rect 71491 10228 71500 10268
rect 71540 10228 71549 10268
rect 71491 10227 71549 10228
rect 72931 10268 72989 10269
rect 72931 10228 72940 10268
rect 72980 10228 72989 10268
rect 72931 10227 72989 10228
rect 73131 10268 73173 10277
rect 73131 10228 73132 10268
rect 73172 10228 73173 10268
rect 73131 10219 73173 10228
rect 73315 10268 73373 10269
rect 73315 10228 73324 10268
rect 73364 10228 73373 10268
rect 73315 10227 73373 10228
rect 73507 10268 73565 10269
rect 73507 10228 73516 10268
rect 73556 10228 73565 10268
rect 73507 10227 73565 10228
rect 73795 10268 73853 10269
rect 73795 10228 73804 10268
rect 73844 10228 73853 10268
rect 73795 10227 73853 10228
rect 73987 10268 74045 10269
rect 73987 10228 73996 10268
rect 74036 10228 74045 10268
rect 73987 10227 74045 10228
rect 74275 10268 74333 10269
rect 74275 10228 74284 10268
rect 74324 10228 74333 10268
rect 74275 10227 74333 10228
rect 74475 10268 74517 10277
rect 74475 10228 74476 10268
rect 74516 10228 74517 10268
rect 74475 10219 74517 10228
rect 76483 10268 76541 10269
rect 76483 10228 76492 10268
rect 76532 10228 76541 10268
rect 76483 10227 76541 10228
rect 76683 10268 76725 10277
rect 76683 10228 76684 10268
rect 76724 10228 76725 10268
rect 76683 10219 76725 10228
rect 76875 10268 76917 10277
rect 76875 10228 76876 10268
rect 76916 10228 76917 10268
rect 76875 10219 76917 10228
rect 77059 10268 77117 10269
rect 77059 10228 77068 10268
rect 77108 10228 77117 10268
rect 77059 10227 77117 10228
rect 77251 10268 77309 10269
rect 77251 10228 77260 10268
rect 77300 10228 77309 10268
rect 77251 10227 77309 10228
rect 77451 10268 77493 10277
rect 77451 10228 77452 10268
rect 77492 10228 77493 10268
rect 77451 10219 77493 10228
rect 77635 10268 77693 10269
rect 77635 10228 77644 10268
rect 77684 10228 77693 10268
rect 77635 10227 77693 10228
rect 77835 10268 77877 10277
rect 77835 10228 77836 10268
rect 77876 10228 77877 10268
rect 77835 10219 77877 10228
rect 82531 10268 82589 10269
rect 82531 10228 82540 10268
rect 82580 10228 82589 10268
rect 82531 10227 82589 10228
rect 82731 10268 82773 10277
rect 82731 10228 82732 10268
rect 82772 10228 82773 10268
rect 82731 10219 82773 10228
rect 83203 10268 83261 10269
rect 83203 10228 83212 10268
rect 83252 10228 83261 10268
rect 83203 10227 83261 10228
rect 83403 10268 83445 10277
rect 83403 10228 83404 10268
rect 83444 10228 83445 10268
rect 83403 10219 83445 10228
rect 83587 10268 83645 10269
rect 83587 10228 83596 10268
rect 83636 10228 83645 10268
rect 83587 10227 83645 10228
rect 83787 10268 83829 10277
rect 83787 10228 83788 10268
rect 83828 10228 83829 10268
rect 83787 10219 83829 10228
rect 83971 10268 84029 10269
rect 83971 10228 83980 10268
rect 84020 10228 84029 10268
rect 83971 10227 84029 10228
rect 84171 10268 84213 10277
rect 84171 10228 84172 10268
rect 84212 10228 84213 10268
rect 84171 10219 84213 10228
rect 87819 10268 87861 10277
rect 87819 10228 87820 10268
rect 87860 10228 87861 10268
rect 87819 10219 87861 10228
rect 88003 10268 88061 10269
rect 88003 10228 88012 10268
rect 88052 10228 88061 10268
rect 88003 10227 88061 10228
rect 88203 10268 88245 10277
rect 88203 10228 88204 10268
rect 88244 10228 88245 10268
rect 88203 10219 88245 10228
rect 88387 10268 88445 10269
rect 88387 10228 88396 10268
rect 88436 10228 88445 10268
rect 88387 10227 88445 10228
rect 88579 10268 88637 10269
rect 88579 10228 88588 10268
rect 88628 10228 88637 10268
rect 88579 10227 88637 10228
rect 88683 10268 88725 10277
rect 88683 10228 88684 10268
rect 88724 10228 88725 10268
rect 88683 10219 88725 10228
rect 88779 10268 88821 10277
rect 88779 10228 88780 10268
rect 88820 10228 88821 10268
rect 89155 10268 89213 10269
rect 88779 10219 88821 10228
rect 88962 10253 89004 10262
rect 20130 10204 20172 10213
rect 88962 10213 88963 10253
rect 89003 10213 89004 10253
rect 89155 10228 89164 10268
rect 89204 10228 89213 10268
rect 89155 10227 89213 10228
rect 89451 10268 89493 10277
rect 89451 10228 89452 10268
rect 89492 10228 89493 10268
rect 89451 10219 89493 10228
rect 89635 10268 89693 10269
rect 89635 10228 89644 10268
rect 89684 10228 89693 10268
rect 89635 10227 89693 10228
rect 88962 10204 89004 10213
rect 12843 10184 12885 10193
rect 12843 10144 12844 10184
rect 12884 10144 12885 10184
rect 12843 10135 12885 10144
rect 21483 10184 21525 10193
rect 21483 10144 21484 10184
rect 21524 10144 21525 10184
rect 21483 10135 21525 10144
rect 25227 10184 25269 10193
rect 25227 10144 25228 10184
rect 25268 10144 25269 10184
rect 25227 10135 25269 10144
rect 32235 10184 32277 10193
rect 32235 10144 32236 10184
rect 32276 10144 32277 10184
rect 32235 10135 32277 10144
rect 15435 10100 15477 10109
rect 15435 10060 15436 10100
rect 15476 10060 15477 10100
rect 15435 10051 15477 10060
rect 16203 10100 16245 10109
rect 16203 10060 16204 10100
rect 16244 10060 16245 10100
rect 16203 10051 16245 10060
rect 21579 10100 21621 10109
rect 21579 10060 21580 10100
rect 21620 10060 21621 10100
rect 21579 10051 21621 10060
rect 25323 10100 25365 10109
rect 25323 10060 25324 10100
rect 25364 10060 25365 10100
rect 25323 10051 25365 10060
rect 30315 10100 30357 10109
rect 30315 10060 30316 10100
rect 30356 10060 30357 10100
rect 30315 10051 30357 10060
rect 30699 10100 30741 10109
rect 30699 10060 30700 10100
rect 30740 10060 30741 10100
rect 30699 10051 30741 10060
rect 37899 10100 37941 10109
rect 37899 10060 37900 10100
rect 37940 10060 37941 10100
rect 37899 10051 37941 10060
rect 58155 10100 58197 10109
rect 58155 10060 58156 10100
rect 58196 10060 58197 10100
rect 58155 10051 58197 10060
rect 58443 10100 58485 10109
rect 58443 10060 58444 10100
rect 58484 10060 58485 10100
rect 58443 10051 58485 10060
rect 58635 10100 58677 10109
rect 58635 10060 58636 10100
rect 58676 10060 58677 10100
rect 58635 10051 58677 10060
rect 60075 10100 60117 10109
rect 60075 10060 60076 10100
rect 60116 10060 60117 10100
rect 60075 10051 60117 10060
rect 69099 10100 69141 10109
rect 69099 10060 69100 10100
rect 69140 10060 69141 10100
rect 69099 10051 69141 10060
rect 74379 10100 74421 10109
rect 74379 10060 74380 10100
rect 74420 10060 74421 10100
rect 74379 10051 74421 10060
rect 87915 10100 87957 10109
rect 87915 10060 87916 10100
rect 87956 10060 87957 10100
rect 87915 10051 87957 10060
rect 89067 10100 89109 10109
rect 89067 10060 89068 10100
rect 89108 10060 89109 10100
rect 89067 10051 89109 10060
rect 11307 10016 11349 10025
rect 11307 9976 11308 10016
rect 11348 9976 11349 10016
rect 11307 9967 11349 9976
rect 11691 10016 11733 10025
rect 11691 9976 11692 10016
rect 11732 9976 11733 10016
rect 11691 9967 11733 9976
rect 12075 10016 12117 10025
rect 12075 9976 12076 10016
rect 12116 9976 12117 10016
rect 12075 9967 12117 9976
rect 12459 10016 12501 10025
rect 12459 9976 12460 10016
rect 12500 9976 12501 10016
rect 12459 9967 12501 9976
rect 14667 10016 14709 10025
rect 14667 9976 14668 10016
rect 14708 9976 14709 10016
rect 14667 9967 14709 9976
rect 15051 10016 15093 10025
rect 15051 9976 15052 10016
rect 15092 9976 15093 10016
rect 15051 9967 15093 9976
rect 15819 10016 15861 10025
rect 15819 9976 15820 10016
rect 15860 9976 15861 10016
rect 15819 9967 15861 9976
rect 18699 10016 18741 10025
rect 18699 9976 18700 10016
rect 18740 9976 18741 10016
rect 18699 9967 18741 9976
rect 19467 10016 19509 10025
rect 19467 9976 19468 10016
rect 19508 9976 19509 10016
rect 19467 9967 19509 9976
rect 20235 10016 20277 10025
rect 20235 9976 20236 10016
rect 20276 9976 20277 10016
rect 20235 9967 20277 9976
rect 24267 10016 24309 10025
rect 24267 9976 24268 10016
rect 24308 9976 24309 10016
rect 24267 9967 24309 9976
rect 24651 10016 24693 10025
rect 24651 9976 24652 10016
rect 24692 9976 24693 10016
rect 24651 9967 24693 9976
rect 31083 10016 31125 10025
rect 31083 9976 31084 10016
rect 31124 9976 31125 10016
rect 31083 9967 31125 9976
rect 31467 10016 31509 10025
rect 31467 9976 31468 10016
rect 31508 9976 31509 10016
rect 31467 9967 31509 9976
rect 32043 10016 32085 10025
rect 32043 9976 32044 10016
rect 32084 9976 32085 10016
rect 32043 9967 32085 9976
rect 35691 10016 35733 10025
rect 35691 9976 35692 10016
rect 35732 9976 35733 10016
rect 35691 9967 35733 9976
rect 36843 10016 36885 10025
rect 36843 9976 36844 10016
rect 36884 9976 36885 10016
rect 36843 9967 36885 9976
rect 37515 10016 37557 10025
rect 37515 9976 37516 10016
rect 37556 9976 37557 10016
rect 37515 9967 37557 9976
rect 38283 10016 38325 10025
rect 38283 9976 38284 10016
rect 38324 9976 38325 10016
rect 38283 9967 38325 9976
rect 38667 10016 38709 10025
rect 38667 9976 38668 10016
rect 38708 9976 38709 10016
rect 38667 9967 38709 9976
rect 39051 10016 39093 10025
rect 39051 9976 39052 10016
rect 39092 9976 39093 10016
rect 39051 9967 39093 9976
rect 57963 10016 58005 10025
rect 57963 9976 57964 10016
rect 58004 9976 58005 10016
rect 57963 9967 58005 9976
rect 59115 10016 59157 10025
rect 59115 9976 59116 10016
rect 59156 9976 59157 10016
rect 59115 9967 59157 9976
rect 60459 10016 60501 10025
rect 60459 9976 60460 10016
rect 60500 9976 60501 10016
rect 60459 9967 60501 9976
rect 71403 10016 71445 10025
rect 71403 9976 71404 10016
rect 71444 9976 71445 10016
rect 71403 9967 71445 9976
rect 73035 10016 73077 10025
rect 73035 9976 73036 10016
rect 73076 9976 73077 10016
rect 73035 9967 73077 9976
rect 76587 10016 76629 10025
rect 76587 9976 76588 10016
rect 76628 9976 76629 10016
rect 76587 9967 76629 9976
rect 76971 10016 77013 10025
rect 76971 9976 76972 10016
rect 77012 9976 77013 10016
rect 76971 9967 77013 9976
rect 77355 10016 77397 10025
rect 77355 9976 77356 10016
rect 77396 9976 77397 10016
rect 77355 9967 77397 9976
rect 77739 10016 77781 10025
rect 77739 9976 77740 10016
rect 77780 9976 77781 10016
rect 77739 9967 77781 9976
rect 82635 10016 82677 10025
rect 82635 9976 82636 10016
rect 82676 9976 82677 10016
rect 82635 9967 82677 9976
rect 83307 10016 83349 10025
rect 83307 9976 83308 10016
rect 83348 9976 83349 10016
rect 83307 9967 83349 9976
rect 83691 10016 83733 10025
rect 83691 9976 83692 10016
rect 83732 9976 83733 10016
rect 83691 9967 83733 9976
rect 89547 10016 89589 10025
rect 89547 9976 89548 10016
rect 89588 9976 89589 10016
rect 89547 9967 89589 9976
rect 1152 9848 98784 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 64168 9848
rect 64208 9808 64250 9848
rect 64290 9808 64332 9848
rect 64372 9808 64414 9848
rect 64454 9808 64496 9848
rect 64536 9808 79288 9848
rect 79328 9808 79370 9848
rect 79410 9808 79452 9848
rect 79492 9808 79534 9848
rect 79574 9808 79616 9848
rect 79656 9808 94408 9848
rect 94448 9808 94490 9848
rect 94530 9808 94572 9848
rect 94612 9808 94654 9848
rect 94694 9808 94736 9848
rect 94776 9808 98784 9848
rect 1152 9784 98784 9808
rect 34539 9680 34581 9689
rect 34539 9640 34540 9680
rect 34580 9640 34581 9680
rect 34539 9631 34581 9640
rect 56235 9680 56277 9689
rect 56235 9640 56236 9680
rect 56276 9640 56277 9680
rect 56235 9631 56277 9640
rect 56619 9680 56661 9689
rect 56619 9640 56620 9680
rect 56660 9640 56661 9680
rect 56619 9631 56661 9640
rect 73803 9680 73845 9689
rect 73803 9640 73804 9680
rect 73844 9640 73845 9680
rect 73803 9631 73845 9640
rect 77451 9680 77493 9689
rect 77451 9640 77452 9680
rect 77492 9640 77493 9680
rect 77451 9631 77493 9640
rect 36363 9596 36405 9605
rect 36363 9556 36364 9596
rect 36404 9556 36405 9596
rect 36363 9547 36405 9556
rect 48459 9596 48501 9605
rect 48459 9556 48460 9596
rect 48500 9556 48501 9596
rect 48459 9547 48501 9556
rect 48651 9596 48693 9605
rect 48651 9556 48652 9596
rect 48692 9556 48693 9596
rect 48651 9547 48693 9556
rect 51147 9596 51189 9605
rect 51147 9556 51148 9596
rect 51188 9556 51189 9596
rect 51147 9547 51189 9556
rect 52299 9596 52341 9605
rect 52299 9556 52300 9596
rect 52340 9556 52341 9596
rect 52299 9547 52341 9556
rect 55851 9596 55893 9605
rect 55851 9556 55852 9596
rect 55892 9556 55893 9596
rect 55851 9547 55893 9556
rect 58731 9596 58773 9605
rect 58731 9556 58732 9596
rect 58772 9556 58773 9596
rect 58731 9547 58773 9556
rect 59883 9596 59925 9605
rect 59883 9556 59884 9596
rect 59924 9556 59925 9596
rect 59883 9547 59925 9556
rect 60363 9596 60405 9605
rect 60363 9556 60364 9596
rect 60404 9556 60405 9596
rect 60363 9547 60405 9556
rect 60843 9596 60885 9605
rect 60843 9556 60844 9596
rect 60884 9556 60885 9596
rect 60843 9547 60885 9556
rect 72075 9596 72117 9605
rect 72075 9556 72076 9596
rect 72116 9556 72117 9596
rect 72075 9547 72117 9556
rect 40683 9512 40725 9521
rect 40683 9472 40684 9512
rect 40724 9472 40725 9512
rect 40683 9463 40725 9472
rect 48259 9512 48317 9513
rect 48259 9472 48268 9512
rect 48308 9472 48317 9512
rect 48259 9471 48317 9472
rect 49803 9512 49845 9521
rect 49803 9472 49804 9512
rect 49844 9472 49845 9512
rect 49803 9463 49845 9472
rect 11595 9428 11637 9437
rect 11595 9388 11596 9428
rect 11636 9388 11637 9428
rect 11595 9379 11637 9388
rect 11779 9428 11837 9429
rect 11779 9388 11788 9428
rect 11828 9388 11837 9428
rect 11779 9387 11837 9388
rect 12067 9428 12125 9429
rect 12067 9388 12076 9428
rect 12116 9388 12125 9428
rect 12067 9387 12125 9388
rect 12259 9428 12317 9429
rect 12259 9388 12268 9428
rect 12308 9388 12317 9428
rect 12259 9387 12317 9388
rect 14571 9428 14613 9437
rect 14571 9388 14572 9428
rect 14612 9388 14613 9428
rect 14571 9379 14613 9388
rect 14667 9428 14709 9437
rect 14667 9388 14668 9428
rect 14708 9388 14709 9428
rect 14667 9379 14709 9388
rect 14755 9428 14813 9429
rect 14755 9388 14764 9428
rect 14804 9388 14813 9428
rect 14755 9387 14813 9388
rect 14955 9428 14997 9437
rect 14955 9388 14956 9428
rect 14996 9388 14997 9428
rect 14955 9379 14997 9388
rect 15139 9428 15197 9429
rect 15139 9388 15148 9428
rect 15188 9388 15197 9428
rect 15139 9387 15197 9388
rect 15339 9428 15381 9437
rect 15339 9388 15340 9428
rect 15380 9388 15381 9428
rect 15339 9379 15381 9388
rect 15523 9428 15581 9429
rect 15523 9388 15532 9428
rect 15572 9388 15581 9428
rect 15523 9387 15581 9388
rect 15715 9428 15773 9429
rect 15715 9388 15724 9428
rect 15764 9388 15773 9428
rect 15715 9387 15773 9388
rect 15915 9428 15957 9437
rect 15915 9388 15916 9428
rect 15956 9388 15957 9428
rect 15915 9379 15957 9388
rect 16107 9428 16149 9437
rect 16107 9388 16108 9428
rect 16148 9388 16149 9428
rect 16107 9379 16149 9388
rect 16291 9428 16349 9429
rect 16291 9388 16300 9428
rect 16340 9388 16349 9428
rect 16291 9387 16349 9388
rect 18987 9428 19029 9437
rect 18987 9388 18988 9428
rect 19028 9388 19029 9428
rect 18987 9379 19029 9388
rect 19171 9428 19229 9429
rect 19171 9388 19180 9428
rect 19220 9388 19229 9428
rect 19171 9387 19229 9388
rect 19371 9428 19413 9437
rect 19371 9388 19372 9428
rect 19412 9388 19413 9428
rect 19371 9379 19413 9388
rect 19555 9428 19613 9429
rect 19555 9388 19564 9428
rect 19604 9388 19613 9428
rect 19555 9387 19613 9388
rect 19747 9428 19805 9429
rect 19747 9388 19756 9428
rect 19796 9388 19805 9428
rect 19747 9387 19805 9388
rect 19947 9428 19989 9437
rect 19947 9388 19948 9428
rect 19988 9388 19989 9428
rect 19947 9379 19989 9388
rect 24171 9428 24213 9437
rect 24171 9388 24172 9428
rect 24212 9388 24213 9428
rect 24171 9379 24213 9388
rect 24355 9428 24413 9429
rect 24355 9388 24364 9428
rect 24404 9388 24413 9428
rect 24355 9387 24413 9388
rect 24555 9428 24597 9437
rect 24555 9388 24556 9428
rect 24596 9388 24597 9428
rect 24555 9379 24597 9388
rect 24739 9428 24797 9429
rect 24739 9388 24748 9428
rect 24788 9388 24797 9428
rect 24739 9387 24797 9388
rect 25219 9428 25277 9429
rect 25219 9388 25228 9428
rect 25268 9388 25277 9428
rect 25219 9387 25277 9388
rect 25411 9428 25469 9429
rect 25411 9388 25420 9428
rect 25460 9388 25469 9428
rect 25411 9387 25469 9388
rect 30019 9428 30077 9429
rect 30019 9388 30028 9428
rect 30068 9388 30077 9428
rect 30019 9387 30077 9388
rect 30211 9428 30269 9429
rect 30211 9388 30220 9428
rect 30260 9388 30269 9428
rect 30211 9387 30269 9388
rect 30603 9428 30645 9437
rect 30603 9388 30604 9428
rect 30644 9388 30645 9428
rect 30603 9379 30645 9388
rect 30787 9428 30845 9429
rect 30787 9388 30796 9428
rect 30836 9388 30845 9428
rect 31083 9428 31125 9437
rect 30787 9387 30845 9388
rect 30987 9415 31029 9424
rect 30987 9375 30988 9415
rect 31028 9375 31029 9415
rect 31083 9388 31084 9428
rect 31124 9388 31125 9428
rect 31083 9379 31125 9388
rect 31171 9428 31229 9429
rect 31171 9388 31180 9428
rect 31220 9388 31229 9428
rect 31171 9387 31229 9388
rect 34443 9428 34485 9437
rect 34443 9388 34444 9428
rect 34484 9388 34485 9428
rect 34443 9379 34485 9388
rect 34627 9428 34685 9429
rect 34627 9388 34636 9428
rect 34676 9388 34685 9428
rect 34627 9387 34685 9388
rect 34827 9428 34869 9437
rect 34827 9388 34828 9428
rect 34868 9388 34869 9428
rect 34827 9379 34869 9388
rect 35011 9428 35069 9429
rect 35011 9388 35020 9428
rect 35060 9388 35069 9428
rect 35011 9387 35069 9388
rect 36267 9428 36309 9437
rect 36267 9388 36268 9428
rect 36308 9388 36309 9428
rect 36267 9379 36309 9388
rect 36451 9428 36509 9429
rect 36451 9388 36460 9428
rect 36500 9388 36509 9428
rect 36451 9387 36509 9388
rect 36651 9428 36693 9437
rect 36651 9388 36652 9428
rect 36692 9388 36693 9428
rect 36651 9379 36693 9388
rect 36835 9428 36893 9429
rect 36835 9388 36844 9428
rect 36884 9388 36893 9428
rect 36835 9387 36893 9388
rect 37123 9428 37181 9429
rect 37123 9388 37132 9428
rect 37172 9388 37181 9428
rect 37123 9387 37181 9388
rect 37315 9428 37373 9429
rect 37315 9388 37324 9428
rect 37364 9388 37373 9428
rect 37315 9387 37373 9388
rect 37995 9428 38037 9437
rect 37995 9388 37996 9428
rect 38036 9388 38037 9428
rect 37995 9379 38037 9388
rect 38179 9428 38237 9429
rect 38179 9388 38188 9428
rect 38228 9388 38237 9428
rect 38179 9387 38237 9388
rect 38379 9428 38421 9437
rect 38379 9388 38380 9428
rect 38420 9388 38421 9428
rect 38379 9379 38421 9388
rect 38563 9428 38621 9429
rect 38563 9388 38572 9428
rect 38612 9388 38621 9428
rect 38563 9387 38621 9388
rect 38763 9428 38805 9437
rect 38763 9388 38764 9428
rect 38804 9388 38805 9428
rect 38763 9379 38805 9388
rect 38947 9428 39005 9429
rect 38947 9388 38956 9428
rect 38996 9388 39005 9428
rect 38947 9387 39005 9388
rect 39331 9428 39389 9429
rect 39331 9388 39340 9428
rect 39380 9388 39389 9428
rect 39331 9387 39389 9388
rect 40291 9428 40349 9429
rect 40291 9388 40300 9428
rect 40340 9388 40349 9428
rect 40291 9387 40349 9388
rect 41539 9428 41597 9429
rect 41539 9388 41548 9428
rect 41588 9388 41597 9428
rect 41539 9387 41597 9388
rect 42307 9428 42365 9429
rect 42307 9388 42316 9428
rect 42356 9388 42365 9428
rect 42307 9387 42365 9388
rect 43267 9428 43325 9429
rect 43267 9388 43276 9428
rect 43316 9388 43325 9428
rect 43267 9387 43325 9388
rect 48843 9428 48885 9437
rect 48843 9388 48844 9428
rect 48884 9388 48885 9428
rect 48843 9379 48885 9388
rect 48939 9428 48981 9437
rect 48939 9388 48940 9428
rect 48980 9388 48981 9428
rect 48939 9379 48981 9388
rect 49515 9428 49557 9437
rect 49515 9388 49516 9428
rect 49556 9388 49557 9428
rect 49515 9379 49557 9388
rect 49611 9428 49653 9437
rect 49611 9388 49612 9428
rect 49652 9388 49653 9428
rect 49611 9379 49653 9388
rect 51339 9428 51381 9437
rect 51339 9388 51340 9428
rect 51380 9388 51381 9428
rect 51339 9379 51381 9388
rect 51435 9428 51477 9437
rect 51435 9388 51436 9428
rect 51476 9388 51477 9428
rect 51435 9379 51477 9388
rect 52011 9428 52053 9437
rect 52011 9388 52012 9428
rect 52052 9388 52053 9428
rect 52011 9379 52053 9388
rect 52107 9428 52149 9437
rect 52107 9388 52108 9428
rect 52148 9388 52149 9428
rect 52107 9379 52149 9388
rect 52483 9428 52541 9429
rect 52483 9388 52492 9428
rect 52532 9388 52541 9428
rect 52483 9387 52541 9388
rect 53443 9428 53501 9429
rect 53443 9388 53452 9428
rect 53492 9388 53501 9428
rect 53443 9387 53501 9388
rect 54787 9428 54845 9429
rect 54787 9388 54796 9428
rect 54836 9388 54845 9428
rect 54787 9387 54845 9388
rect 54987 9428 55029 9437
rect 54987 9388 54988 9428
rect 55028 9388 55029 9428
rect 54987 9379 55029 9388
rect 55755 9428 55797 9437
rect 55755 9388 55756 9428
rect 55796 9388 55797 9428
rect 55755 9379 55797 9388
rect 55939 9428 55997 9429
rect 55939 9388 55948 9428
rect 55988 9388 55997 9428
rect 55939 9387 55997 9388
rect 56139 9428 56181 9437
rect 56139 9388 56140 9428
rect 56180 9388 56181 9428
rect 56139 9379 56181 9388
rect 56323 9428 56381 9429
rect 56323 9388 56332 9428
rect 56372 9388 56381 9428
rect 56323 9387 56381 9388
rect 56523 9428 56565 9437
rect 56523 9388 56524 9428
rect 56564 9388 56565 9428
rect 56523 9379 56565 9388
rect 56707 9428 56765 9429
rect 56707 9388 56716 9428
rect 56756 9388 56765 9428
rect 56707 9387 56765 9388
rect 58731 9428 58773 9437
rect 58731 9388 58732 9428
rect 58772 9388 58773 9428
rect 58731 9379 58773 9388
rect 59019 9428 59061 9437
rect 59019 9388 59020 9428
rect 59060 9388 59061 9428
rect 59019 9379 59061 9388
rect 59211 9428 59253 9437
rect 59211 9388 59212 9428
rect 59252 9388 59253 9428
rect 59211 9379 59253 9388
rect 59403 9428 59445 9437
rect 59403 9388 59404 9428
rect 59444 9388 59445 9428
rect 59403 9379 59445 9388
rect 59595 9428 59637 9437
rect 59595 9388 59596 9428
rect 59636 9388 59637 9428
rect 59595 9379 59637 9388
rect 59883 9428 59925 9437
rect 59883 9388 59884 9428
rect 59924 9388 59925 9428
rect 59883 9379 59925 9388
rect 60363 9428 60405 9437
rect 60363 9388 60364 9428
rect 60404 9388 60405 9428
rect 60363 9379 60405 9388
rect 60843 9428 60885 9437
rect 60843 9388 60844 9428
rect 60884 9388 60885 9428
rect 60843 9379 60885 9388
rect 62083 9428 62141 9429
rect 62083 9388 62092 9428
rect 62132 9388 62141 9428
rect 62083 9387 62141 9388
rect 65155 9428 65213 9429
rect 65155 9388 65164 9428
rect 65204 9388 65213 9428
rect 65155 9387 65213 9388
rect 66115 9428 66173 9429
rect 66115 9388 66124 9428
rect 66164 9388 66173 9428
rect 66115 9387 66173 9388
rect 70531 9428 70589 9429
rect 70531 9388 70540 9428
rect 70580 9388 70589 9428
rect 70531 9387 70589 9388
rect 70723 9428 70781 9429
rect 70723 9388 70732 9428
rect 70772 9388 70781 9428
rect 70723 9387 70781 9388
rect 71587 9428 71645 9429
rect 71587 9388 71596 9428
rect 71636 9388 71645 9428
rect 71587 9387 71645 9388
rect 71787 9428 71829 9437
rect 71787 9388 71788 9428
rect 71828 9388 71829 9428
rect 71787 9379 71829 9388
rect 71971 9428 72029 9429
rect 71971 9388 71980 9428
rect 72020 9388 72029 9428
rect 71971 9387 72029 9388
rect 72171 9428 72213 9437
rect 72171 9388 72172 9428
rect 72212 9388 72213 9428
rect 72171 9379 72213 9388
rect 73123 9428 73181 9429
rect 73123 9388 73132 9428
rect 73172 9388 73181 9428
rect 73123 9387 73181 9388
rect 73323 9428 73365 9437
rect 73323 9388 73324 9428
rect 73364 9388 73365 9428
rect 73323 9379 73365 9388
rect 73699 9428 73757 9429
rect 73699 9388 73708 9428
rect 73748 9388 73757 9428
rect 73699 9387 73757 9388
rect 73899 9428 73941 9437
rect 73899 9388 73900 9428
rect 73940 9388 73941 9428
rect 73899 9379 73941 9388
rect 76963 9428 77021 9429
rect 76963 9388 76972 9428
rect 77012 9388 77021 9428
rect 76963 9387 77021 9388
rect 77163 9428 77205 9437
rect 77163 9388 77164 9428
rect 77204 9388 77205 9428
rect 77163 9379 77205 9388
rect 77347 9428 77405 9429
rect 77347 9388 77356 9428
rect 77396 9388 77405 9428
rect 77347 9387 77405 9388
rect 77547 9428 77589 9437
rect 77547 9388 77548 9428
rect 77588 9388 77589 9428
rect 77547 9379 77589 9388
rect 77739 9428 77781 9437
rect 77739 9388 77740 9428
rect 77780 9388 77781 9428
rect 77739 9379 77781 9388
rect 77923 9428 77981 9429
rect 77923 9388 77932 9428
rect 77972 9388 77981 9428
rect 77923 9387 77981 9388
rect 78307 9428 78365 9429
rect 78307 9388 78316 9428
rect 78356 9388 78365 9428
rect 78307 9387 78365 9388
rect 78507 9428 78549 9437
rect 78507 9388 78508 9428
rect 78548 9388 78549 9428
rect 78507 9379 78549 9388
rect 79267 9428 79325 9429
rect 79267 9388 79276 9428
rect 79316 9388 79325 9428
rect 79267 9387 79325 9388
rect 80227 9428 80285 9429
rect 80227 9388 80236 9428
rect 80276 9388 80285 9428
rect 80227 9387 80285 9388
rect 80611 9428 80669 9429
rect 80611 9388 80620 9428
rect 80660 9388 80669 9428
rect 80611 9387 80669 9388
rect 80811 9428 80853 9437
rect 80811 9388 80812 9428
rect 80852 9388 80853 9428
rect 80811 9379 80853 9388
rect 81003 9428 81045 9437
rect 81003 9388 81004 9428
rect 81044 9388 81045 9428
rect 81003 9379 81045 9388
rect 81187 9428 81245 9429
rect 81187 9388 81196 9428
rect 81236 9388 81245 9428
rect 81187 9387 81245 9388
rect 81859 9428 81917 9429
rect 81859 9388 81868 9428
rect 81908 9388 81917 9428
rect 81859 9387 81917 9388
rect 82059 9428 82101 9437
rect 82059 9388 82060 9428
rect 82100 9388 82101 9428
rect 82059 9379 82101 9388
rect 87139 9428 87197 9429
rect 87139 9388 87148 9428
rect 87188 9388 87197 9428
rect 87139 9387 87197 9388
rect 87339 9428 87381 9437
rect 87339 9388 87340 9428
rect 87380 9388 87381 9428
rect 87339 9379 87381 9388
rect 87723 9428 87765 9437
rect 87723 9388 87724 9428
rect 87764 9388 87765 9428
rect 87723 9379 87765 9388
rect 87819 9428 87861 9437
rect 87819 9388 87820 9428
rect 87860 9388 87861 9428
rect 87819 9379 87861 9388
rect 87907 9428 87965 9429
rect 87907 9388 87916 9428
rect 87956 9388 87965 9428
rect 87907 9387 87965 9388
rect 88195 9428 88253 9429
rect 88195 9388 88204 9428
rect 88244 9388 88253 9428
rect 88195 9387 88253 9388
rect 88395 9428 88437 9437
rect 88395 9388 88396 9428
rect 88436 9388 88437 9428
rect 88395 9379 88437 9388
rect 88579 9428 88637 9429
rect 88579 9388 88588 9428
rect 88628 9388 88637 9428
rect 88579 9387 88637 9388
rect 88779 9428 88821 9437
rect 88779 9388 88780 9428
rect 88820 9388 88821 9428
rect 88779 9379 88821 9388
rect 88971 9428 89013 9437
rect 88971 9388 88972 9428
rect 89012 9388 89013 9428
rect 88971 9379 89013 9388
rect 89155 9428 89213 9429
rect 89155 9388 89164 9428
rect 89204 9388 89213 9428
rect 89155 9387 89213 9388
rect 89347 9428 89405 9429
rect 89347 9388 89356 9428
rect 89396 9388 89405 9428
rect 89347 9387 89405 9388
rect 89547 9428 89589 9437
rect 89547 9388 89548 9428
rect 89588 9388 89589 9428
rect 89547 9379 89589 9388
rect 89739 9428 89781 9437
rect 89739 9388 89740 9428
rect 89780 9388 89781 9428
rect 89739 9379 89781 9388
rect 89923 9428 89981 9429
rect 89923 9388 89932 9428
rect 89972 9388 89981 9428
rect 89923 9387 89981 9388
rect 30987 9366 31029 9375
rect 11691 9344 11733 9353
rect 11691 9304 11692 9344
rect 11732 9304 11733 9344
rect 11691 9295 11733 9304
rect 15051 9344 15093 9353
rect 15051 9304 15052 9344
rect 15092 9304 15093 9344
rect 15051 9295 15093 9304
rect 15435 9344 15477 9353
rect 15435 9304 15436 9344
rect 15476 9304 15477 9344
rect 15435 9295 15477 9304
rect 15819 9344 15861 9353
rect 15819 9304 15820 9344
rect 15860 9304 15861 9344
rect 15819 9295 15861 9304
rect 16203 9344 16245 9353
rect 16203 9304 16204 9344
rect 16244 9304 16245 9344
rect 16203 9295 16245 9304
rect 19083 9344 19125 9353
rect 19083 9304 19084 9344
rect 19124 9304 19125 9344
rect 19083 9295 19125 9304
rect 19467 9344 19509 9353
rect 19467 9304 19468 9344
rect 19508 9304 19509 9344
rect 19467 9295 19509 9304
rect 19851 9344 19893 9353
rect 19851 9304 19852 9344
rect 19892 9304 19893 9344
rect 19851 9295 19893 9304
rect 24267 9344 24309 9353
rect 24267 9304 24268 9344
rect 24308 9304 24309 9344
rect 24267 9295 24309 9304
rect 24651 9344 24693 9353
rect 24651 9304 24652 9344
rect 24692 9304 24693 9344
rect 24651 9295 24693 9304
rect 30699 9344 30741 9353
rect 30699 9304 30700 9344
rect 30740 9304 30741 9344
rect 30699 9295 30741 9304
rect 34923 9344 34965 9353
rect 34923 9304 34924 9344
rect 34964 9304 34965 9344
rect 34923 9295 34965 9304
rect 36747 9344 36789 9353
rect 36747 9304 36748 9344
rect 36788 9304 36789 9344
rect 36747 9295 36789 9304
rect 38091 9344 38133 9353
rect 38091 9304 38092 9344
rect 38132 9304 38133 9344
rect 38091 9295 38133 9304
rect 38475 9344 38517 9353
rect 38475 9304 38476 9344
rect 38516 9304 38517 9344
rect 38475 9295 38517 9304
rect 38859 9344 38901 9353
rect 38859 9304 38860 9344
rect 38900 9304 38901 9344
rect 38859 9295 38901 9304
rect 54891 9344 54933 9353
rect 54891 9304 54892 9344
rect 54932 9304 54933 9344
rect 54891 9295 54933 9304
rect 62947 9344 63005 9345
rect 62947 9304 62956 9344
rect 62996 9304 63005 9344
rect 62947 9303 63005 9304
rect 71691 9344 71733 9353
rect 71691 9304 71692 9344
rect 71732 9304 71733 9344
rect 71691 9295 71733 9304
rect 73227 9344 73269 9353
rect 73227 9304 73228 9344
rect 73268 9304 73269 9344
rect 73227 9295 73269 9304
rect 77067 9344 77109 9353
rect 77067 9304 77068 9344
rect 77108 9304 77109 9344
rect 77067 9295 77109 9304
rect 77835 9344 77877 9353
rect 77835 9304 77836 9344
rect 77876 9304 77877 9344
rect 77835 9295 77877 9304
rect 78411 9344 78453 9353
rect 78411 9304 78412 9344
rect 78452 9304 78453 9344
rect 78411 9295 78453 9304
rect 80715 9344 80757 9353
rect 80715 9304 80716 9344
rect 80756 9304 80757 9344
rect 80715 9295 80757 9304
rect 81099 9344 81141 9353
rect 81099 9304 81100 9344
rect 81140 9304 81141 9344
rect 81099 9295 81141 9304
rect 81963 9344 82005 9353
rect 81963 9304 81964 9344
rect 82004 9304 82005 9344
rect 81963 9295 82005 9304
rect 87243 9344 87285 9353
rect 87243 9304 87244 9344
rect 87284 9304 87285 9344
rect 87243 9295 87285 9304
rect 88299 9344 88341 9353
rect 88299 9304 88300 9344
rect 88340 9304 88341 9344
rect 88299 9295 88341 9304
rect 88683 9344 88725 9353
rect 88683 9304 88684 9344
rect 88724 9304 88725 9344
rect 88683 9295 88725 9304
rect 89067 9344 89109 9353
rect 89067 9304 89068 9344
rect 89108 9304 89109 9344
rect 89067 9295 89109 9304
rect 89451 9344 89493 9353
rect 89451 9304 89452 9344
rect 89492 9304 89493 9344
rect 89451 9295 89493 9304
rect 89835 9344 89877 9353
rect 89835 9304 89836 9344
rect 89876 9304 89877 9344
rect 89835 9295 89877 9304
rect 48931 9260 48989 9261
rect 48931 9220 48940 9260
rect 48980 9220 48989 9260
rect 48931 9219 48989 9220
rect 49507 9260 49565 9261
rect 49507 9220 49516 9260
rect 49556 9220 49565 9260
rect 49507 9219 49565 9220
rect 51427 9260 51485 9261
rect 51427 9220 51436 9260
rect 51476 9220 51485 9260
rect 51427 9219 51485 9220
rect 52003 9260 52061 9261
rect 52003 9220 52012 9260
rect 52052 9220 52061 9260
rect 52003 9219 52061 9220
rect 58539 9260 58581 9269
rect 58539 9220 58540 9260
rect 58580 9220 58581 9260
rect 58539 9211 58581 9220
rect 59115 9260 59157 9269
rect 59115 9220 59116 9260
rect 59156 9220 59157 9260
rect 59115 9211 59157 9220
rect 59499 9260 59541 9269
rect 59499 9220 59500 9260
rect 59540 9220 59541 9260
rect 59499 9211 59541 9220
rect 60075 9260 60117 9269
rect 60075 9220 60076 9260
rect 60116 9220 60117 9260
rect 60075 9211 60117 9220
rect 60555 9260 60597 9269
rect 60555 9220 60556 9260
rect 60596 9220 60597 9260
rect 60555 9211 60597 9220
rect 61035 9260 61077 9269
rect 61035 9220 61036 9260
rect 61076 9220 61077 9260
rect 61035 9211 61077 9220
rect 1152 9092 98784 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 65408 9092
rect 65448 9052 65490 9092
rect 65530 9052 65572 9092
rect 65612 9052 65654 9092
rect 65694 9052 65736 9092
rect 65776 9052 80528 9092
rect 80568 9052 80610 9092
rect 80650 9052 80692 9092
rect 80732 9052 80774 9092
rect 80814 9052 80856 9092
rect 80896 9052 95648 9092
rect 95688 9052 95730 9092
rect 95770 9052 95812 9092
rect 95852 9052 95894 9092
rect 95934 9052 95976 9092
rect 96016 9052 98784 9092
rect 1152 9028 98784 9052
rect 15339 8924 15381 8933
rect 15339 8884 15340 8924
rect 15380 8884 15381 8924
rect 15339 8875 15381 8884
rect 31947 8924 31989 8933
rect 31947 8884 31948 8924
rect 31988 8884 31989 8924
rect 31947 8875 31989 8884
rect 45187 8924 45245 8925
rect 45187 8884 45196 8924
rect 45236 8884 45245 8924
rect 45187 8883 45245 8884
rect 49315 8924 49373 8925
rect 49315 8884 49324 8924
rect 49364 8884 49373 8924
rect 49315 8883 49373 8884
rect 49891 8924 49949 8925
rect 49891 8884 49900 8924
rect 49940 8884 49949 8924
rect 49891 8883 49949 8884
rect 52579 8924 52637 8925
rect 52579 8884 52588 8924
rect 52628 8884 52637 8924
rect 52579 8883 52637 8884
rect 55467 8924 55509 8933
rect 55467 8884 55468 8924
rect 55508 8884 55509 8924
rect 55467 8875 55509 8884
rect 58731 8924 58773 8933
rect 58731 8884 58732 8924
rect 58772 8884 58773 8924
rect 58731 8875 58773 8884
rect 9771 8840 9813 8849
rect 9771 8800 9772 8840
rect 9812 8800 9813 8840
rect 9771 8791 9813 8800
rect 11595 8840 11637 8849
rect 11595 8800 11596 8840
rect 11636 8800 11637 8840
rect 11595 8791 11637 8800
rect 11979 8840 12021 8849
rect 11979 8800 11980 8840
rect 12020 8800 12021 8840
rect 11979 8791 12021 8800
rect 12363 8840 12405 8849
rect 12363 8800 12364 8840
rect 12404 8800 12405 8840
rect 12363 8791 12405 8800
rect 18699 8840 18741 8849
rect 18699 8800 18700 8840
rect 18740 8800 18741 8840
rect 18699 8791 18741 8800
rect 25035 8840 25077 8849
rect 25035 8800 25036 8840
rect 25076 8800 25077 8840
rect 25035 8791 25077 8800
rect 27915 8840 27957 8849
rect 27915 8800 27916 8840
rect 27956 8800 27957 8840
rect 27915 8791 27957 8800
rect 28299 8840 28341 8849
rect 28299 8800 28300 8840
rect 28340 8800 28341 8840
rect 28299 8791 28341 8800
rect 28683 8840 28725 8849
rect 28683 8800 28684 8840
rect 28724 8800 28725 8840
rect 28683 8791 28725 8800
rect 34827 8840 34869 8849
rect 34827 8800 34828 8840
rect 34868 8800 34869 8840
rect 34827 8791 34869 8800
rect 50179 8840 50237 8841
rect 50179 8800 50188 8840
rect 50228 8800 50237 8840
rect 50179 8799 50237 8800
rect 70059 8840 70101 8849
rect 70059 8800 70060 8840
rect 70100 8800 70101 8840
rect 70059 8791 70101 8800
rect 70539 8840 70581 8849
rect 70539 8800 70540 8840
rect 70580 8800 70581 8840
rect 70539 8791 70581 8800
rect 70923 8840 70965 8849
rect 70923 8800 70924 8840
rect 70964 8800 70965 8840
rect 70923 8791 70965 8800
rect 74667 8840 74709 8849
rect 74667 8800 74668 8840
rect 74708 8800 74709 8840
rect 74667 8791 74709 8800
rect 75051 8840 75093 8849
rect 75051 8800 75052 8840
rect 75092 8800 75093 8840
rect 75051 8791 75093 8800
rect 75435 8840 75477 8849
rect 75435 8800 75436 8840
rect 75476 8800 75477 8840
rect 75435 8791 75477 8800
rect 78795 8840 78837 8849
rect 78795 8800 78796 8840
rect 78836 8800 78837 8840
rect 78795 8791 78837 8800
rect 80907 8840 80949 8849
rect 80907 8800 80908 8840
rect 80948 8800 80949 8840
rect 80907 8791 80949 8800
rect 81675 8840 81717 8849
rect 81675 8800 81676 8840
rect 81716 8800 81717 8840
rect 81675 8791 81717 8800
rect 82059 8840 82101 8849
rect 82059 8800 82060 8840
rect 82100 8800 82101 8840
rect 82059 8791 82101 8800
rect 83211 8840 83253 8849
rect 83211 8800 83212 8840
rect 83252 8800 83253 8840
rect 83211 8791 83253 8800
rect 83595 8840 83637 8849
rect 83595 8800 83596 8840
rect 83636 8800 83637 8840
rect 83595 8791 83637 8800
rect 86955 8840 86997 8849
rect 86955 8800 86956 8840
rect 86996 8800 86997 8840
rect 86955 8791 86997 8800
rect 87723 8840 87765 8849
rect 87723 8800 87724 8840
rect 87764 8800 87765 8840
rect 87723 8791 87765 8800
rect 89067 8840 89109 8849
rect 89067 8800 89068 8840
rect 89108 8800 89109 8840
rect 89067 8791 89109 8800
rect 9675 8756 9717 8765
rect 9675 8716 9676 8756
rect 9716 8716 9717 8756
rect 9675 8707 9717 8716
rect 9859 8756 9917 8757
rect 9859 8716 9868 8756
rect 9908 8716 9917 8756
rect 9859 8715 9917 8716
rect 10059 8756 10101 8765
rect 10059 8716 10060 8756
rect 10100 8716 10101 8756
rect 10059 8707 10101 8716
rect 10243 8756 10301 8757
rect 10243 8716 10252 8756
rect 10292 8716 10301 8756
rect 10243 8715 10301 8716
rect 11115 8756 11157 8765
rect 11115 8716 11116 8756
rect 11156 8716 11157 8756
rect 11115 8707 11157 8716
rect 11299 8756 11357 8757
rect 11299 8716 11308 8756
rect 11348 8716 11357 8756
rect 11299 8715 11357 8716
rect 11499 8756 11541 8765
rect 11499 8716 11500 8756
rect 11540 8716 11541 8756
rect 11499 8707 11541 8716
rect 11683 8756 11741 8757
rect 11683 8716 11692 8756
rect 11732 8716 11741 8756
rect 11683 8715 11741 8716
rect 11883 8756 11925 8765
rect 11883 8716 11884 8756
rect 11924 8716 11925 8756
rect 11883 8707 11925 8716
rect 12067 8756 12125 8757
rect 12067 8716 12076 8756
rect 12116 8716 12125 8756
rect 12067 8715 12125 8716
rect 12267 8756 12309 8765
rect 12267 8716 12268 8756
rect 12308 8716 12309 8756
rect 12267 8707 12309 8716
rect 12451 8756 12509 8757
rect 12451 8716 12460 8756
rect 12500 8716 12509 8756
rect 12451 8715 12509 8716
rect 15723 8756 15765 8765
rect 15723 8716 15724 8756
rect 15764 8716 15765 8756
rect 15723 8707 15765 8716
rect 18595 8756 18653 8757
rect 18595 8716 18604 8756
rect 18644 8716 18653 8756
rect 18595 8715 18653 8716
rect 18795 8756 18837 8765
rect 18795 8716 18796 8756
rect 18836 8716 18837 8756
rect 18795 8707 18837 8716
rect 20611 8756 20669 8757
rect 20611 8716 20620 8756
rect 20660 8716 20669 8756
rect 20611 8715 20669 8716
rect 20803 8756 20861 8757
rect 20803 8716 20812 8756
rect 20852 8716 20861 8756
rect 20803 8715 20861 8716
rect 24163 8756 24221 8757
rect 24163 8716 24172 8756
rect 24212 8716 24221 8756
rect 24163 8715 24221 8716
rect 24363 8756 24405 8765
rect 24363 8716 24364 8756
rect 24404 8716 24405 8756
rect 24363 8707 24405 8716
rect 24555 8756 24597 8765
rect 24555 8716 24556 8756
rect 24596 8716 24597 8756
rect 24555 8707 24597 8716
rect 24739 8756 24797 8757
rect 24739 8716 24748 8756
rect 24788 8716 24797 8756
rect 24739 8715 24797 8716
rect 24939 8756 24981 8765
rect 24939 8716 24940 8756
rect 24980 8716 24981 8756
rect 24939 8707 24981 8716
rect 25123 8756 25181 8757
rect 25123 8716 25132 8756
rect 25172 8716 25181 8756
rect 25123 8715 25181 8716
rect 25411 8756 25469 8757
rect 25411 8716 25420 8756
rect 25460 8716 25469 8756
rect 25411 8715 25469 8716
rect 25603 8756 25661 8757
rect 25603 8716 25612 8756
rect 25652 8716 25661 8756
rect 25603 8715 25661 8716
rect 27427 8756 27485 8757
rect 27427 8716 27436 8756
rect 27476 8716 27485 8756
rect 27427 8715 27485 8716
rect 27627 8756 27669 8765
rect 27627 8716 27628 8756
rect 27668 8716 27669 8756
rect 27627 8707 27669 8716
rect 27819 8756 27861 8765
rect 27819 8716 27820 8756
rect 27860 8716 27861 8756
rect 27819 8707 27861 8716
rect 28003 8756 28061 8757
rect 28003 8716 28012 8756
rect 28052 8716 28061 8756
rect 28003 8715 28061 8716
rect 28203 8756 28245 8765
rect 28203 8716 28204 8756
rect 28244 8716 28245 8756
rect 28203 8707 28245 8716
rect 28387 8756 28445 8757
rect 28387 8716 28396 8756
rect 28436 8716 28445 8756
rect 28387 8715 28445 8716
rect 28587 8756 28629 8765
rect 28587 8716 28588 8756
rect 28628 8716 28629 8756
rect 28587 8707 28629 8716
rect 28771 8756 28829 8757
rect 28771 8716 28780 8756
rect 28820 8716 28829 8756
rect 28771 8715 28829 8716
rect 29347 8756 29405 8757
rect 29347 8716 29356 8756
rect 29396 8716 29405 8756
rect 29347 8715 29405 8716
rect 29539 8756 29597 8757
rect 29539 8716 29548 8756
rect 29588 8716 29597 8756
rect 29539 8715 29597 8716
rect 32331 8756 32373 8765
rect 32331 8716 32332 8756
rect 32372 8716 32373 8756
rect 32331 8707 32373 8716
rect 33963 8756 34005 8765
rect 33963 8716 33964 8756
rect 34004 8716 34005 8756
rect 33963 8707 34005 8716
rect 34155 8756 34197 8765
rect 34155 8716 34156 8756
rect 34196 8716 34197 8756
rect 34155 8707 34197 8716
rect 34347 8756 34389 8765
rect 34347 8716 34348 8756
rect 34388 8716 34389 8756
rect 34347 8707 34389 8716
rect 34531 8756 34589 8757
rect 34531 8716 34540 8756
rect 34580 8716 34589 8756
rect 34531 8715 34589 8716
rect 34731 8756 34773 8765
rect 34731 8716 34732 8756
rect 34772 8716 34773 8756
rect 34731 8707 34773 8716
rect 34915 8756 34973 8757
rect 34915 8716 34924 8756
rect 34964 8716 34973 8756
rect 34915 8715 34973 8716
rect 35115 8756 35157 8765
rect 35115 8716 35116 8756
rect 35156 8716 35157 8756
rect 35115 8707 35157 8716
rect 35299 8756 35357 8757
rect 35299 8716 35308 8756
rect 35348 8716 35357 8756
rect 35299 8715 35357 8716
rect 35499 8756 35541 8765
rect 35499 8716 35500 8756
rect 35540 8716 35541 8756
rect 35499 8707 35541 8716
rect 35683 8756 35741 8757
rect 35683 8716 35692 8756
rect 35732 8716 35741 8756
rect 35683 8715 35741 8716
rect 37027 8756 37085 8757
rect 37027 8716 37036 8756
rect 37076 8716 37085 8756
rect 37027 8715 37085 8716
rect 37219 8756 37277 8757
rect 37219 8716 37228 8756
rect 37268 8716 37277 8756
rect 37219 8715 37277 8716
rect 38275 8756 38333 8757
rect 38275 8716 38284 8756
rect 38324 8716 38333 8756
rect 38275 8715 38333 8716
rect 38467 8756 38525 8757
rect 38467 8716 38476 8756
rect 38516 8716 38525 8756
rect 38467 8715 38525 8716
rect 43363 8756 43421 8757
rect 43363 8716 43372 8756
rect 43412 8716 43421 8756
rect 43363 8715 43421 8716
rect 43651 8756 43709 8757
rect 43651 8716 43660 8756
rect 43700 8716 43709 8756
rect 43651 8715 43709 8716
rect 44611 8756 44669 8757
rect 44611 8716 44620 8756
rect 44660 8716 44669 8756
rect 44611 8715 44669 8716
rect 44907 8756 44949 8765
rect 44907 8716 44908 8756
rect 44948 8716 44949 8756
rect 44907 8707 44949 8716
rect 45099 8756 45141 8765
rect 45099 8716 45100 8756
rect 45140 8716 45141 8756
rect 45099 8707 45141 8716
rect 45195 8756 45237 8765
rect 45195 8716 45196 8756
rect 45236 8716 45237 8756
rect 45195 8707 45237 8716
rect 46147 8756 46205 8757
rect 46147 8716 46156 8756
rect 46196 8716 46205 8756
rect 46147 8715 46205 8716
rect 47107 8756 47165 8757
rect 47107 8716 47116 8756
rect 47156 8716 47165 8756
rect 47107 8715 47165 8716
rect 48355 8756 48413 8757
rect 48355 8716 48364 8756
rect 48404 8716 48413 8756
rect 48355 8715 48413 8716
rect 49323 8756 49365 8765
rect 49323 8716 49324 8756
rect 49364 8716 49365 8756
rect 49323 8707 49365 8716
rect 49419 8756 49461 8765
rect 49419 8716 49420 8756
rect 49460 8716 49461 8756
rect 49419 8707 49461 8716
rect 49611 8756 49653 8765
rect 49611 8716 49612 8756
rect 49652 8716 49653 8756
rect 49611 8707 49653 8716
rect 49987 8756 50045 8757
rect 49987 8716 49996 8756
rect 50036 8716 50045 8756
rect 49987 8715 50045 8716
rect 50467 8756 50525 8757
rect 50467 8716 50476 8756
rect 50516 8716 50525 8756
rect 50467 8715 50525 8716
rect 52587 8756 52629 8765
rect 52587 8716 52588 8756
rect 52628 8716 52629 8756
rect 52587 8707 52629 8716
rect 52683 8756 52725 8765
rect 52683 8716 52684 8756
rect 52724 8716 52725 8756
rect 52683 8707 52725 8716
rect 52875 8756 52917 8765
rect 52875 8716 52876 8756
rect 52916 8716 52917 8756
rect 52875 8707 52917 8716
rect 54315 8756 54357 8765
rect 54315 8716 54316 8756
rect 54356 8716 54357 8756
rect 54315 8707 54357 8716
rect 54507 8756 54549 8765
rect 54507 8716 54508 8756
rect 54548 8716 54549 8756
rect 54507 8707 54549 8716
rect 54891 8764 54933 8773
rect 54891 8724 54892 8764
rect 54932 8724 54933 8764
rect 54891 8715 54933 8724
rect 55275 8756 55317 8765
rect 55275 8716 55276 8756
rect 55316 8716 55317 8756
rect 55275 8707 55317 8716
rect 55947 8756 55989 8765
rect 56811 8764 56853 8773
rect 55947 8716 55948 8756
rect 55988 8716 55989 8756
rect 55947 8707 55989 8716
rect 56131 8756 56189 8757
rect 56131 8716 56140 8756
rect 56180 8716 56189 8756
rect 56131 8715 56189 8716
rect 56811 8724 56812 8764
rect 56852 8724 56853 8764
rect 56811 8715 56853 8724
rect 57195 8764 57237 8773
rect 78315 8769 78357 8778
rect 57195 8724 57196 8764
rect 57236 8724 57237 8764
rect 57195 8715 57237 8724
rect 59203 8756 59261 8757
rect 59203 8716 59212 8756
rect 59252 8716 59261 8756
rect 59203 8715 59261 8716
rect 60075 8756 60117 8765
rect 60075 8716 60076 8756
rect 60116 8716 60117 8756
rect 60075 8707 60117 8716
rect 66979 8756 67037 8757
rect 66979 8716 66988 8756
rect 67028 8716 67037 8756
rect 66979 8715 67037 8716
rect 67171 8756 67229 8757
rect 67171 8716 67180 8756
rect 67220 8716 67229 8756
rect 67171 8715 67229 8716
rect 69955 8756 70013 8757
rect 69955 8716 69964 8756
rect 70004 8716 70013 8756
rect 69955 8715 70013 8716
rect 70155 8756 70197 8765
rect 70155 8716 70156 8756
rect 70196 8716 70197 8756
rect 70155 8707 70197 8716
rect 70435 8756 70493 8757
rect 70435 8716 70444 8756
rect 70484 8716 70493 8756
rect 70435 8715 70493 8716
rect 70635 8756 70677 8765
rect 70635 8716 70636 8756
rect 70676 8716 70677 8756
rect 70635 8707 70677 8716
rect 70819 8756 70877 8757
rect 70819 8716 70828 8756
rect 70868 8716 70877 8756
rect 70819 8715 70877 8716
rect 71019 8756 71061 8765
rect 71019 8716 71020 8756
rect 71060 8716 71061 8756
rect 71019 8707 71061 8716
rect 73219 8756 73277 8757
rect 73219 8716 73228 8756
rect 73268 8716 73277 8756
rect 73219 8715 73277 8716
rect 73419 8756 73461 8765
rect 73419 8716 73420 8756
rect 73460 8716 73461 8756
rect 73419 8707 73461 8716
rect 74563 8756 74621 8757
rect 74563 8716 74572 8756
rect 74612 8716 74621 8756
rect 74563 8715 74621 8716
rect 74763 8756 74805 8765
rect 74763 8716 74764 8756
rect 74804 8716 74805 8756
rect 74763 8707 74805 8716
rect 74947 8756 75005 8757
rect 74947 8716 74956 8756
rect 74996 8716 75005 8756
rect 74947 8715 75005 8716
rect 75147 8756 75189 8765
rect 75147 8716 75148 8756
rect 75188 8716 75189 8756
rect 75147 8707 75189 8716
rect 75331 8756 75389 8757
rect 75331 8716 75340 8756
rect 75380 8716 75389 8756
rect 75331 8715 75389 8716
rect 75531 8756 75573 8765
rect 75531 8716 75532 8756
rect 75572 8716 75573 8756
rect 75531 8707 75573 8716
rect 75907 8756 75965 8757
rect 75907 8716 75916 8756
rect 75956 8716 75965 8756
rect 75907 8715 75965 8716
rect 76099 8756 76157 8757
rect 76099 8716 76108 8756
rect 76148 8716 76157 8756
rect 76099 8715 76157 8716
rect 76683 8756 76725 8765
rect 76683 8716 76684 8756
rect 76724 8716 76725 8756
rect 76683 8707 76725 8716
rect 76867 8756 76925 8757
rect 76867 8716 76876 8756
rect 76916 8716 76925 8756
rect 76867 8715 76925 8716
rect 77931 8756 77973 8765
rect 77931 8716 77932 8756
rect 77972 8716 77973 8756
rect 77931 8707 77973 8716
rect 78115 8756 78173 8757
rect 78115 8716 78124 8756
rect 78164 8716 78173 8756
rect 78315 8729 78316 8769
rect 78356 8729 78357 8769
rect 88203 8769 88245 8778
rect 78315 8720 78357 8729
rect 78499 8756 78557 8757
rect 78115 8715 78173 8716
rect 78499 8716 78508 8756
rect 78548 8716 78557 8756
rect 78499 8715 78557 8716
rect 78691 8756 78749 8757
rect 78691 8716 78700 8756
rect 78740 8716 78749 8756
rect 78691 8715 78749 8716
rect 78891 8756 78933 8765
rect 78891 8716 78892 8756
rect 78932 8716 78933 8756
rect 78891 8707 78933 8716
rect 80811 8756 80853 8765
rect 80811 8716 80812 8756
rect 80852 8716 80853 8756
rect 80811 8707 80853 8716
rect 80995 8756 81053 8757
rect 80995 8716 81004 8756
rect 81044 8716 81053 8756
rect 80995 8715 81053 8716
rect 81195 8756 81237 8765
rect 81195 8716 81196 8756
rect 81236 8716 81237 8756
rect 81195 8707 81237 8716
rect 81291 8756 81333 8765
rect 81291 8716 81292 8756
rect 81332 8716 81333 8756
rect 81291 8707 81333 8716
rect 81379 8756 81437 8757
rect 81379 8716 81388 8756
rect 81428 8716 81437 8756
rect 81379 8715 81437 8716
rect 81579 8756 81621 8765
rect 81579 8716 81580 8756
rect 81620 8716 81621 8756
rect 81579 8707 81621 8716
rect 81763 8756 81821 8757
rect 81763 8716 81772 8756
rect 81812 8716 81821 8756
rect 81763 8715 81821 8716
rect 81963 8756 82005 8765
rect 81963 8716 81964 8756
rect 82004 8716 82005 8756
rect 81963 8707 82005 8716
rect 82147 8756 82205 8757
rect 82147 8716 82156 8756
rect 82196 8716 82205 8756
rect 82147 8715 82205 8716
rect 83115 8756 83157 8765
rect 83115 8716 83116 8756
rect 83156 8716 83157 8756
rect 83115 8707 83157 8716
rect 83299 8756 83357 8757
rect 83299 8716 83308 8756
rect 83348 8716 83357 8756
rect 83299 8715 83357 8716
rect 83499 8756 83541 8765
rect 83499 8716 83500 8756
rect 83540 8716 83541 8756
rect 83499 8707 83541 8716
rect 83683 8756 83741 8757
rect 83683 8716 83692 8756
rect 83732 8716 83741 8756
rect 83683 8715 83741 8716
rect 84075 8756 84117 8765
rect 84075 8716 84076 8756
rect 84116 8716 84117 8756
rect 84075 8707 84117 8716
rect 84259 8756 84317 8757
rect 84259 8716 84268 8756
rect 84308 8716 84317 8756
rect 84259 8715 84317 8716
rect 86851 8756 86909 8757
rect 86851 8716 86860 8756
rect 86900 8716 86909 8756
rect 86851 8715 86909 8716
rect 87051 8756 87093 8765
rect 87051 8716 87052 8756
rect 87092 8716 87093 8756
rect 87051 8707 87093 8716
rect 87235 8756 87293 8757
rect 87235 8716 87244 8756
rect 87284 8716 87293 8756
rect 87235 8715 87293 8716
rect 87435 8756 87477 8765
rect 87435 8716 87436 8756
rect 87476 8716 87477 8756
rect 87435 8707 87477 8716
rect 87619 8756 87677 8757
rect 87619 8716 87628 8756
rect 87668 8716 87677 8756
rect 87619 8715 87677 8716
rect 87819 8756 87861 8765
rect 87819 8716 87820 8756
rect 87860 8716 87861 8756
rect 87819 8707 87861 8716
rect 88003 8756 88061 8757
rect 88003 8716 88012 8756
rect 88052 8716 88061 8756
rect 88203 8729 88204 8769
rect 88244 8729 88245 8769
rect 88203 8720 88245 8729
rect 88971 8756 89013 8765
rect 88003 8715 88061 8716
rect 88971 8716 88972 8756
rect 89012 8716 89013 8756
rect 88971 8707 89013 8716
rect 89155 8756 89213 8757
rect 89155 8716 89164 8756
rect 89204 8716 89213 8756
rect 89155 8715 89213 8716
rect 89355 8756 89397 8765
rect 89355 8716 89356 8756
rect 89396 8716 89397 8756
rect 89355 8707 89397 8716
rect 89539 8756 89597 8757
rect 89539 8716 89548 8756
rect 89588 8716 89597 8756
rect 89539 8715 89597 8716
rect 34059 8672 34101 8681
rect 34059 8632 34060 8672
rect 34100 8632 34101 8672
rect 34059 8623 34101 8632
rect 42507 8672 42549 8681
rect 42507 8632 42508 8672
rect 42548 8632 42549 8672
rect 42507 8623 42549 8632
rect 48739 8672 48797 8673
rect 48739 8632 48748 8672
rect 48788 8632 48797 8672
rect 48739 8631 48797 8632
rect 54411 8672 54453 8681
rect 54411 8632 54412 8672
rect 54452 8632 54453 8672
rect 54411 8623 54453 8632
rect 58915 8672 58973 8673
rect 58915 8632 58924 8672
rect 58964 8632 58973 8672
rect 58915 8631 58973 8632
rect 48075 8588 48117 8597
rect 48075 8548 48076 8588
rect 48116 8548 48117 8588
rect 48075 8539 48117 8548
rect 48939 8588 48981 8597
rect 48939 8548 48940 8588
rect 48980 8548 48981 8588
rect 48939 8539 48981 8548
rect 54891 8588 54933 8597
rect 54891 8548 54892 8588
rect 54932 8548 54933 8588
rect 54891 8539 54933 8548
rect 55275 8588 55317 8597
rect 55275 8548 55276 8588
rect 55316 8548 55317 8588
rect 55275 8539 55317 8548
rect 56043 8588 56085 8597
rect 56043 8548 56044 8588
rect 56084 8548 56085 8588
rect 56043 8539 56085 8548
rect 56619 8588 56661 8597
rect 56619 8548 56620 8588
rect 56660 8548 56661 8588
rect 56619 8539 56661 8548
rect 56811 8588 56853 8597
rect 56811 8548 56812 8588
rect 56852 8548 56853 8588
rect 56811 8539 56853 8548
rect 57195 8588 57237 8597
rect 57195 8548 57196 8588
rect 57236 8548 57237 8588
rect 57195 8539 57237 8548
rect 84171 8588 84213 8597
rect 84171 8548 84172 8588
rect 84212 8548 84213 8588
rect 84171 8539 84213 8548
rect 10155 8504 10197 8513
rect 10155 8464 10156 8504
rect 10196 8464 10197 8504
rect 10155 8455 10197 8464
rect 11211 8504 11253 8513
rect 11211 8464 11212 8504
rect 11252 8464 11253 8504
rect 11211 8455 11253 8464
rect 24267 8504 24309 8513
rect 24267 8464 24268 8504
rect 24308 8464 24309 8504
rect 24267 8455 24309 8464
rect 24651 8504 24693 8513
rect 24651 8464 24652 8504
rect 24692 8464 24693 8504
rect 24651 8455 24693 8464
rect 27531 8504 27573 8513
rect 27531 8464 27532 8504
rect 27572 8464 27573 8504
rect 27531 8455 27573 8464
rect 34443 8504 34485 8513
rect 34443 8464 34444 8504
rect 34484 8464 34485 8504
rect 34443 8455 34485 8464
rect 35211 8504 35253 8513
rect 35211 8464 35212 8504
rect 35252 8464 35253 8504
rect 35211 8455 35253 8464
rect 35595 8504 35637 8513
rect 35595 8464 35596 8504
rect 35636 8464 35637 8504
rect 35595 8455 35637 8464
rect 50955 8504 50997 8513
rect 50955 8464 50956 8504
rect 50996 8464 50997 8504
rect 50955 8455 50997 8464
rect 54699 8504 54741 8513
rect 54699 8464 54700 8504
rect 54740 8464 54741 8504
rect 54699 8455 54741 8464
rect 57387 8504 57429 8513
rect 57387 8464 57388 8504
rect 57428 8464 57429 8504
rect 57387 8455 57429 8464
rect 73323 8504 73365 8513
rect 73323 8464 73324 8504
rect 73364 8464 73365 8504
rect 73323 8455 73365 8464
rect 76779 8504 76821 8513
rect 76779 8464 76780 8504
rect 76820 8464 76821 8504
rect 76779 8455 76821 8464
rect 78027 8504 78069 8513
rect 78027 8464 78028 8504
rect 78068 8464 78069 8504
rect 78027 8455 78069 8464
rect 78411 8504 78453 8513
rect 78411 8464 78412 8504
rect 78452 8464 78453 8504
rect 78411 8455 78453 8464
rect 87339 8504 87381 8513
rect 87339 8464 87340 8504
rect 87380 8464 87381 8504
rect 87339 8455 87381 8464
rect 88107 8504 88149 8513
rect 88107 8464 88108 8504
rect 88148 8464 88149 8504
rect 88107 8455 88149 8464
rect 89451 8504 89493 8513
rect 89451 8464 89452 8504
rect 89492 8464 89493 8504
rect 89451 8455 89493 8464
rect 1152 8336 98784 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 64168 8336
rect 64208 8296 64250 8336
rect 64290 8296 64332 8336
rect 64372 8296 64414 8336
rect 64454 8296 64496 8336
rect 64536 8296 79288 8336
rect 79328 8296 79370 8336
rect 79410 8296 79452 8336
rect 79492 8296 79534 8336
rect 79574 8296 79616 8336
rect 79656 8296 94408 8336
rect 94448 8296 94490 8336
rect 94530 8296 94572 8336
rect 94612 8296 94654 8336
rect 94694 8296 94736 8336
rect 94776 8296 98784 8336
rect 1152 8272 98784 8296
rect 30219 8168 30261 8177
rect 30219 8128 30220 8168
rect 30260 8128 30261 8168
rect 30219 8119 30261 8128
rect 37035 8168 37077 8177
rect 37035 8128 37036 8168
rect 37076 8128 37077 8168
rect 37035 8119 37077 8128
rect 50763 8168 50805 8177
rect 50763 8128 50764 8168
rect 50804 8128 50805 8168
rect 50763 8119 50805 8128
rect 54603 8168 54645 8177
rect 54603 8128 54604 8168
rect 54644 8128 54645 8168
rect 54603 8119 54645 8128
rect 58731 8168 58773 8177
rect 58731 8128 58732 8168
rect 58772 8128 58773 8168
rect 58731 8119 58773 8128
rect 60171 8168 60213 8177
rect 60171 8128 60172 8168
rect 60212 8128 60213 8168
rect 60171 8119 60213 8128
rect 72547 8168 72605 8169
rect 72547 8128 72556 8168
rect 72596 8128 72605 8168
rect 72547 8127 72605 8128
rect 75043 8168 75101 8169
rect 75043 8128 75052 8168
rect 75092 8128 75101 8168
rect 75043 8127 75101 8128
rect 81579 8168 81621 8177
rect 81579 8128 81580 8168
rect 81620 8128 81621 8168
rect 81579 8119 81621 8128
rect 83691 8168 83733 8177
rect 83691 8128 83692 8168
rect 83732 8128 83733 8168
rect 83691 8119 83733 8128
rect 86955 8168 86997 8177
rect 86955 8128 86956 8168
rect 86996 8128 86997 8168
rect 86955 8119 86997 8128
rect 12459 8084 12501 8093
rect 12459 8044 12460 8084
rect 12500 8044 12501 8084
rect 12459 8035 12501 8044
rect 22347 8084 22389 8093
rect 22347 8044 22348 8084
rect 22388 8044 22389 8084
rect 22347 8035 22389 8044
rect 37707 8084 37749 8093
rect 37707 8044 37708 8084
rect 37748 8044 37749 8084
rect 37707 8035 37749 8044
rect 46251 8084 46293 8093
rect 46251 8044 46252 8084
rect 46292 8044 46293 8084
rect 46251 8035 46293 8044
rect 48171 8084 48213 8093
rect 48171 8044 48172 8084
rect 48212 8044 48213 8084
rect 48171 8035 48213 8044
rect 51435 8084 51477 8093
rect 51435 8044 51436 8084
rect 51476 8044 51477 8084
rect 51435 8035 51477 8044
rect 58923 8084 58965 8093
rect 58923 8044 58924 8084
rect 58964 8044 58965 8084
rect 58923 8035 58965 8044
rect 85227 8084 85269 8093
rect 85227 8044 85228 8084
rect 85268 8044 85269 8084
rect 85227 8035 85269 8044
rect 16299 8000 16341 8009
rect 16299 7960 16300 8000
rect 16340 7960 16341 8000
rect 16299 7951 16341 7960
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 34923 8000 34965 8009
rect 34923 7960 34924 8000
rect 34964 7960 34965 8000
rect 34923 7951 34965 7960
rect 35307 8000 35349 8009
rect 35307 7960 35308 8000
rect 35348 7960 35349 8000
rect 35307 7951 35349 7960
rect 45579 8000 45621 8009
rect 45579 7960 45580 8000
rect 45620 7960 45621 8000
rect 45579 7951 45621 7960
rect 50563 8000 50621 8001
rect 50563 7960 50572 8000
rect 50612 7960 50621 8000
rect 50563 7959 50621 7960
rect 54403 8000 54461 8001
rect 54403 7960 54412 8000
rect 54452 7960 54461 8000
rect 54403 7959 54461 7960
rect 58347 8000 58389 8009
rect 58347 7960 58348 8000
rect 58388 7960 58389 8000
rect 58347 7951 58389 7960
rect 59971 8000 60029 8001
rect 59971 7960 59980 8000
rect 60020 7960 60029 8000
rect 59971 7959 60029 7960
rect 84843 8000 84885 8009
rect 84843 7960 84844 8000
rect 84884 7960 84885 8000
rect 84843 7951 84885 7960
rect 87531 8000 87573 8009
rect 87531 7960 87532 8000
rect 87572 7960 87573 8000
rect 87531 7951 87573 7960
rect 82435 7939 82493 7940
rect 8907 7916 8949 7925
rect 8907 7876 8908 7916
rect 8948 7876 8949 7916
rect 8907 7867 8949 7876
rect 9091 7916 9149 7917
rect 9091 7876 9100 7916
rect 9140 7876 9149 7916
rect 9091 7875 9149 7876
rect 9291 7916 9333 7925
rect 9291 7876 9292 7916
rect 9332 7876 9333 7916
rect 9291 7867 9333 7876
rect 9475 7916 9533 7917
rect 9475 7876 9484 7916
rect 9524 7876 9533 7916
rect 9475 7875 9533 7876
rect 9667 7916 9725 7917
rect 9667 7876 9676 7916
rect 9716 7876 9725 7916
rect 9667 7875 9725 7876
rect 9867 7916 9909 7925
rect 9867 7876 9868 7916
rect 9908 7876 9909 7916
rect 9867 7867 9909 7876
rect 10051 7916 10109 7917
rect 10051 7876 10060 7916
rect 10100 7876 10109 7916
rect 10051 7875 10109 7876
rect 10251 7916 10293 7925
rect 10251 7876 10252 7916
rect 10292 7876 10293 7916
rect 10251 7867 10293 7876
rect 10435 7916 10493 7917
rect 10435 7876 10444 7916
rect 10484 7876 10493 7916
rect 10435 7875 10493 7876
rect 10635 7916 10677 7925
rect 10635 7876 10636 7916
rect 10676 7876 10677 7916
rect 10635 7867 10677 7876
rect 11587 7916 11645 7917
rect 11587 7876 11596 7916
rect 11636 7876 11645 7916
rect 11587 7875 11645 7876
rect 11787 7916 11829 7925
rect 11787 7876 11788 7916
rect 11828 7876 11829 7916
rect 11787 7867 11829 7876
rect 11979 7916 12021 7925
rect 11979 7876 11980 7916
rect 12020 7876 12021 7916
rect 11979 7867 12021 7876
rect 12163 7916 12221 7917
rect 12163 7876 12172 7916
rect 12212 7876 12221 7916
rect 12163 7875 12221 7876
rect 12355 7916 12413 7917
rect 12355 7876 12364 7916
rect 12404 7876 12413 7916
rect 12355 7875 12413 7876
rect 12555 7916 12597 7925
rect 12555 7876 12556 7916
rect 12596 7876 12597 7916
rect 12555 7867 12597 7876
rect 12747 7916 12789 7925
rect 12747 7876 12748 7916
rect 12788 7876 12789 7916
rect 12747 7867 12789 7876
rect 12931 7916 12989 7917
rect 12931 7876 12940 7916
rect 12980 7876 12989 7916
rect 12931 7875 12989 7876
rect 13131 7916 13173 7925
rect 13131 7876 13132 7916
rect 13172 7876 13173 7916
rect 13131 7867 13173 7876
rect 13315 7916 13373 7917
rect 13315 7876 13324 7916
rect 13364 7876 13373 7916
rect 13315 7875 13373 7876
rect 13515 7916 13557 7925
rect 13515 7876 13516 7916
rect 13556 7876 13557 7916
rect 13515 7867 13557 7876
rect 13699 7916 13757 7917
rect 13699 7876 13708 7916
rect 13748 7876 13757 7916
rect 13699 7875 13757 7876
rect 14179 7916 14237 7917
rect 14179 7876 14188 7916
rect 14228 7876 14237 7916
rect 14179 7875 14237 7876
rect 14371 7916 14429 7917
rect 14371 7876 14380 7916
rect 14420 7876 14429 7916
rect 14371 7875 14429 7876
rect 17155 7916 17213 7917
rect 17155 7876 17164 7916
rect 17204 7876 17213 7916
rect 17155 7875 17213 7876
rect 17827 7916 17885 7917
rect 17827 7876 17836 7916
rect 17876 7876 17885 7916
rect 17827 7875 17885 7876
rect 18027 7916 18069 7925
rect 18027 7876 18028 7916
rect 18068 7876 18069 7916
rect 18027 7867 18069 7876
rect 18219 7916 18261 7925
rect 18219 7876 18220 7916
rect 18260 7876 18261 7916
rect 18219 7867 18261 7876
rect 18403 7916 18461 7917
rect 18403 7876 18412 7916
rect 18452 7876 18461 7916
rect 18403 7875 18461 7876
rect 18603 7916 18645 7925
rect 18603 7876 18604 7916
rect 18644 7876 18645 7916
rect 18603 7867 18645 7876
rect 18787 7916 18845 7917
rect 18787 7876 18796 7916
rect 18836 7876 18845 7916
rect 18787 7875 18845 7876
rect 18987 7916 19029 7925
rect 18987 7876 18988 7916
rect 19028 7876 19029 7916
rect 18987 7867 19029 7876
rect 19171 7916 19229 7917
rect 19171 7876 19180 7916
rect 19220 7876 19229 7916
rect 19171 7875 19229 7876
rect 19371 7916 19413 7925
rect 19371 7876 19372 7916
rect 19412 7876 19413 7916
rect 19371 7867 19413 7876
rect 19555 7916 19613 7917
rect 19555 7876 19564 7916
rect 19604 7876 19613 7916
rect 19555 7875 19613 7876
rect 19747 7916 19805 7917
rect 19747 7876 19756 7916
rect 19796 7876 19805 7916
rect 20419 7916 20477 7917
rect 19747 7875 19805 7876
rect 19947 7903 19989 7912
rect 19947 7863 19948 7903
rect 19988 7863 19989 7903
rect 20419 7876 20428 7916
rect 20468 7876 20477 7916
rect 20419 7875 20477 7876
rect 20611 7916 20669 7917
rect 20611 7876 20620 7916
rect 20660 7876 20669 7916
rect 20611 7875 20669 7876
rect 22539 7916 22581 7925
rect 22539 7876 22540 7916
rect 22580 7876 22581 7916
rect 22539 7867 22581 7876
rect 22635 7916 22677 7925
rect 22635 7876 22636 7916
rect 22676 7876 22677 7916
rect 22635 7867 22677 7876
rect 23211 7916 23253 7925
rect 23211 7876 23212 7916
rect 23252 7876 23253 7916
rect 23211 7867 23253 7876
rect 23307 7916 23349 7925
rect 23307 7876 23308 7916
rect 23348 7876 23349 7916
rect 23307 7867 23349 7876
rect 24547 7916 24605 7917
rect 24547 7876 24556 7916
rect 24596 7876 24605 7916
rect 24547 7875 24605 7876
rect 24747 7916 24789 7925
rect 24747 7876 24748 7916
rect 24788 7876 24789 7916
rect 24747 7867 24789 7876
rect 24939 7916 24981 7925
rect 24939 7876 24940 7916
rect 24980 7876 24981 7916
rect 24939 7867 24981 7876
rect 25123 7916 25181 7917
rect 25123 7876 25132 7916
rect 25172 7876 25181 7916
rect 25123 7875 25181 7876
rect 25315 7916 25373 7917
rect 25315 7876 25324 7916
rect 25364 7876 25373 7916
rect 25315 7875 25373 7876
rect 25515 7916 25557 7925
rect 25515 7876 25516 7916
rect 25556 7876 25557 7916
rect 25515 7867 25557 7876
rect 25707 7916 25749 7925
rect 25707 7876 25708 7916
rect 25748 7876 25749 7916
rect 25707 7867 25749 7876
rect 25891 7916 25949 7917
rect 25891 7876 25900 7916
rect 25940 7876 25949 7916
rect 25891 7875 25949 7876
rect 27627 7916 27669 7925
rect 27627 7876 27628 7916
rect 27668 7876 27669 7916
rect 27627 7867 27669 7876
rect 27811 7916 27869 7917
rect 27811 7876 27820 7916
rect 27860 7876 27869 7916
rect 27811 7875 27869 7876
rect 28011 7916 28053 7925
rect 28011 7876 28012 7916
rect 28052 7876 28053 7916
rect 28011 7867 28053 7876
rect 28195 7916 28253 7917
rect 28195 7876 28204 7916
rect 28244 7876 28253 7916
rect 28195 7875 28253 7876
rect 28395 7916 28437 7925
rect 28395 7876 28396 7916
rect 28436 7876 28437 7916
rect 28395 7867 28437 7876
rect 28579 7916 28637 7917
rect 28579 7876 28588 7916
rect 28628 7876 28637 7916
rect 28579 7875 28637 7876
rect 28779 7916 28821 7925
rect 28779 7876 28780 7916
rect 28820 7876 28821 7916
rect 28779 7867 28821 7876
rect 28963 7916 29021 7917
rect 28963 7876 28972 7916
rect 29012 7876 29021 7916
rect 28963 7875 29021 7876
rect 29931 7916 29973 7925
rect 29931 7876 29932 7916
rect 29972 7876 29973 7916
rect 29931 7867 29973 7876
rect 30027 7916 30069 7925
rect 30027 7876 30028 7916
rect 30068 7876 30069 7916
rect 30027 7867 30069 7876
rect 30787 7916 30845 7917
rect 30787 7876 30796 7916
rect 30836 7876 30845 7916
rect 30787 7875 30845 7876
rect 30987 7916 31029 7925
rect 30987 7876 30988 7916
rect 31028 7876 31029 7916
rect 30987 7867 31029 7876
rect 31179 7916 31221 7925
rect 31179 7876 31180 7916
rect 31220 7876 31221 7916
rect 31179 7867 31221 7876
rect 31363 7916 31421 7917
rect 31363 7876 31372 7916
rect 31412 7876 31421 7916
rect 31363 7875 31421 7876
rect 31563 7916 31605 7925
rect 31563 7876 31564 7916
rect 31604 7876 31605 7916
rect 31563 7867 31605 7876
rect 31747 7916 31805 7917
rect 31747 7876 31756 7916
rect 31796 7876 31805 7916
rect 31747 7875 31805 7876
rect 31947 7916 31989 7925
rect 31947 7876 31948 7916
rect 31988 7876 31989 7916
rect 31947 7867 31989 7876
rect 32131 7916 32189 7917
rect 32131 7876 32140 7916
rect 32180 7876 32189 7916
rect 32131 7875 32189 7876
rect 32331 7916 32373 7925
rect 32331 7876 32332 7916
rect 32372 7876 32373 7916
rect 32331 7867 32373 7876
rect 32515 7916 32573 7917
rect 32515 7876 32524 7916
rect 32564 7876 32573 7916
rect 32515 7875 32573 7876
rect 32715 7916 32757 7925
rect 32715 7876 32716 7916
rect 32756 7876 32757 7916
rect 32715 7867 32757 7876
rect 32811 7916 32853 7925
rect 32811 7876 32812 7916
rect 32852 7876 32853 7916
rect 32811 7867 32853 7876
rect 32899 7916 32957 7917
rect 32899 7876 32908 7916
rect 32948 7876 32957 7916
rect 32899 7875 32957 7876
rect 33099 7916 33141 7925
rect 33099 7876 33100 7916
rect 33140 7876 33141 7916
rect 33099 7867 33141 7876
rect 33195 7916 33237 7925
rect 33195 7876 33196 7916
rect 33236 7876 33237 7916
rect 33195 7867 33237 7876
rect 33283 7916 33341 7917
rect 33283 7876 33292 7916
rect 33332 7876 33341 7916
rect 33283 7875 33341 7876
rect 33571 7916 33629 7917
rect 33571 7876 33580 7916
rect 33620 7876 33629 7916
rect 33571 7875 33629 7876
rect 33763 7916 33821 7917
rect 33763 7876 33772 7916
rect 33812 7876 33821 7916
rect 33763 7875 33821 7876
rect 34443 7916 34485 7925
rect 34443 7876 34444 7916
rect 34484 7876 34485 7916
rect 34443 7867 34485 7876
rect 34627 7916 34685 7917
rect 34627 7876 34636 7916
rect 34676 7876 34685 7916
rect 34627 7875 34685 7876
rect 34827 7916 34869 7925
rect 34827 7876 34828 7916
rect 34868 7876 34869 7916
rect 34827 7867 34869 7876
rect 35011 7916 35069 7917
rect 35011 7876 35020 7916
rect 35060 7876 35069 7916
rect 35011 7875 35069 7876
rect 36163 7916 36221 7917
rect 36163 7876 36172 7916
rect 36212 7876 36221 7916
rect 36163 7875 36221 7876
rect 36747 7916 36789 7925
rect 36747 7876 36748 7916
rect 36788 7876 36789 7916
rect 36747 7867 36789 7876
rect 37419 7916 37461 7925
rect 37419 7876 37420 7916
rect 37460 7876 37461 7916
rect 36835 7874 36893 7875
rect 19947 7854 19989 7863
rect 9003 7832 9045 7841
rect 9003 7792 9004 7832
rect 9044 7792 9045 7832
rect 9003 7783 9045 7792
rect 9387 7832 9429 7841
rect 9387 7792 9388 7832
rect 9428 7792 9429 7832
rect 9387 7783 9429 7792
rect 9771 7832 9813 7841
rect 9771 7792 9772 7832
rect 9812 7792 9813 7832
rect 9771 7783 9813 7792
rect 10155 7832 10197 7841
rect 10155 7792 10156 7832
rect 10196 7792 10197 7832
rect 10155 7783 10197 7792
rect 10539 7832 10581 7841
rect 10539 7792 10540 7832
rect 10580 7792 10581 7832
rect 10539 7783 10581 7792
rect 11691 7832 11733 7841
rect 11691 7792 11692 7832
rect 11732 7792 11733 7832
rect 11691 7783 11733 7792
rect 12075 7832 12117 7841
rect 12075 7792 12076 7832
rect 12116 7792 12117 7832
rect 12075 7783 12117 7792
rect 12843 7832 12885 7841
rect 12843 7792 12844 7832
rect 12884 7792 12885 7832
rect 12843 7783 12885 7792
rect 13227 7832 13269 7841
rect 13227 7792 13228 7832
rect 13268 7792 13269 7832
rect 13227 7783 13269 7792
rect 13611 7832 13653 7841
rect 13611 7792 13612 7832
rect 13652 7792 13653 7832
rect 13611 7783 13653 7792
rect 17931 7832 17973 7841
rect 17931 7792 17932 7832
rect 17972 7792 17973 7832
rect 17931 7783 17973 7792
rect 18315 7832 18357 7841
rect 18315 7792 18316 7832
rect 18356 7792 18357 7832
rect 18315 7783 18357 7792
rect 18699 7832 18741 7841
rect 18699 7792 18700 7832
rect 18740 7792 18741 7832
rect 18699 7783 18741 7792
rect 19083 7832 19125 7841
rect 19083 7792 19084 7832
rect 19124 7792 19125 7832
rect 19083 7783 19125 7792
rect 19467 7832 19509 7841
rect 19467 7792 19468 7832
rect 19508 7792 19509 7832
rect 19467 7783 19509 7792
rect 19851 7832 19893 7841
rect 19851 7792 19852 7832
rect 19892 7792 19893 7832
rect 19851 7783 19893 7792
rect 23011 7832 23069 7833
rect 23011 7792 23020 7832
rect 23060 7792 23069 7832
rect 23011 7791 23069 7792
rect 24651 7832 24693 7841
rect 24651 7792 24652 7832
rect 24692 7792 24693 7832
rect 24651 7783 24693 7792
rect 25035 7832 25077 7841
rect 25035 7792 25036 7832
rect 25076 7792 25077 7832
rect 25035 7783 25077 7792
rect 25419 7832 25461 7841
rect 25419 7792 25420 7832
rect 25460 7792 25461 7832
rect 25419 7783 25461 7792
rect 25803 7832 25845 7841
rect 25803 7792 25804 7832
rect 25844 7792 25845 7832
rect 25803 7783 25845 7792
rect 27723 7832 27765 7841
rect 27723 7792 27724 7832
rect 27764 7792 27765 7832
rect 27723 7783 27765 7792
rect 28107 7832 28149 7841
rect 28107 7792 28108 7832
rect 28148 7792 28149 7832
rect 28107 7783 28149 7792
rect 28491 7832 28533 7841
rect 28491 7792 28492 7832
rect 28532 7792 28533 7832
rect 28491 7783 28533 7792
rect 28875 7832 28917 7841
rect 28875 7792 28876 7832
rect 28916 7792 28917 7832
rect 28875 7783 28917 7792
rect 30891 7832 30933 7841
rect 30891 7792 30892 7832
rect 30932 7792 30933 7832
rect 30891 7783 30933 7792
rect 31275 7832 31317 7841
rect 31275 7792 31276 7832
rect 31316 7792 31317 7832
rect 31275 7783 31317 7792
rect 31659 7832 31701 7841
rect 31659 7792 31660 7832
rect 31700 7792 31701 7832
rect 31659 7783 31701 7792
rect 32043 7832 32085 7841
rect 32043 7792 32044 7832
rect 32084 7792 32085 7832
rect 32043 7783 32085 7792
rect 34539 7832 34581 7841
rect 36835 7834 36844 7874
rect 36884 7834 36893 7874
rect 37419 7867 37461 7876
rect 37515 7916 37557 7925
rect 37515 7876 37516 7916
rect 37556 7876 37557 7916
rect 37515 7867 37557 7876
rect 39427 7916 39485 7917
rect 39427 7876 39436 7916
rect 39476 7876 39485 7916
rect 39427 7875 39485 7876
rect 39531 7916 39573 7925
rect 39531 7876 39532 7916
rect 39572 7876 39573 7916
rect 39531 7867 39573 7876
rect 39715 7916 39773 7917
rect 39715 7876 39724 7916
rect 39764 7876 39773 7916
rect 39715 7875 39773 7876
rect 39907 7916 39965 7917
rect 39907 7876 39916 7916
rect 39956 7876 39965 7916
rect 39907 7875 39965 7876
rect 40867 7916 40925 7917
rect 40867 7876 40876 7916
rect 40916 7876 40925 7916
rect 40867 7875 40925 7876
rect 41155 7916 41213 7917
rect 41155 7876 41164 7916
rect 41204 7876 41213 7916
rect 41155 7875 41213 7876
rect 42027 7916 42069 7925
rect 42027 7876 42028 7916
rect 42068 7876 42069 7916
rect 42027 7867 42069 7876
rect 42403 7916 42461 7917
rect 42403 7876 42412 7916
rect 42452 7876 42461 7916
rect 42403 7875 42461 7876
rect 43363 7916 43421 7917
rect 43363 7876 43372 7916
rect 43412 7876 43421 7916
rect 43363 7875 43421 7876
rect 44043 7916 44085 7925
rect 44043 7876 44044 7916
rect 44084 7876 44085 7916
rect 44043 7867 44085 7876
rect 44235 7916 44277 7925
rect 44235 7876 44236 7916
rect 44276 7876 44277 7916
rect 44235 7867 44277 7876
rect 44331 7916 44373 7925
rect 44331 7876 44332 7916
rect 44372 7876 44373 7916
rect 44331 7867 44373 7876
rect 44907 7916 44949 7925
rect 44907 7876 44908 7916
rect 44948 7876 44949 7916
rect 44907 7867 44949 7876
rect 45003 7916 45045 7925
rect 45003 7876 45004 7916
rect 45044 7876 45045 7916
rect 45003 7867 45045 7876
rect 45195 7916 45237 7925
rect 45195 7876 45196 7916
rect 45236 7876 45237 7916
rect 45195 7867 45237 7876
rect 45771 7916 45813 7925
rect 45771 7876 45772 7916
rect 45812 7876 45813 7916
rect 45771 7867 45813 7876
rect 45867 7916 45909 7925
rect 45867 7876 45868 7916
rect 45908 7876 45909 7916
rect 45867 7867 45909 7876
rect 46443 7916 46485 7925
rect 46443 7876 46444 7916
rect 46484 7876 46485 7916
rect 46443 7867 46485 7876
rect 46539 7916 46581 7925
rect 46539 7876 46540 7916
rect 46580 7876 46581 7916
rect 46539 7867 46581 7876
rect 46923 7916 46965 7925
rect 46923 7876 46924 7916
rect 46964 7876 46965 7916
rect 46923 7867 46965 7876
rect 47115 7916 47157 7925
rect 47115 7876 47116 7916
rect 47156 7876 47157 7916
rect 47115 7867 47157 7876
rect 47211 7916 47253 7925
rect 47211 7876 47212 7916
rect 47252 7876 47253 7916
rect 47211 7867 47253 7876
rect 48363 7916 48405 7925
rect 48363 7876 48364 7916
rect 48404 7876 48405 7916
rect 48363 7867 48405 7876
rect 48459 7916 48501 7925
rect 48459 7876 48460 7916
rect 48500 7876 48501 7916
rect 48459 7867 48501 7876
rect 49219 7916 49277 7917
rect 49219 7876 49228 7916
rect 49268 7876 49277 7916
rect 49219 7875 49277 7876
rect 50179 7916 50237 7917
rect 50179 7876 50188 7916
rect 50228 7876 50237 7916
rect 50179 7875 50237 7876
rect 51243 7916 51285 7925
rect 51243 7876 51244 7916
rect 51284 7876 51285 7916
rect 51243 7867 51285 7876
rect 51435 7916 51477 7925
rect 51435 7876 51436 7916
rect 51476 7876 51477 7916
rect 51435 7867 51477 7876
rect 51619 7916 51677 7917
rect 51619 7876 51628 7916
rect 51668 7876 51677 7916
rect 51619 7875 51677 7876
rect 51811 7916 51869 7917
rect 51811 7876 51820 7916
rect 51860 7876 51869 7916
rect 51811 7875 51869 7876
rect 54795 7916 54837 7925
rect 54795 7876 54796 7916
rect 54836 7876 54837 7916
rect 54795 7867 54837 7876
rect 54987 7916 55029 7925
rect 54987 7876 54988 7916
rect 55028 7876 55029 7916
rect 54987 7867 55029 7876
rect 56043 7916 56085 7925
rect 56043 7876 56044 7916
rect 56084 7876 56085 7916
rect 56043 7867 56085 7876
rect 56139 7916 56181 7925
rect 56139 7876 56140 7916
rect 56180 7876 56181 7916
rect 56139 7867 56181 7876
rect 56227 7916 56285 7917
rect 56227 7876 56236 7916
rect 56276 7876 56285 7916
rect 56227 7875 56285 7876
rect 56427 7916 56469 7925
rect 56427 7876 56428 7916
rect 56468 7876 56469 7916
rect 56427 7867 56469 7876
rect 56619 7916 56661 7925
rect 56619 7876 56620 7916
rect 56660 7876 56661 7916
rect 56619 7867 56661 7876
rect 56811 7916 56853 7925
rect 56811 7876 56812 7916
rect 56852 7876 56853 7916
rect 56811 7867 56853 7876
rect 57003 7916 57045 7925
rect 57003 7876 57004 7916
rect 57044 7876 57045 7916
rect 57003 7867 57045 7876
rect 57675 7916 57717 7925
rect 57675 7876 57676 7916
rect 57716 7876 57717 7916
rect 57675 7867 57717 7876
rect 57867 7916 57909 7925
rect 57867 7876 57868 7916
rect 57908 7876 57909 7916
rect 57867 7867 57909 7876
rect 58251 7916 58293 7925
rect 58251 7876 58252 7916
rect 58292 7876 58293 7916
rect 58251 7867 58293 7876
rect 58443 7916 58485 7925
rect 58443 7876 58444 7916
rect 58484 7876 58485 7916
rect 58443 7867 58485 7876
rect 58923 7916 58965 7925
rect 58923 7876 58924 7916
rect 58964 7876 58965 7916
rect 58923 7867 58965 7876
rect 59491 7916 59549 7917
rect 59491 7876 59500 7916
rect 59540 7876 59549 7916
rect 59491 7875 59549 7876
rect 59683 7916 59741 7917
rect 59683 7876 59692 7916
rect 59732 7876 59741 7916
rect 59683 7875 59741 7876
rect 62659 7916 62717 7917
rect 62659 7876 62668 7916
rect 62708 7876 62717 7916
rect 62659 7875 62717 7876
rect 63619 7916 63677 7917
rect 63619 7876 63628 7916
rect 63668 7876 63677 7916
rect 63619 7875 63677 7876
rect 64003 7916 64061 7917
rect 64003 7876 64012 7916
rect 64052 7876 64061 7916
rect 64003 7875 64061 7876
rect 64963 7916 65021 7917
rect 64963 7876 64972 7916
rect 65012 7876 65021 7916
rect 64963 7875 65021 7876
rect 65251 7916 65309 7917
rect 65251 7876 65260 7916
rect 65300 7876 65309 7916
rect 65251 7875 65309 7876
rect 66211 7916 66269 7917
rect 66211 7876 66220 7916
rect 66260 7876 66269 7916
rect 66211 7875 66269 7876
rect 67171 7916 67229 7917
rect 67171 7876 67180 7916
rect 67220 7876 67229 7916
rect 67171 7875 67229 7876
rect 67363 7916 67421 7917
rect 67363 7876 67372 7916
rect 67412 7876 67421 7916
rect 67363 7875 67421 7876
rect 67651 7916 67709 7917
rect 67651 7876 67660 7916
rect 67700 7876 67709 7916
rect 67651 7875 67709 7876
rect 67843 7916 67901 7917
rect 67843 7876 67852 7916
rect 67892 7876 67901 7916
rect 67843 7875 67901 7876
rect 68707 7916 68765 7917
rect 68707 7876 68716 7916
rect 68756 7876 68765 7916
rect 68707 7875 68765 7876
rect 68899 7916 68957 7917
rect 68899 7876 68908 7916
rect 68948 7876 68957 7916
rect 68899 7875 68957 7876
rect 69771 7916 69813 7925
rect 69771 7876 69772 7916
rect 69812 7876 69813 7916
rect 69771 7867 69813 7876
rect 69955 7916 70013 7917
rect 69955 7876 69964 7916
rect 70004 7876 70013 7916
rect 69955 7875 70013 7876
rect 70147 7916 70205 7917
rect 70147 7876 70156 7916
rect 70196 7876 70205 7916
rect 70147 7875 70205 7876
rect 70347 7916 70389 7925
rect 70347 7876 70348 7916
rect 70388 7876 70389 7916
rect 70347 7867 70389 7876
rect 70531 7916 70589 7917
rect 70531 7876 70540 7916
rect 70580 7876 70589 7916
rect 70531 7875 70589 7876
rect 70731 7916 70773 7925
rect 70731 7876 70732 7916
rect 70772 7876 70773 7916
rect 70731 7867 70773 7876
rect 70915 7916 70973 7917
rect 70915 7876 70924 7916
rect 70964 7876 70973 7916
rect 70915 7875 70973 7876
rect 71115 7916 71157 7925
rect 71115 7876 71116 7916
rect 71156 7876 71157 7916
rect 71115 7867 71157 7876
rect 71683 7916 71741 7917
rect 71683 7876 71692 7916
rect 71732 7876 71741 7916
rect 71683 7875 71741 7876
rect 71875 7916 71933 7917
rect 71875 7876 71884 7916
rect 71924 7876 71933 7916
rect 71875 7875 71933 7876
rect 72067 7916 72125 7917
rect 72067 7876 72076 7916
rect 72116 7876 72125 7916
rect 72067 7875 72125 7876
rect 72259 7916 72317 7917
rect 72259 7876 72268 7916
rect 72308 7876 72317 7916
rect 72259 7875 72317 7876
rect 72739 7916 72797 7917
rect 72739 7876 72748 7916
rect 72788 7876 72797 7916
rect 72739 7875 72797 7876
rect 73987 7916 74045 7917
rect 73987 7876 73996 7916
rect 74036 7876 74045 7916
rect 73987 7875 74045 7876
rect 74187 7916 74229 7925
rect 74187 7876 74188 7916
rect 74228 7876 74229 7916
rect 74187 7867 74229 7876
rect 74371 7916 74429 7917
rect 74371 7876 74380 7916
rect 74420 7876 74429 7916
rect 74371 7875 74429 7876
rect 74571 7916 74613 7925
rect 74571 7876 74572 7916
rect 74612 7876 74613 7916
rect 74571 7867 74613 7876
rect 74851 7916 74909 7917
rect 74851 7876 74860 7916
rect 74900 7876 74909 7916
rect 74851 7875 74909 7876
rect 75235 7916 75293 7917
rect 75235 7876 75244 7916
rect 75284 7876 75293 7916
rect 75235 7875 75293 7876
rect 75427 7916 75485 7917
rect 75427 7876 75436 7916
rect 75476 7876 75485 7916
rect 75427 7875 75485 7876
rect 75723 7916 75765 7925
rect 75723 7876 75724 7916
rect 75764 7876 75765 7916
rect 75723 7867 75765 7876
rect 75907 7916 75965 7917
rect 75907 7876 75916 7916
rect 75956 7876 75965 7916
rect 75907 7875 75965 7876
rect 77539 7916 77597 7917
rect 77539 7876 77548 7916
rect 77588 7876 77597 7916
rect 77539 7875 77597 7876
rect 77739 7916 77781 7925
rect 77739 7876 77740 7916
rect 77780 7876 77781 7916
rect 77739 7867 77781 7876
rect 77923 7916 77981 7917
rect 77923 7876 77932 7916
rect 77972 7876 77981 7916
rect 77923 7875 77981 7876
rect 78123 7916 78165 7925
rect 78123 7876 78124 7916
rect 78164 7876 78165 7916
rect 78123 7867 78165 7876
rect 78403 7916 78461 7917
rect 78403 7876 78412 7916
rect 78452 7876 78461 7916
rect 78403 7875 78461 7876
rect 78595 7916 78653 7917
rect 78595 7876 78604 7916
rect 78644 7876 78653 7916
rect 78595 7875 78653 7876
rect 78795 7916 78837 7925
rect 78795 7876 78796 7916
rect 78836 7876 78837 7916
rect 78795 7867 78837 7876
rect 78979 7916 79037 7917
rect 78979 7876 78988 7916
rect 79028 7876 79037 7916
rect 78979 7875 79037 7876
rect 80715 7916 80757 7925
rect 80715 7876 80716 7916
rect 80756 7876 80757 7916
rect 80715 7867 80757 7876
rect 80899 7916 80957 7917
rect 80899 7876 80908 7916
rect 80948 7876 80957 7916
rect 80899 7875 80957 7876
rect 81099 7916 81141 7925
rect 81099 7876 81100 7916
rect 81140 7876 81141 7916
rect 81099 7867 81141 7876
rect 81283 7916 81341 7917
rect 81283 7876 81292 7916
rect 81332 7876 81341 7916
rect 81283 7875 81341 7876
rect 81483 7916 81525 7925
rect 81483 7876 81484 7916
rect 81524 7876 81525 7916
rect 81483 7867 81525 7876
rect 81667 7916 81725 7917
rect 81667 7876 81676 7916
rect 81716 7876 81725 7916
rect 81667 7875 81725 7876
rect 81867 7916 81909 7925
rect 81867 7876 81868 7916
rect 81908 7876 81909 7916
rect 81867 7867 81909 7876
rect 82051 7916 82109 7917
rect 82051 7876 82060 7916
rect 82100 7876 82109 7916
rect 82435 7899 82444 7939
rect 82484 7899 82493 7939
rect 89254 7939 89312 7940
rect 82435 7898 82493 7899
rect 82635 7916 82677 7925
rect 82051 7875 82109 7876
rect 82635 7876 82636 7916
rect 82676 7876 82677 7916
rect 82635 7867 82677 7876
rect 82819 7916 82877 7917
rect 82819 7876 82828 7916
rect 82868 7876 82877 7916
rect 82819 7875 82877 7876
rect 83019 7916 83061 7925
rect 83019 7876 83020 7916
rect 83060 7876 83061 7916
rect 83019 7867 83061 7876
rect 83211 7916 83253 7925
rect 83211 7876 83212 7916
rect 83252 7876 83253 7916
rect 83211 7867 83253 7876
rect 83395 7916 83453 7917
rect 83395 7876 83404 7916
rect 83444 7876 83453 7916
rect 83395 7875 83453 7876
rect 83587 7916 83645 7917
rect 83587 7876 83596 7916
rect 83636 7876 83645 7916
rect 83587 7875 83645 7876
rect 83787 7916 83829 7925
rect 83787 7876 83788 7916
rect 83828 7876 83829 7916
rect 83787 7867 83829 7876
rect 83971 7916 84029 7917
rect 83971 7876 83980 7916
rect 84020 7876 84029 7916
rect 83971 7875 84029 7876
rect 84171 7916 84213 7925
rect 84171 7876 84172 7916
rect 84212 7876 84213 7916
rect 84171 7867 84213 7876
rect 84355 7916 84413 7917
rect 84355 7876 84364 7916
rect 84404 7876 84413 7916
rect 84355 7875 84413 7876
rect 84555 7916 84597 7925
rect 84555 7876 84556 7916
rect 84596 7876 84597 7916
rect 84555 7867 84597 7876
rect 84739 7916 84797 7917
rect 84739 7876 84748 7916
rect 84788 7876 84797 7916
rect 84739 7875 84797 7876
rect 84939 7916 84981 7925
rect 84939 7876 84940 7916
rect 84980 7876 84981 7916
rect 84939 7867 84981 7876
rect 85123 7916 85181 7917
rect 85123 7876 85132 7916
rect 85172 7876 85181 7916
rect 85123 7875 85181 7876
rect 85323 7916 85365 7925
rect 85323 7876 85324 7916
rect 85364 7876 85365 7916
rect 85323 7867 85365 7876
rect 86763 7916 86805 7925
rect 86763 7876 86764 7916
rect 86804 7876 86805 7916
rect 86763 7867 86805 7876
rect 87811 7916 87869 7917
rect 87811 7876 87820 7916
rect 87860 7876 87869 7916
rect 87811 7875 87869 7876
rect 88011 7916 88053 7925
rect 88011 7876 88012 7916
rect 88052 7876 88053 7916
rect 88011 7867 88053 7876
rect 88203 7916 88245 7925
rect 88203 7876 88204 7916
rect 88244 7876 88245 7916
rect 88203 7867 88245 7876
rect 88387 7916 88445 7917
rect 88387 7876 88396 7916
rect 88436 7876 88445 7916
rect 88387 7875 88445 7876
rect 88579 7916 88637 7917
rect 88579 7876 88588 7916
rect 88628 7876 88637 7916
rect 88579 7875 88637 7876
rect 88683 7916 88725 7925
rect 88683 7876 88684 7916
rect 88724 7876 88725 7916
rect 89067 7916 89109 7925
rect 88683 7867 88725 7876
rect 88788 7903 88830 7912
rect 88788 7863 88789 7903
rect 88829 7863 88830 7903
rect 89067 7876 89068 7916
rect 89108 7876 89109 7916
rect 89254 7899 89263 7939
rect 89303 7899 89312 7939
rect 89635 7916 89693 7917
rect 89254 7898 89312 7899
rect 89451 7903 89493 7912
rect 89067 7867 89109 7876
rect 88788 7854 88830 7863
rect 89451 7863 89452 7903
rect 89492 7863 89493 7903
rect 89635 7876 89644 7916
rect 89684 7876 89693 7916
rect 89635 7875 89693 7876
rect 89451 7854 89493 7863
rect 36835 7833 36893 7834
rect 34539 7792 34540 7832
rect 34580 7792 34581 7832
rect 34539 7783 34581 7792
rect 49419 7832 49461 7841
rect 49419 7792 49420 7832
rect 49460 7792 49461 7832
rect 49419 7783 49461 7792
rect 49995 7832 50037 7841
rect 49995 7792 49996 7832
rect 50036 7792 50037 7832
rect 49995 7783 50037 7792
rect 69867 7832 69909 7841
rect 69867 7792 69868 7832
rect 69908 7792 69909 7832
rect 69867 7783 69909 7792
rect 70251 7832 70293 7841
rect 70251 7792 70252 7832
rect 70292 7792 70293 7832
rect 70251 7783 70293 7792
rect 70635 7832 70677 7841
rect 70635 7792 70636 7832
rect 70676 7792 70677 7832
rect 70635 7783 70677 7792
rect 71019 7832 71061 7841
rect 71019 7792 71020 7832
rect 71060 7792 71061 7832
rect 71019 7783 71061 7792
rect 74091 7832 74133 7841
rect 74091 7792 74092 7832
rect 74132 7792 74133 7832
rect 74091 7783 74133 7792
rect 74475 7832 74517 7841
rect 74475 7792 74476 7832
rect 74516 7792 74517 7832
rect 74475 7783 74517 7792
rect 75819 7832 75861 7841
rect 75819 7792 75820 7832
rect 75860 7792 75861 7832
rect 75819 7783 75861 7792
rect 77643 7832 77685 7841
rect 77643 7792 77644 7832
rect 77684 7792 77685 7832
rect 77643 7783 77685 7792
rect 78027 7832 78069 7841
rect 78027 7792 78028 7832
rect 78068 7792 78069 7832
rect 78027 7783 78069 7792
rect 78891 7832 78933 7841
rect 78891 7792 78892 7832
rect 78932 7792 78933 7832
rect 78891 7783 78933 7792
rect 80811 7832 80853 7841
rect 80811 7792 80812 7832
rect 80852 7792 80853 7832
rect 80811 7783 80853 7792
rect 81195 7832 81237 7841
rect 81195 7792 81196 7832
rect 81236 7792 81237 7832
rect 81195 7783 81237 7792
rect 81963 7832 82005 7841
rect 81963 7792 81964 7832
rect 82004 7792 82005 7832
rect 81963 7783 82005 7792
rect 82539 7832 82581 7841
rect 82539 7792 82540 7832
rect 82580 7792 82581 7832
rect 82539 7783 82581 7792
rect 82923 7832 82965 7841
rect 82923 7792 82924 7832
rect 82964 7792 82965 7832
rect 82923 7783 82965 7792
rect 83307 7832 83349 7841
rect 83307 7792 83308 7832
rect 83348 7792 83349 7832
rect 83307 7783 83349 7792
rect 84075 7832 84117 7841
rect 84075 7792 84076 7832
rect 84116 7792 84117 7832
rect 84075 7783 84117 7792
rect 84459 7832 84501 7841
rect 84459 7792 84460 7832
rect 84500 7792 84501 7832
rect 84459 7783 84501 7792
rect 87915 7832 87957 7841
rect 87915 7792 87916 7832
rect 87956 7792 87957 7832
rect 87915 7783 87957 7792
rect 88299 7832 88341 7841
rect 88299 7792 88300 7832
rect 88340 7792 88341 7832
rect 88299 7783 88341 7792
rect 89163 7832 89205 7841
rect 89163 7792 89164 7832
rect 89204 7792 89205 7832
rect 89163 7783 89205 7792
rect 89547 7832 89589 7841
rect 89547 7792 89548 7832
rect 89588 7792 89589 7832
rect 89547 7783 89589 7792
rect 22627 7748 22685 7749
rect 22627 7708 22636 7748
rect 22676 7708 22685 7748
rect 22627 7707 22685 7708
rect 23299 7748 23357 7749
rect 23299 7708 23308 7748
rect 23348 7708 23357 7748
rect 36739 7748 36797 7749
rect 23299 7707 23357 7708
rect 29739 7706 29781 7715
rect 36739 7708 36748 7748
rect 36788 7708 36797 7748
rect 36739 7707 36797 7708
rect 37411 7748 37469 7749
rect 37411 7708 37420 7748
rect 37460 7708 37469 7748
rect 37411 7707 37469 7708
rect 39723 7748 39765 7757
rect 39723 7708 39724 7748
rect 39764 7708 39765 7748
rect 45859 7748 45917 7749
rect 29739 7666 29740 7706
rect 29780 7666 29781 7706
rect 39723 7699 39765 7708
rect 44523 7706 44565 7715
rect 29739 7657 29781 7666
rect 44523 7666 44524 7706
rect 44564 7666 44565 7706
rect 44523 7657 44565 7666
rect 44715 7706 44757 7715
rect 45859 7708 45868 7748
rect 45908 7708 45917 7748
rect 45859 7707 45917 7708
rect 46531 7748 46589 7749
rect 46531 7708 46540 7748
rect 46580 7708 46589 7748
rect 46531 7707 46589 7708
rect 47203 7748 47261 7749
rect 47203 7708 47212 7748
rect 47252 7708 47261 7748
rect 47203 7707 47261 7708
rect 48451 7748 48509 7749
rect 48451 7708 48460 7748
rect 48500 7708 48509 7748
rect 48451 7707 48509 7708
rect 49603 7748 49661 7749
rect 49603 7708 49612 7748
rect 49652 7708 49661 7748
rect 54603 7748 54645 7757
rect 49603 7707 49661 7708
rect 44715 7666 44716 7706
rect 44756 7666 44757 7706
rect 44715 7657 44757 7666
rect 49803 7706 49845 7715
rect 49803 7666 49804 7706
rect 49844 7666 49845 7706
rect 54603 7708 54604 7748
rect 54644 7708 54645 7748
rect 54603 7699 54645 7708
rect 54891 7748 54933 7757
rect 54891 7708 54892 7748
rect 54932 7708 54933 7748
rect 54891 7699 54933 7708
rect 56523 7748 56565 7757
rect 56523 7708 56524 7748
rect 56564 7708 56565 7748
rect 56523 7699 56565 7708
rect 56907 7748 56949 7757
rect 56907 7708 56908 7748
rect 56948 7708 56949 7748
rect 56907 7699 56949 7708
rect 57771 7748 57813 7757
rect 57771 7708 57772 7748
rect 57812 7708 57813 7748
rect 57771 7699 57813 7708
rect 72835 7748 72893 7749
rect 72835 7708 72844 7748
rect 72884 7708 72893 7748
rect 72835 7707 72893 7708
rect 74755 7748 74813 7749
rect 74755 7708 74764 7748
rect 74804 7708 74813 7748
rect 74755 7707 74813 7708
rect 49803 7657 49845 7666
rect 1152 7580 98784 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 65408 7580
rect 65448 7540 65490 7580
rect 65530 7540 65572 7580
rect 65612 7540 65654 7580
rect 65694 7540 65736 7580
rect 65776 7540 80528 7580
rect 80568 7540 80610 7580
rect 80650 7540 80692 7580
rect 80732 7540 80774 7580
rect 80814 7540 80856 7580
rect 80896 7540 95648 7580
rect 95688 7540 95730 7580
rect 95770 7540 95812 7580
rect 95852 7540 95894 7580
rect 95934 7540 95976 7580
rect 96016 7540 98784 7580
rect 1152 7516 98784 7540
rect 77067 7454 77109 7463
rect 23011 7412 23069 7413
rect 23011 7372 23020 7412
rect 23060 7372 23069 7412
rect 23011 7371 23069 7372
rect 36651 7412 36693 7421
rect 36651 7372 36652 7412
rect 36692 7372 36693 7412
rect 36651 7363 36693 7372
rect 42987 7412 43029 7421
rect 42987 7372 42988 7412
rect 43028 7372 43029 7412
rect 42987 7363 43029 7372
rect 44611 7412 44669 7413
rect 44611 7372 44620 7412
rect 44660 7372 44669 7412
rect 44611 7371 44669 7372
rect 46627 7412 46685 7413
rect 46627 7372 46636 7412
rect 46676 7372 46685 7412
rect 46627 7371 46685 7372
rect 51339 7412 51381 7421
rect 51339 7372 51340 7412
rect 51380 7372 51381 7412
rect 51339 7363 51381 7372
rect 59787 7412 59829 7421
rect 59787 7372 59788 7412
rect 59828 7372 59829 7412
rect 59787 7363 59829 7372
rect 60547 7412 60605 7413
rect 60547 7372 60556 7412
rect 60596 7372 60605 7412
rect 60547 7371 60605 7372
rect 60843 7412 60885 7421
rect 77067 7414 77068 7454
rect 77108 7414 77109 7454
rect 60843 7372 60844 7412
rect 60884 7372 60885 7412
rect 60843 7363 60885 7372
rect 61795 7412 61853 7413
rect 61795 7372 61804 7412
rect 61844 7372 61853 7412
rect 61795 7371 61853 7372
rect 62083 7412 62141 7413
rect 62083 7372 62092 7412
rect 62132 7372 62141 7412
rect 77067 7405 77109 7414
rect 78403 7412 78461 7413
rect 62083 7371 62141 7372
rect 78403 7372 78412 7412
rect 78452 7372 78461 7412
rect 78403 7371 78461 7372
rect 78883 7412 78941 7413
rect 78883 7372 78892 7412
rect 78932 7372 78941 7412
rect 78883 7371 78941 7372
rect 79171 7412 79229 7413
rect 79171 7372 79180 7412
rect 79220 7372 79229 7412
rect 79171 7371 79229 7372
rect 86859 7412 86901 7421
rect 86859 7372 86860 7412
rect 86900 7372 86901 7412
rect 86859 7363 86901 7372
rect 89067 7412 89109 7421
rect 89067 7372 89068 7412
rect 89108 7372 89109 7412
rect 89067 7363 89109 7372
rect 60451 7328 60509 7329
rect 60451 7288 60460 7328
rect 60500 7288 60509 7328
rect 60451 7287 60509 7288
rect 78691 7328 78749 7329
rect 78691 7288 78700 7328
rect 78740 7288 78749 7328
rect 78691 7287 78749 7288
rect 85707 7328 85749 7337
rect 85707 7288 85708 7328
rect 85748 7288 85749 7328
rect 85707 7279 85749 7288
rect 10827 7257 10869 7266
rect 9667 7244 9725 7245
rect 9667 7204 9676 7244
rect 9716 7204 9725 7244
rect 9667 7203 9725 7204
rect 9867 7244 9909 7253
rect 9867 7204 9868 7244
rect 9908 7204 9909 7244
rect 9867 7195 9909 7204
rect 10051 7244 10109 7245
rect 10051 7204 10060 7244
rect 10100 7204 10109 7244
rect 10051 7203 10109 7204
rect 10251 7244 10293 7253
rect 10251 7204 10252 7244
rect 10292 7204 10293 7244
rect 10251 7195 10293 7204
rect 10627 7244 10685 7245
rect 10627 7204 10636 7244
rect 10676 7204 10685 7244
rect 10827 7217 10828 7257
rect 10868 7217 10869 7257
rect 70531 7265 70589 7266
rect 10827 7208 10869 7217
rect 11011 7244 11069 7245
rect 10627 7203 10685 7204
rect 11011 7204 11020 7244
rect 11060 7204 11069 7244
rect 11011 7203 11069 7204
rect 11211 7244 11253 7253
rect 11211 7204 11212 7244
rect 11252 7204 11253 7244
rect 11211 7195 11253 7204
rect 11875 7244 11933 7245
rect 11875 7204 11884 7244
rect 11924 7204 11933 7244
rect 11875 7203 11933 7204
rect 12075 7244 12117 7253
rect 12075 7204 12076 7244
rect 12116 7204 12117 7244
rect 12075 7195 12117 7204
rect 12547 7244 12605 7245
rect 12547 7204 12556 7244
rect 12596 7204 12605 7244
rect 12547 7203 12605 7204
rect 12747 7244 12789 7253
rect 12747 7204 12748 7244
rect 12788 7204 12789 7244
rect 12747 7195 12789 7204
rect 13411 7244 13469 7245
rect 13411 7204 13420 7244
rect 13460 7204 13469 7244
rect 13411 7203 13469 7204
rect 13603 7244 13661 7245
rect 13603 7204 13612 7244
rect 13652 7204 13661 7244
rect 13603 7203 13661 7204
rect 18699 7244 18741 7253
rect 18699 7204 18700 7244
rect 18740 7204 18741 7244
rect 18699 7195 18741 7204
rect 18883 7244 18941 7245
rect 18883 7204 18892 7244
rect 18932 7204 18941 7244
rect 18883 7203 18941 7204
rect 22731 7244 22773 7253
rect 22731 7204 22732 7244
rect 22772 7204 22773 7244
rect 22731 7195 22773 7204
rect 22923 7244 22965 7253
rect 22923 7204 22924 7244
rect 22964 7204 22965 7244
rect 22923 7195 22965 7204
rect 23019 7244 23061 7253
rect 23019 7204 23020 7244
rect 23060 7204 23061 7244
rect 23019 7195 23061 7204
rect 23979 7244 24021 7253
rect 23979 7204 23980 7244
rect 24020 7204 24021 7244
rect 23979 7195 24021 7204
rect 24171 7244 24213 7253
rect 24171 7204 24172 7244
rect 24212 7204 24213 7244
rect 24171 7195 24213 7204
rect 24363 7244 24405 7253
rect 24363 7204 24364 7244
rect 24404 7204 24405 7244
rect 24363 7195 24405 7204
rect 24555 7244 24597 7253
rect 24555 7204 24556 7244
rect 24596 7204 24597 7244
rect 24555 7195 24597 7204
rect 25035 7244 25077 7253
rect 25035 7204 25036 7244
rect 25076 7204 25077 7244
rect 25035 7195 25077 7204
rect 25131 7244 25173 7253
rect 25131 7204 25132 7244
rect 25172 7204 25173 7244
rect 25131 7195 25173 7204
rect 25219 7244 25277 7245
rect 25219 7204 25228 7244
rect 25268 7204 25277 7244
rect 25219 7203 25277 7204
rect 26955 7244 26997 7253
rect 26955 7204 26956 7244
rect 26996 7204 26997 7244
rect 26955 7195 26997 7204
rect 27147 7244 27189 7253
rect 27147 7204 27148 7244
rect 27188 7204 27189 7244
rect 27147 7195 27189 7204
rect 30019 7244 30077 7245
rect 30019 7204 30028 7244
rect 30068 7204 30077 7244
rect 30019 7203 30077 7204
rect 31179 7244 31221 7253
rect 31179 7204 31180 7244
rect 31220 7204 31221 7244
rect 31179 7195 31221 7204
rect 31651 7244 31709 7245
rect 32331 7244 32373 7253
rect 31651 7204 31660 7244
rect 31700 7204 31709 7244
rect 31651 7203 31709 7204
rect 31851 7243 31909 7244
rect 31851 7203 31860 7243
rect 31900 7203 31909 7243
rect 31851 7202 31909 7203
rect 32331 7204 32332 7244
rect 32372 7204 32373 7244
rect 32331 7195 32373 7204
rect 32619 7244 32661 7253
rect 32619 7204 32620 7244
rect 32660 7204 32661 7244
rect 32619 7195 32661 7204
rect 32803 7244 32861 7245
rect 32803 7204 32812 7244
rect 32852 7204 32861 7244
rect 32803 7203 32861 7204
rect 33867 7244 33909 7253
rect 33867 7204 33868 7244
rect 33908 7204 33909 7244
rect 33867 7195 33909 7204
rect 34059 7244 34101 7253
rect 34059 7204 34060 7244
rect 34100 7204 34101 7244
rect 34059 7195 34101 7204
rect 34251 7244 34293 7253
rect 34251 7204 34252 7244
rect 34292 7204 34293 7244
rect 34251 7195 34293 7204
rect 34443 7244 34485 7253
rect 34443 7204 34444 7244
rect 34484 7204 34485 7244
rect 34443 7195 34485 7204
rect 37323 7244 37365 7253
rect 37323 7204 37324 7244
rect 37364 7204 37365 7244
rect 37323 7195 37365 7204
rect 37515 7244 37557 7253
rect 37515 7204 37516 7244
rect 37556 7204 37557 7244
rect 37515 7195 37557 7204
rect 37707 7244 37749 7253
rect 37707 7204 37708 7244
rect 37748 7204 37749 7244
rect 37707 7195 37749 7204
rect 37899 7244 37941 7253
rect 37899 7204 37900 7244
rect 37940 7204 37941 7244
rect 37899 7195 37941 7204
rect 39139 7244 39197 7245
rect 39139 7204 39148 7244
rect 39188 7204 39197 7244
rect 39139 7203 39197 7204
rect 40099 7244 40157 7245
rect 40099 7204 40108 7244
rect 40148 7204 40157 7244
rect 40099 7203 40157 7204
rect 40387 7244 40445 7245
rect 40387 7204 40396 7244
rect 40436 7204 40445 7244
rect 40387 7203 40445 7204
rect 41347 7244 41405 7245
rect 41347 7204 41356 7244
rect 41396 7204 41405 7244
rect 41347 7203 41405 7204
rect 43459 7244 43517 7245
rect 43459 7204 43468 7244
rect 43508 7204 43517 7244
rect 43459 7203 43517 7204
rect 44331 7244 44373 7253
rect 44331 7204 44332 7244
rect 44372 7204 44373 7244
rect 44331 7195 44373 7204
rect 44523 7245 44565 7254
rect 44523 7205 44524 7245
rect 44564 7205 44565 7245
rect 44523 7196 44565 7205
rect 44619 7244 44661 7253
rect 44619 7204 44620 7244
rect 44660 7204 44661 7244
rect 44619 7195 44661 7204
rect 45763 7244 45821 7245
rect 45763 7204 45772 7244
rect 45812 7204 45821 7244
rect 45763 7203 45821 7204
rect 45955 7244 46013 7245
rect 45955 7204 45964 7244
rect 46004 7204 46013 7244
rect 45955 7203 46013 7204
rect 46539 7244 46581 7253
rect 46539 7204 46540 7244
rect 46580 7204 46581 7244
rect 46539 7195 46581 7204
rect 46635 7244 46677 7253
rect 46635 7204 46636 7244
rect 46676 7204 46677 7244
rect 46635 7195 46677 7204
rect 47107 7244 47165 7245
rect 47107 7204 47116 7244
rect 47156 7204 47165 7244
rect 47107 7203 47165 7204
rect 47299 7244 47357 7245
rect 47299 7204 47308 7244
rect 47348 7204 47357 7244
rect 47299 7203 47357 7204
rect 48547 7244 48605 7245
rect 48547 7204 48556 7244
rect 48596 7204 48605 7244
rect 48547 7203 48605 7204
rect 48739 7244 48797 7245
rect 48739 7204 48748 7244
rect 48788 7204 48797 7244
rect 48739 7203 48797 7204
rect 49027 7244 49085 7245
rect 49027 7204 49036 7244
rect 49076 7204 49085 7244
rect 49027 7203 49085 7204
rect 49227 7244 49269 7253
rect 49227 7204 49228 7244
rect 49268 7204 49269 7244
rect 49227 7195 49269 7204
rect 49315 7244 49373 7245
rect 49315 7204 49324 7244
rect 49364 7204 49373 7244
rect 49315 7203 49373 7204
rect 49515 7244 49557 7253
rect 49515 7204 49516 7244
rect 49556 7204 49557 7244
rect 49515 7195 49557 7204
rect 49707 7244 49749 7253
rect 49707 7204 49708 7244
rect 49748 7204 49749 7244
rect 49707 7195 49749 7204
rect 50083 7244 50141 7245
rect 50083 7204 50092 7244
rect 50132 7204 50141 7244
rect 50083 7203 50141 7204
rect 50371 7244 50429 7245
rect 50371 7204 50380 7244
rect 50420 7204 50429 7244
rect 50371 7203 50429 7204
rect 50563 7244 50621 7245
rect 50563 7204 50572 7244
rect 50612 7204 50621 7244
rect 50563 7203 50621 7204
rect 50755 7244 50813 7245
rect 50755 7204 50764 7244
rect 50804 7204 50813 7244
rect 50755 7203 50813 7204
rect 50947 7244 51005 7245
rect 50947 7204 50956 7244
rect 50996 7204 51005 7244
rect 50947 7203 51005 7204
rect 51243 7244 51285 7253
rect 51243 7204 51244 7244
rect 51284 7204 51285 7244
rect 51243 7195 51285 7204
rect 51531 7244 51573 7253
rect 51531 7204 51532 7244
rect 51572 7204 51573 7244
rect 51531 7195 51573 7204
rect 51715 7244 51773 7245
rect 51715 7204 51724 7244
rect 51764 7204 51773 7244
rect 51715 7203 51773 7204
rect 51819 7244 51861 7253
rect 51819 7204 51820 7244
rect 51860 7204 51861 7244
rect 51819 7195 51861 7204
rect 52003 7244 52061 7245
rect 52003 7204 52012 7244
rect 52052 7204 52061 7244
rect 52003 7203 52061 7204
rect 52291 7244 52349 7245
rect 52291 7204 52300 7244
rect 52340 7204 52349 7244
rect 52291 7203 52349 7204
rect 54307 7244 54365 7245
rect 54307 7204 54316 7244
rect 54356 7204 54365 7244
rect 54307 7203 54365 7204
rect 54507 7244 54549 7253
rect 54507 7204 54508 7244
rect 54548 7204 54549 7244
rect 54507 7195 54549 7204
rect 58347 7244 58389 7253
rect 58347 7204 58348 7244
rect 58388 7204 58389 7244
rect 58347 7195 58389 7204
rect 59203 7244 59261 7245
rect 59203 7204 59212 7244
rect 59252 7204 59261 7244
rect 59203 7203 59261 7204
rect 59395 7244 59453 7245
rect 59395 7204 59404 7244
rect 59444 7204 59453 7244
rect 59395 7203 59453 7204
rect 59779 7244 59837 7245
rect 59779 7204 59788 7244
rect 59828 7204 59837 7244
rect 59779 7203 59837 7204
rect 59979 7244 60021 7253
rect 59979 7204 59980 7244
rect 60020 7204 60021 7244
rect 59979 7195 60021 7204
rect 60067 7244 60125 7245
rect 60067 7204 60076 7244
rect 60116 7204 60125 7244
rect 60067 7203 60125 7204
rect 60267 7244 60309 7253
rect 60267 7204 60268 7244
rect 60308 7204 60309 7244
rect 60267 7195 60309 7204
rect 60363 7244 60405 7253
rect 60363 7204 60364 7244
rect 60404 7204 60405 7244
rect 60363 7195 60405 7204
rect 61891 7244 61949 7245
rect 61891 7204 61900 7244
rect 61940 7204 61949 7244
rect 61891 7203 61949 7204
rect 63043 7244 63101 7245
rect 63043 7204 63052 7244
rect 63092 7204 63101 7244
rect 63043 7203 63101 7204
rect 64003 7244 64061 7245
rect 64003 7204 64012 7244
rect 64052 7204 64061 7244
rect 64003 7203 64061 7204
rect 64483 7244 64541 7245
rect 64483 7204 64492 7244
rect 64532 7204 64541 7244
rect 64483 7203 64541 7204
rect 64675 7244 64733 7245
rect 64675 7204 64684 7244
rect 64724 7204 64733 7244
rect 64675 7203 64733 7204
rect 64963 7244 65021 7245
rect 64963 7204 64972 7244
rect 65012 7204 65021 7244
rect 64963 7203 65021 7204
rect 65155 7244 65213 7245
rect 65155 7204 65164 7244
rect 65204 7204 65213 7244
rect 65155 7203 65213 7204
rect 66787 7244 66845 7245
rect 66787 7204 66796 7244
rect 66836 7204 66845 7244
rect 66787 7203 66845 7204
rect 66979 7244 67037 7245
rect 66979 7204 66988 7244
rect 67028 7204 67037 7244
rect 66979 7203 67037 7204
rect 68043 7244 68085 7253
rect 68043 7204 68044 7244
rect 68084 7204 68085 7244
rect 68043 7195 68085 7204
rect 68235 7244 68277 7253
rect 68235 7204 68236 7244
rect 68276 7204 68277 7244
rect 68235 7195 68277 7204
rect 68523 7244 68565 7253
rect 68523 7204 68524 7244
rect 68564 7204 68565 7244
rect 68523 7195 68565 7204
rect 68715 7244 68757 7253
rect 68715 7204 68716 7244
rect 68756 7204 68757 7244
rect 68715 7195 68757 7204
rect 69003 7244 69045 7253
rect 69003 7204 69004 7244
rect 69044 7204 69045 7244
rect 69003 7195 69045 7204
rect 69195 7244 69237 7253
rect 69195 7204 69196 7244
rect 69236 7204 69237 7244
rect 70531 7225 70540 7265
rect 70580 7225 70589 7265
rect 70531 7224 70589 7225
rect 70731 7244 70773 7253
rect 69195 7195 69237 7204
rect 70731 7204 70732 7244
rect 70772 7204 70773 7244
rect 70731 7195 70773 7204
rect 74283 7244 74325 7253
rect 74283 7204 74284 7244
rect 74324 7204 74325 7244
rect 74283 7195 74325 7204
rect 74475 7244 74517 7253
rect 74475 7204 74476 7244
rect 74516 7204 74517 7244
rect 74475 7195 74517 7204
rect 74851 7244 74909 7245
rect 74851 7204 74860 7244
rect 74900 7204 74909 7244
rect 74851 7203 74909 7204
rect 75051 7244 75093 7253
rect 75051 7204 75052 7244
rect 75092 7204 75093 7244
rect 75051 7195 75093 7204
rect 75235 7244 75293 7245
rect 75235 7204 75244 7244
rect 75284 7204 75293 7244
rect 75235 7203 75293 7204
rect 75435 7244 75477 7253
rect 75435 7204 75436 7244
rect 75476 7204 75477 7244
rect 75435 7195 75477 7204
rect 77259 7244 77301 7253
rect 77259 7204 77260 7244
rect 77300 7204 77301 7244
rect 77259 7195 77301 7204
rect 77355 7244 77397 7253
rect 77355 7204 77356 7244
rect 77396 7204 77397 7244
rect 77355 7195 77397 7204
rect 77547 7244 77589 7253
rect 77547 7204 77548 7244
rect 77588 7204 77589 7244
rect 78219 7244 78261 7253
rect 77547 7195 77589 7204
rect 78019 7221 78077 7222
rect 78019 7181 78028 7221
rect 78068 7181 78077 7221
rect 78219 7204 78220 7244
rect 78260 7204 78261 7244
rect 78219 7195 78261 7204
rect 78499 7244 78557 7245
rect 78499 7204 78508 7244
rect 78548 7204 78557 7244
rect 78499 7203 78557 7204
rect 78979 7244 79037 7245
rect 78979 7204 78988 7244
rect 79028 7204 79037 7244
rect 78979 7203 79037 7204
rect 80803 7244 80861 7245
rect 80803 7204 80812 7244
rect 80852 7204 80861 7244
rect 80803 7203 80861 7204
rect 80995 7244 81053 7245
rect 80995 7204 81004 7244
rect 81044 7204 81053 7244
rect 80995 7203 81053 7204
rect 82635 7244 82677 7253
rect 82635 7204 82636 7244
rect 82676 7204 82677 7244
rect 82635 7195 82677 7204
rect 82827 7244 82869 7253
rect 82827 7204 82828 7244
rect 82868 7204 82869 7244
rect 82827 7195 82869 7204
rect 83019 7244 83061 7253
rect 83019 7204 83020 7244
rect 83060 7204 83061 7244
rect 83019 7195 83061 7204
rect 83203 7244 83261 7245
rect 83203 7204 83212 7244
rect 83252 7204 83261 7244
rect 83203 7203 83261 7204
rect 83403 7244 83445 7253
rect 83403 7204 83404 7244
rect 83444 7204 83445 7244
rect 83403 7195 83445 7204
rect 83587 7244 83645 7245
rect 83587 7204 83596 7244
rect 83636 7204 83645 7244
rect 83587 7203 83645 7204
rect 83787 7244 83829 7253
rect 83787 7204 83788 7244
rect 83828 7204 83829 7244
rect 83787 7195 83829 7204
rect 83971 7244 84029 7245
rect 83971 7204 83980 7244
rect 84020 7204 84029 7244
rect 83971 7203 84029 7204
rect 84171 7244 84213 7253
rect 84171 7204 84172 7244
rect 84212 7204 84213 7244
rect 84171 7195 84213 7204
rect 84355 7244 84413 7245
rect 84355 7204 84364 7244
rect 84404 7204 84413 7244
rect 84355 7203 84413 7204
rect 85611 7244 85653 7253
rect 85611 7204 85612 7244
rect 85652 7204 85653 7244
rect 85611 7195 85653 7204
rect 85795 7244 85853 7245
rect 85795 7204 85804 7244
rect 85844 7204 85853 7244
rect 85795 7203 85853 7204
rect 86371 7244 86429 7245
rect 86371 7204 86380 7244
rect 86420 7204 86429 7244
rect 86371 7203 86429 7204
rect 87523 7244 87581 7245
rect 87523 7204 87532 7244
rect 87572 7204 87581 7244
rect 87523 7203 87581 7204
rect 87715 7244 87773 7245
rect 87715 7204 87724 7244
rect 87764 7204 87773 7244
rect 87715 7203 87773 7204
rect 88003 7244 88061 7245
rect 88003 7204 88012 7244
rect 88052 7204 88061 7244
rect 88003 7203 88061 7204
rect 88203 7244 88245 7253
rect 88203 7204 88204 7244
rect 88244 7204 88245 7244
rect 88203 7195 88245 7204
rect 89451 7244 89493 7253
rect 89451 7204 89452 7244
rect 89492 7204 89493 7244
rect 89451 7195 89493 7204
rect 78019 7180 78077 7181
rect 30411 7160 30453 7169
rect 30411 7120 30412 7160
rect 30452 7120 30453 7160
rect 30411 7111 30453 7120
rect 33963 7160 34005 7169
rect 33963 7120 33964 7160
rect 34004 7120 34005 7160
rect 33963 7111 34005 7120
rect 36451 7160 36509 7161
rect 36451 7120 36460 7160
rect 36500 7120 36509 7160
rect 36451 7119 36509 7120
rect 46347 7160 46389 7169
rect 46347 7120 46348 7160
rect 46388 7120 46389 7160
rect 46347 7111 46389 7120
rect 56227 7160 56285 7161
rect 56227 7120 56236 7160
rect 56276 7120 56285 7160
rect 56227 7119 56285 7120
rect 56611 7160 56669 7161
rect 56611 7120 56620 7160
rect 56660 7120 56669 7160
rect 56611 7119 56669 7120
rect 57187 7160 57245 7161
rect 57187 7120 57196 7160
rect 57236 7120 57245 7160
rect 57187 7119 57245 7120
rect 61027 7160 61085 7161
rect 61027 7120 61036 7160
rect 61076 7120 61085 7160
rect 61027 7119 61085 7120
rect 11979 7076 12021 7085
rect 11979 7036 11980 7076
rect 12020 7036 12021 7076
rect 11979 7027 12021 7036
rect 29739 7076 29781 7085
rect 29739 7036 29740 7076
rect 29780 7036 29781 7076
rect 29739 7027 29781 7036
rect 31851 7076 31893 7085
rect 31851 7036 31852 7076
rect 31892 7036 31893 7076
rect 31851 7027 31893 7036
rect 32331 7076 32373 7085
rect 32331 7036 32332 7076
rect 32372 7036 32373 7076
rect 32331 7027 32373 7036
rect 51811 7076 51869 7077
rect 51811 7036 51820 7076
rect 51860 7036 51869 7076
rect 51811 7035 51869 7036
rect 58347 7076 58389 7085
rect 58347 7036 58348 7076
rect 58388 7036 58389 7076
rect 58347 7027 58389 7036
rect 9771 6992 9813 7001
rect 9771 6952 9772 6992
rect 9812 6952 9813 6992
rect 9771 6943 9813 6952
rect 10155 6992 10197 7001
rect 10155 6952 10156 6992
rect 10196 6952 10197 6992
rect 10155 6943 10197 6952
rect 10731 6992 10773 7001
rect 10731 6952 10732 6992
rect 10772 6952 10773 6992
rect 10731 6943 10773 6952
rect 11115 6992 11157 7001
rect 11115 6952 11116 6992
rect 11156 6952 11157 6992
rect 11115 6943 11157 6952
rect 12651 6992 12693 7001
rect 12651 6952 12652 6992
rect 12692 6952 12693 6992
rect 12651 6943 12693 6952
rect 18795 6992 18837 7001
rect 18795 6952 18796 6992
rect 18836 6952 18837 6992
rect 18795 6943 18837 6952
rect 23979 6992 24021 7001
rect 23979 6952 23980 6992
rect 24020 6952 24021 6992
rect 23979 6943 24021 6952
rect 24363 6992 24405 7001
rect 24363 6952 24364 6992
rect 24404 6952 24405 6992
rect 24363 6943 24405 6952
rect 27147 6992 27189 7001
rect 27147 6952 27148 6992
rect 27188 6952 27189 6992
rect 27147 6943 27189 6952
rect 32139 6992 32181 7001
rect 32139 6952 32140 6992
rect 32180 6952 32181 6992
rect 32139 6943 32181 6952
rect 32715 6992 32757 7001
rect 32715 6952 32716 6992
rect 32756 6952 32757 6992
rect 32715 6943 32757 6952
rect 34443 6992 34485 7001
rect 34443 6952 34444 6992
rect 34484 6952 34485 6992
rect 34443 6943 34485 6952
rect 36651 6992 36693 7001
rect 36651 6952 36652 6992
rect 36692 6952 36693 6992
rect 36651 6943 36693 6952
rect 37515 6992 37557 7001
rect 37515 6952 37516 6992
rect 37556 6952 37557 6992
rect 37515 6943 37557 6952
rect 37899 6992 37941 7001
rect 37899 6952 37900 6992
rect 37940 6952 37941 6992
rect 37899 6943 37941 6952
rect 49035 6992 49077 7001
rect 49035 6952 49036 6992
rect 49076 6952 49077 6992
rect 49035 6943 49077 6952
rect 49515 6992 49557 7001
rect 49515 6952 49516 6992
rect 49556 6952 49557 6992
rect 49515 6943 49557 6952
rect 52587 6992 52629 7001
rect 52587 6952 52588 6992
rect 52628 6952 52629 6992
rect 52587 6943 52629 6952
rect 54411 6992 54453 7001
rect 54411 6952 54412 6992
rect 54452 6952 54453 6992
rect 54411 6943 54453 6952
rect 56043 6992 56085 7001
rect 56043 6952 56044 6992
rect 56084 6952 56085 6992
rect 56043 6943 56085 6952
rect 56427 6992 56469 7001
rect 56427 6952 56428 6992
rect 56468 6952 56469 6992
rect 56427 6943 56469 6952
rect 57003 6992 57045 7001
rect 57003 6952 57004 6992
rect 57044 6952 57045 6992
rect 57003 6943 57045 6952
rect 58539 6992 58581 7001
rect 58539 6952 58540 6992
rect 58580 6952 58581 6992
rect 58539 6943 58581 6952
rect 60555 6992 60597 7001
rect 60555 6952 60556 6992
rect 60596 6952 60597 6992
rect 60555 6943 60597 6952
rect 68235 6992 68277 7001
rect 68235 6952 68236 6992
rect 68276 6952 68277 6992
rect 68235 6943 68277 6952
rect 68523 6992 68565 7001
rect 68523 6952 68524 6992
rect 68564 6952 68565 6992
rect 68523 6943 68565 6952
rect 69003 6992 69045 7001
rect 69003 6952 69004 6992
rect 69044 6952 69045 6992
rect 69003 6943 69045 6952
rect 70635 6992 70677 7001
rect 70635 6952 70636 6992
rect 70676 6952 70677 6992
rect 70635 6943 70677 6952
rect 74475 6992 74517 7001
rect 74475 6952 74476 6992
rect 74516 6952 74517 6992
rect 74475 6943 74517 6952
rect 74955 6992 74997 7001
rect 74955 6952 74956 6992
rect 74996 6952 74997 6992
rect 74955 6943 74997 6952
rect 75339 6992 75381 7001
rect 75339 6952 75340 6992
rect 75380 6952 75381 6992
rect 75339 6943 75381 6952
rect 78123 6992 78165 7001
rect 78123 6952 78124 6992
rect 78164 6952 78165 6992
rect 78123 6943 78165 6952
rect 82827 6992 82869 7001
rect 82827 6952 82828 6992
rect 82868 6952 82869 6992
rect 82827 6943 82869 6952
rect 83115 6992 83157 7001
rect 83115 6952 83116 6992
rect 83156 6952 83157 6992
rect 83115 6943 83157 6952
rect 83499 6992 83541 7001
rect 83499 6952 83500 6992
rect 83540 6952 83541 6992
rect 83499 6943 83541 6952
rect 83883 6992 83925 7001
rect 83883 6952 83884 6992
rect 83924 6952 83925 6992
rect 83883 6943 83925 6952
rect 84267 6992 84309 7001
rect 84267 6952 84268 6992
rect 84308 6952 84309 6992
rect 84267 6943 84309 6952
rect 88107 6992 88149 7001
rect 88107 6952 88108 6992
rect 88148 6952 88149 6992
rect 88107 6943 88149 6952
rect 1152 6824 98784 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 64168 6824
rect 64208 6784 64250 6824
rect 64290 6784 64332 6824
rect 64372 6784 64414 6824
rect 64454 6784 64496 6824
rect 64536 6784 79288 6824
rect 79328 6784 79370 6824
rect 79410 6784 79452 6824
rect 79492 6784 79534 6824
rect 79574 6784 79616 6824
rect 79656 6784 94408 6824
rect 94448 6784 94490 6824
rect 94530 6784 94572 6824
rect 94612 6784 94654 6824
rect 94694 6784 94736 6824
rect 94776 6784 98784 6824
rect 1152 6760 98784 6784
rect 15819 6656 15861 6665
rect 15819 6616 15820 6656
rect 15860 6616 15861 6656
rect 15819 6607 15861 6616
rect 36651 6656 36693 6665
rect 36651 6616 36652 6656
rect 36692 6616 36693 6656
rect 36651 6607 36693 6616
rect 48651 6656 48693 6665
rect 48651 6616 48652 6656
rect 48692 6616 48693 6656
rect 48651 6607 48693 6616
rect 51435 6656 51477 6665
rect 51435 6616 51436 6656
rect 51476 6616 51477 6656
rect 51435 6607 51477 6616
rect 51915 6656 51957 6665
rect 51915 6616 51916 6656
rect 51956 6616 51957 6656
rect 51915 6607 51957 6616
rect 52107 6656 52149 6665
rect 52107 6616 52108 6656
rect 52148 6616 52149 6656
rect 52107 6607 52149 6616
rect 52587 6656 52629 6665
rect 52587 6616 52588 6656
rect 52628 6616 52629 6656
rect 52587 6607 52629 6616
rect 59307 6656 59349 6665
rect 59307 6616 59308 6656
rect 59348 6616 59349 6656
rect 59307 6607 59349 6616
rect 62467 6656 62525 6657
rect 62467 6616 62476 6656
rect 62516 6616 62525 6656
rect 62467 6615 62525 6616
rect 74187 6656 74229 6665
rect 74187 6616 74188 6656
rect 74228 6616 74229 6656
rect 74187 6607 74229 6616
rect 77451 6656 77493 6665
rect 77451 6616 77452 6656
rect 77492 6616 77493 6656
rect 77451 6607 77493 6616
rect 79467 6656 79509 6665
rect 79467 6616 79468 6656
rect 79508 6616 79509 6656
rect 79467 6607 79509 6616
rect 87723 6656 87765 6665
rect 87723 6616 87724 6656
rect 87764 6616 87765 6656
rect 87723 6607 87765 6616
rect 16395 6572 16437 6581
rect 16395 6532 16396 6572
rect 16436 6532 16437 6572
rect 16395 6523 16437 6532
rect 18507 6572 18549 6581
rect 18507 6532 18508 6572
rect 18548 6532 18549 6572
rect 18507 6523 18549 6532
rect 29923 6572 29981 6573
rect 29923 6532 29932 6572
rect 29972 6532 29981 6572
rect 29923 6531 29981 6532
rect 32811 6572 32853 6581
rect 32811 6532 32812 6572
rect 32852 6532 32853 6572
rect 32811 6523 32853 6532
rect 35499 6572 35541 6581
rect 35499 6532 35500 6572
rect 35540 6532 35541 6572
rect 35499 6523 35541 6532
rect 35971 6572 36029 6573
rect 35971 6532 35980 6572
rect 36020 6532 36029 6572
rect 35971 6531 36029 6532
rect 47883 6572 47925 6581
rect 47883 6532 47884 6572
rect 47924 6532 47925 6572
rect 47883 6523 47925 6532
rect 49035 6572 49077 6581
rect 49035 6532 49036 6572
rect 49076 6532 49077 6572
rect 49035 6523 49077 6532
rect 53259 6572 53301 6581
rect 53259 6532 53260 6572
rect 53300 6532 53301 6572
rect 53259 6523 53301 6532
rect 54411 6572 54453 6581
rect 54411 6532 54412 6572
rect 54452 6532 54453 6572
rect 54411 6523 54453 6532
rect 54987 6572 55029 6581
rect 54987 6532 54988 6572
rect 55028 6532 55029 6572
rect 54987 6523 55029 6532
rect 57003 6572 57045 6581
rect 57003 6532 57004 6572
rect 57044 6532 57045 6572
rect 57003 6523 57045 6532
rect 61227 6572 61269 6581
rect 61227 6532 61228 6572
rect 61268 6532 61269 6572
rect 61227 6523 61269 6532
rect 62275 6572 62333 6573
rect 62275 6532 62284 6572
rect 62324 6532 62333 6572
rect 62275 6531 62333 6532
rect 67275 6572 67317 6581
rect 67275 6532 67276 6572
rect 67316 6532 67317 6572
rect 67275 6523 67317 6532
rect 71979 6572 72021 6581
rect 71979 6532 71980 6572
rect 72020 6532 72021 6572
rect 71979 6523 72021 6532
rect 79275 6572 79317 6581
rect 79275 6532 79276 6572
rect 79316 6532 79317 6572
rect 79275 6523 79317 6532
rect 79851 6572 79893 6581
rect 79851 6532 79852 6572
rect 79892 6532 79893 6572
rect 79851 6523 79893 6532
rect 80235 6572 80277 6581
rect 80235 6532 80236 6572
rect 80276 6532 80277 6572
rect 80235 6523 80277 6532
rect 82347 6572 82389 6581
rect 82347 6532 82348 6572
rect 82388 6532 82389 6572
rect 82347 6523 82389 6532
rect 83307 6572 83349 6581
rect 83307 6532 83308 6572
rect 83348 6532 83349 6572
rect 83307 6523 83349 6532
rect 1411 6488 1469 6489
rect 1411 6448 1420 6488
rect 1460 6448 1469 6488
rect 1411 6447 1469 6448
rect 19459 6488 19517 6489
rect 19459 6448 19468 6488
rect 19508 6448 19517 6488
rect 19459 6447 19517 6448
rect 20707 6488 20765 6489
rect 20707 6448 20716 6488
rect 20756 6448 20765 6488
rect 20707 6447 20765 6448
rect 21091 6488 21149 6489
rect 21091 6448 21100 6488
rect 21140 6448 21149 6488
rect 35683 6488 35741 6489
rect 21091 6447 21149 6448
rect 24651 6446 24693 6455
rect 35683 6448 35692 6488
rect 35732 6448 35741 6488
rect 38763 6488 38805 6497
rect 35683 6447 35741 6448
rect 10435 6404 10493 6405
rect 10435 6364 10444 6404
rect 10484 6364 10493 6404
rect 10435 6363 10493 6364
rect 10635 6404 10677 6413
rect 10635 6364 10636 6404
rect 10676 6364 10677 6404
rect 10635 6355 10677 6364
rect 15627 6404 15669 6413
rect 15627 6364 15628 6404
rect 15668 6364 15669 6404
rect 15627 6355 15669 6364
rect 15819 6404 15861 6413
rect 15819 6364 15820 6404
rect 15860 6364 15861 6404
rect 15819 6355 15861 6364
rect 16011 6404 16053 6413
rect 16011 6364 16012 6404
rect 16052 6364 16053 6404
rect 16011 6355 16053 6364
rect 16208 6401 16250 6410
rect 16208 6361 16209 6401
rect 16249 6361 16250 6401
rect 16208 6352 16250 6361
rect 16395 6404 16437 6413
rect 16395 6364 16396 6404
rect 16436 6364 16437 6404
rect 16395 6355 16437 6364
rect 16587 6404 16629 6413
rect 16587 6364 16588 6404
rect 16628 6364 16629 6404
rect 16587 6355 16629 6364
rect 17739 6404 17781 6413
rect 17739 6364 17740 6404
rect 17780 6364 17781 6404
rect 17739 6355 17781 6364
rect 17931 6404 17973 6413
rect 17931 6364 17932 6404
rect 17972 6364 17973 6404
rect 17931 6355 17973 6364
rect 18123 6404 18165 6413
rect 18123 6364 18124 6404
rect 18164 6364 18165 6404
rect 18123 6355 18165 6364
rect 18315 6404 18357 6413
rect 18315 6364 18316 6404
rect 18356 6364 18357 6404
rect 18315 6355 18357 6364
rect 18507 6404 18549 6413
rect 18507 6364 18508 6404
rect 18548 6364 18549 6404
rect 18507 6355 18549 6364
rect 18699 6404 18741 6413
rect 18699 6364 18700 6404
rect 18740 6364 18741 6404
rect 18699 6355 18741 6364
rect 18891 6404 18933 6413
rect 18891 6364 18892 6404
rect 18932 6364 18933 6404
rect 18891 6355 18933 6364
rect 19083 6404 19125 6413
rect 19083 6364 19084 6404
rect 19124 6364 19125 6404
rect 19083 6355 19125 6364
rect 19659 6404 19701 6413
rect 19659 6364 19660 6404
rect 19700 6364 19701 6404
rect 19659 6355 19701 6364
rect 19851 6404 19893 6413
rect 19851 6364 19852 6404
rect 19892 6364 19893 6404
rect 19851 6355 19893 6364
rect 23211 6404 23253 6413
rect 23211 6364 23212 6404
rect 23252 6364 23253 6404
rect 23211 6355 23253 6364
rect 23403 6404 23445 6413
rect 23403 6364 23404 6404
rect 23444 6364 23445 6404
rect 23403 6355 23445 6364
rect 23595 6404 23637 6413
rect 23595 6364 23596 6404
rect 23636 6364 23637 6404
rect 23595 6355 23637 6364
rect 23787 6404 23829 6413
rect 24651 6406 24652 6446
rect 24692 6406 24693 6446
rect 37803 6446 37845 6455
rect 27915 6417 27957 6426
rect 23787 6364 23788 6404
rect 23828 6364 23829 6404
rect 23787 6355 23829 6364
rect 24067 6404 24125 6405
rect 24067 6364 24076 6404
rect 24116 6364 24125 6404
rect 24067 6363 24125 6364
rect 24259 6404 24317 6405
rect 24259 6364 24268 6404
rect 24308 6364 24317 6404
rect 24259 6363 24317 6364
rect 24451 6404 24509 6405
rect 24451 6364 24460 6404
rect 24500 6364 24509 6404
rect 24651 6397 24693 6406
rect 24941 6405 24999 6406
rect 24451 6363 24509 6364
rect 24739 6390 24797 6391
rect 24739 6350 24748 6390
rect 24788 6350 24797 6390
rect 24941 6365 24950 6405
rect 24990 6365 24999 6405
rect 24941 6364 24999 6365
rect 25131 6404 25173 6413
rect 25131 6364 25132 6404
rect 25172 6364 25173 6404
rect 25131 6355 25173 6364
rect 25323 6404 25365 6413
rect 25323 6364 25324 6404
rect 25364 6364 25365 6404
rect 25323 6355 25365 6364
rect 25515 6404 25557 6413
rect 25515 6364 25516 6404
rect 25556 6364 25557 6404
rect 25515 6355 25557 6364
rect 26187 6404 26229 6413
rect 26187 6364 26188 6404
rect 26228 6364 26229 6404
rect 26187 6355 26229 6364
rect 26379 6404 26421 6413
rect 26379 6364 26380 6404
rect 26420 6364 26421 6404
rect 26379 6355 26421 6364
rect 26571 6404 26613 6413
rect 26571 6364 26572 6404
rect 26612 6364 26613 6404
rect 26571 6355 26613 6364
rect 26763 6404 26805 6413
rect 26763 6364 26764 6404
rect 26804 6364 26805 6404
rect 26763 6355 26805 6364
rect 26955 6404 26997 6413
rect 26955 6364 26956 6404
rect 26996 6364 26997 6404
rect 26955 6355 26997 6364
rect 27147 6404 27189 6413
rect 27147 6364 27148 6404
rect 27188 6364 27189 6404
rect 27147 6355 27189 6364
rect 27339 6404 27381 6413
rect 27339 6364 27340 6404
rect 27380 6364 27381 6404
rect 27339 6355 27381 6364
rect 27531 6404 27573 6413
rect 27531 6364 27532 6404
rect 27572 6364 27573 6404
rect 27531 6355 27573 6364
rect 27723 6404 27765 6413
rect 27723 6364 27724 6404
rect 27764 6364 27765 6404
rect 27915 6377 27916 6417
rect 27956 6377 27957 6417
rect 32235 6417 32277 6426
rect 27915 6368 27957 6377
rect 28483 6404 28541 6405
rect 27723 6355 27765 6364
rect 28483 6364 28492 6404
rect 28532 6364 28541 6404
rect 28483 6363 28541 6364
rect 28675 6404 28733 6405
rect 28675 6364 28684 6404
rect 28724 6364 28733 6404
rect 28675 6363 28733 6364
rect 29731 6404 29789 6405
rect 29731 6364 29740 6404
rect 29780 6364 29789 6404
rect 29731 6363 29789 6364
rect 29931 6404 29973 6413
rect 29931 6364 29932 6404
rect 29972 6364 29973 6404
rect 29931 6355 29973 6364
rect 30019 6404 30077 6405
rect 30019 6364 30028 6404
rect 30068 6364 30077 6404
rect 30019 6363 30077 6364
rect 31467 6404 31509 6413
rect 31467 6364 31468 6404
rect 31508 6364 31509 6404
rect 31467 6355 31509 6364
rect 31659 6404 31701 6413
rect 31659 6364 31660 6404
rect 31700 6364 31701 6404
rect 31659 6355 31701 6364
rect 31851 6404 31893 6413
rect 31851 6364 31852 6404
rect 31892 6364 31893 6404
rect 31851 6355 31893 6364
rect 32043 6404 32085 6413
rect 32043 6364 32044 6404
rect 32084 6364 32085 6404
rect 32235 6377 32236 6417
rect 32276 6377 32277 6417
rect 32235 6368 32277 6377
rect 32427 6404 32469 6413
rect 32043 6355 32085 6364
rect 32427 6364 32428 6404
rect 32468 6364 32469 6404
rect 32427 6355 32469 6364
rect 32619 6404 32661 6413
rect 32619 6364 32620 6404
rect 32660 6364 32661 6404
rect 32619 6355 32661 6364
rect 32811 6404 32853 6413
rect 32811 6364 32812 6404
rect 32852 6364 32853 6404
rect 32811 6355 32853 6364
rect 33195 6404 33237 6413
rect 33195 6364 33196 6404
rect 33236 6364 33237 6404
rect 33195 6355 33237 6364
rect 33291 6404 33333 6413
rect 33291 6364 33292 6404
rect 33332 6364 33333 6404
rect 33291 6355 33333 6364
rect 33675 6404 33717 6413
rect 33675 6364 33676 6404
rect 33716 6364 33717 6404
rect 33675 6355 33717 6364
rect 33867 6404 33909 6413
rect 33867 6364 33868 6404
rect 33908 6364 33909 6404
rect 33867 6355 33909 6364
rect 34059 6404 34101 6413
rect 34059 6364 34060 6404
rect 34100 6364 34101 6404
rect 34059 6355 34101 6364
rect 34251 6404 34293 6413
rect 34251 6364 34252 6404
rect 34292 6364 34293 6404
rect 34251 6355 34293 6364
rect 34443 6404 34485 6413
rect 34443 6364 34444 6404
rect 34484 6364 34485 6404
rect 34827 6404 34869 6413
rect 34443 6355 34485 6364
rect 34635 6393 34677 6402
rect 24739 6349 24797 6350
rect 34635 6353 34636 6393
rect 34676 6353 34677 6393
rect 34827 6364 34828 6404
rect 34868 6364 34869 6404
rect 34827 6355 34869 6364
rect 35019 6404 35061 6413
rect 35019 6364 35020 6404
rect 35060 6364 35061 6404
rect 35019 6355 35061 6364
rect 35875 6404 35933 6405
rect 35875 6364 35884 6404
rect 35924 6364 35933 6404
rect 35875 6363 35933 6364
rect 35979 6404 36021 6413
rect 37803 6406 37804 6446
rect 37844 6406 37845 6446
rect 38763 6448 38764 6488
rect 38804 6448 38805 6488
rect 38763 6439 38805 6448
rect 46627 6488 46685 6489
rect 46627 6448 46636 6488
rect 46676 6448 46685 6488
rect 46627 6447 46685 6448
rect 47203 6488 47261 6489
rect 47203 6448 47212 6488
rect 47252 6448 47261 6488
rect 47203 6447 47261 6448
rect 47587 6488 47645 6489
rect 47587 6448 47596 6488
rect 47636 6448 47645 6488
rect 47587 6447 47645 6448
rect 53059 6488 53117 6489
rect 53059 6448 53068 6488
rect 53108 6448 53117 6488
rect 53059 6447 53117 6448
rect 57483 6488 57525 6497
rect 57483 6448 57484 6488
rect 57524 6448 57525 6488
rect 57483 6439 57525 6448
rect 57955 6488 58013 6489
rect 57955 6448 57964 6488
rect 58004 6448 58013 6488
rect 57955 6447 58013 6448
rect 58819 6488 58877 6489
rect 58819 6448 58828 6488
rect 58868 6448 58877 6488
rect 58819 6447 58877 6448
rect 75715 6488 75773 6489
rect 75715 6448 75724 6488
rect 75764 6448 75773 6488
rect 75715 6447 75773 6448
rect 78795 6488 78837 6497
rect 78795 6448 78796 6488
rect 78836 6448 78837 6488
rect 77443 6446 77501 6447
rect 35979 6364 35980 6404
rect 36020 6364 36021 6404
rect 35979 6355 36021 6364
rect 36163 6404 36221 6405
rect 36163 6364 36172 6404
rect 36212 6364 36221 6404
rect 36163 6363 36221 6364
rect 36355 6404 36413 6405
rect 36355 6364 36364 6404
rect 36404 6364 36413 6404
rect 36355 6363 36413 6364
rect 37315 6404 37373 6405
rect 37315 6364 37324 6404
rect 37364 6364 37373 6404
rect 37315 6363 37373 6364
rect 37603 6404 37661 6405
rect 37603 6364 37612 6404
rect 37652 6364 37661 6404
rect 37803 6397 37845 6406
rect 37891 6404 37949 6405
rect 37603 6363 37661 6364
rect 37891 6364 37900 6404
rect 37940 6364 37949 6404
rect 37891 6363 37949 6364
rect 38091 6404 38133 6413
rect 38091 6364 38092 6404
rect 38132 6364 38133 6404
rect 38091 6355 38133 6364
rect 38283 6404 38325 6413
rect 38283 6364 38284 6404
rect 38324 6364 38325 6404
rect 38283 6355 38325 6364
rect 38667 6404 38709 6413
rect 38667 6364 38668 6404
rect 38708 6364 38709 6404
rect 38667 6355 38709 6364
rect 38859 6404 38901 6413
rect 38859 6364 38860 6404
rect 38900 6364 38901 6404
rect 38859 6355 38901 6364
rect 39331 6404 39389 6405
rect 39331 6364 39340 6404
rect 39380 6364 39389 6404
rect 39331 6363 39389 6364
rect 40203 6404 40245 6413
rect 40203 6364 40204 6404
rect 40244 6364 40245 6404
rect 40203 6355 40245 6364
rect 41635 6404 41693 6405
rect 41635 6364 41644 6404
rect 41684 6364 41693 6404
rect 41635 6363 41693 6364
rect 41923 6404 41981 6405
rect 41923 6364 41932 6404
rect 41972 6364 41981 6404
rect 41923 6363 41981 6364
rect 42795 6404 42837 6413
rect 42795 6364 42796 6404
rect 42836 6364 42837 6404
rect 42795 6355 42837 6364
rect 43459 6404 43517 6405
rect 43459 6364 43468 6404
rect 43508 6364 43517 6404
rect 43459 6363 43517 6364
rect 44331 6404 44373 6413
rect 44331 6364 44332 6404
rect 44372 6364 44373 6404
rect 44331 6355 44373 6364
rect 44707 6404 44765 6405
rect 44707 6364 44716 6404
rect 44756 6364 44765 6404
rect 44707 6363 44765 6364
rect 45667 6404 45725 6405
rect 45667 6364 45676 6404
rect 45716 6364 45725 6404
rect 45667 6363 45725 6364
rect 46147 6404 46205 6405
rect 46147 6364 46156 6404
rect 46196 6364 46205 6404
rect 46147 6363 46205 6364
rect 46339 6404 46397 6405
rect 46339 6364 46348 6404
rect 46388 6364 46397 6404
rect 46339 6363 46397 6364
rect 47875 6404 47933 6405
rect 47875 6364 47884 6404
rect 47924 6364 47933 6404
rect 47875 6363 47933 6364
rect 48075 6404 48117 6413
rect 48075 6364 48076 6404
rect 48116 6364 48117 6404
rect 48075 6355 48117 6364
rect 48163 6404 48221 6405
rect 48163 6364 48172 6404
rect 48212 6364 48221 6404
rect 48163 6363 48221 6364
rect 49315 6404 49373 6405
rect 49315 6364 49324 6404
rect 49364 6364 49373 6404
rect 49315 6363 49373 6364
rect 50371 6404 50429 6405
rect 50371 6364 50380 6404
rect 50420 6364 50429 6404
rect 50371 6363 50429 6364
rect 50659 6404 50717 6405
rect 50659 6364 50668 6404
rect 50708 6364 50717 6404
rect 50659 6363 50717 6364
rect 50851 6404 50909 6405
rect 50851 6364 50860 6404
rect 50900 6364 50909 6404
rect 50851 6363 50909 6364
rect 51139 6404 51197 6405
rect 51139 6364 51148 6404
rect 51188 6364 51197 6404
rect 51139 6363 51197 6364
rect 51243 6404 51285 6413
rect 51243 6364 51244 6404
rect 51284 6364 51285 6404
rect 51243 6355 51285 6364
rect 51427 6404 51485 6405
rect 51427 6364 51436 6404
rect 51476 6364 51485 6404
rect 51427 6363 51485 6364
rect 51627 6404 51669 6413
rect 51627 6364 51628 6404
rect 51668 6364 51669 6404
rect 51627 6355 51669 6364
rect 51915 6404 51957 6413
rect 51915 6364 51916 6404
rect 51956 6364 51957 6404
rect 52299 6404 52341 6413
rect 51915 6355 51957 6364
rect 52099 6390 52157 6391
rect 34635 6344 34677 6353
rect 52099 6350 52108 6390
rect 52148 6350 52157 6390
rect 52299 6364 52300 6404
rect 52340 6364 52341 6404
rect 52299 6355 52341 6364
rect 52387 6404 52445 6405
rect 52387 6364 52396 6404
rect 52436 6364 52445 6404
rect 52387 6363 52445 6364
rect 52579 6404 52637 6405
rect 52579 6364 52588 6404
rect 52628 6364 52637 6404
rect 52579 6363 52637 6364
rect 52779 6404 52821 6413
rect 52779 6364 52780 6404
rect 52820 6364 52821 6404
rect 52779 6355 52821 6364
rect 52867 6404 52925 6405
rect 52867 6364 52876 6404
rect 52916 6364 52925 6404
rect 52867 6363 52925 6364
rect 53923 6404 53981 6405
rect 53923 6364 53932 6404
rect 53972 6364 53981 6404
rect 53923 6363 53981 6364
rect 54115 6404 54173 6405
rect 54115 6364 54124 6404
rect 54164 6364 54173 6404
rect 54115 6363 54173 6364
rect 54411 6404 54453 6413
rect 54411 6364 54412 6404
rect 54452 6364 54453 6404
rect 54411 6355 54453 6364
rect 54987 6404 55029 6413
rect 54987 6364 54988 6404
rect 55028 6364 55029 6404
rect 54987 6355 55029 6364
rect 55555 6404 55613 6405
rect 55555 6364 55564 6404
rect 55604 6364 55613 6404
rect 55555 6363 55613 6364
rect 55747 6404 55805 6405
rect 55747 6364 55756 6404
rect 55796 6364 55805 6404
rect 55747 6363 55805 6364
rect 56043 6404 56085 6413
rect 56043 6364 56044 6404
rect 56084 6364 56085 6404
rect 56043 6355 56085 6364
rect 56227 6404 56285 6405
rect 56227 6364 56236 6404
rect 56276 6364 56285 6404
rect 56227 6363 56285 6364
rect 56523 6404 56565 6413
rect 56523 6364 56524 6404
rect 56564 6364 56565 6404
rect 56523 6355 56565 6364
rect 56715 6404 56757 6413
rect 56715 6364 56716 6404
rect 56756 6364 56757 6404
rect 56715 6355 56757 6364
rect 57003 6404 57045 6413
rect 57003 6364 57004 6404
rect 57044 6364 57045 6404
rect 57003 6355 57045 6364
rect 57387 6404 57429 6413
rect 57387 6364 57388 6404
rect 57428 6364 57429 6404
rect 57387 6355 57429 6364
rect 57579 6404 57621 6413
rect 57579 6364 57580 6404
rect 57620 6364 57621 6404
rect 57579 6355 57621 6364
rect 58243 6404 58301 6405
rect 58243 6364 58252 6404
rect 58292 6364 58301 6404
rect 58243 6363 58301 6364
rect 58435 6404 58493 6405
rect 58435 6364 58444 6404
rect 58484 6364 58493 6404
rect 58435 6363 58493 6364
rect 59883 6404 59925 6413
rect 59883 6364 59884 6404
rect 59924 6364 59925 6404
rect 59883 6355 59925 6364
rect 60267 6404 60309 6413
rect 60267 6364 60268 6404
rect 60308 6364 60309 6404
rect 60267 6355 60309 6364
rect 61027 6404 61085 6405
rect 61027 6364 61036 6404
rect 61076 6364 61085 6404
rect 61027 6363 61085 6364
rect 61219 6404 61277 6405
rect 61219 6364 61228 6404
rect 61268 6364 61277 6404
rect 61219 6363 61277 6364
rect 61803 6404 61845 6413
rect 61803 6364 61804 6404
rect 61844 6364 61845 6404
rect 61803 6355 61845 6364
rect 61899 6404 61941 6413
rect 61899 6364 61900 6404
rect 61940 6364 61941 6404
rect 61899 6355 61941 6364
rect 61995 6404 62037 6413
rect 61995 6364 61996 6404
rect 62036 6364 62037 6404
rect 61995 6355 62037 6364
rect 62091 6404 62133 6413
rect 62091 6364 62092 6404
rect 62132 6364 62133 6404
rect 62091 6355 62133 6364
rect 62659 6404 62717 6405
rect 62659 6364 62668 6404
rect 62708 6364 62717 6404
rect 62659 6363 62717 6364
rect 62947 6404 63005 6405
rect 62947 6364 62956 6404
rect 62996 6364 63005 6404
rect 62947 6363 63005 6364
rect 63147 6404 63189 6413
rect 63147 6364 63148 6404
rect 63188 6364 63189 6404
rect 63147 6355 63189 6364
rect 64003 6404 64061 6405
rect 64003 6364 64012 6404
rect 64052 6364 64061 6404
rect 64003 6363 64061 6364
rect 64963 6404 65021 6405
rect 64963 6364 64972 6404
rect 65012 6364 65021 6404
rect 64963 6363 65021 6364
rect 65251 6404 65309 6405
rect 65251 6364 65260 6404
rect 65300 6364 65309 6404
rect 65251 6363 65309 6364
rect 66211 6404 66269 6405
rect 66211 6364 66220 6404
rect 66260 6364 66269 6404
rect 66211 6363 66269 6364
rect 66403 6404 66461 6405
rect 66403 6364 66412 6404
rect 66452 6364 66461 6404
rect 66403 6363 66461 6364
rect 66595 6404 66653 6405
rect 66595 6364 66604 6404
rect 66644 6364 66653 6404
rect 66595 6363 66653 6364
rect 67179 6404 67221 6413
rect 67179 6364 67180 6404
rect 67220 6364 67221 6404
rect 67179 6355 67221 6364
rect 67363 6404 67421 6405
rect 67363 6364 67372 6404
rect 67412 6364 67421 6404
rect 67363 6363 67421 6364
rect 67555 6404 67613 6405
rect 67555 6364 67564 6404
rect 67604 6364 67613 6404
rect 67555 6363 67613 6364
rect 67747 6404 67805 6405
rect 67747 6364 67756 6404
rect 67796 6364 67805 6404
rect 67747 6363 67805 6364
rect 68043 6404 68085 6413
rect 68043 6364 68044 6404
rect 68084 6364 68085 6404
rect 68043 6355 68085 6364
rect 68235 6404 68277 6413
rect 68235 6364 68236 6404
rect 68276 6364 68277 6404
rect 68235 6355 68277 6364
rect 68611 6404 68669 6405
rect 68611 6364 68620 6404
rect 68660 6364 68669 6404
rect 68611 6363 68669 6364
rect 68803 6404 68861 6405
rect 68803 6364 68812 6404
rect 68852 6364 68861 6404
rect 68803 6363 68861 6364
rect 69099 6404 69141 6413
rect 69099 6364 69100 6404
rect 69140 6364 69141 6404
rect 69099 6355 69141 6364
rect 69291 6404 69333 6413
rect 69291 6364 69292 6404
rect 69332 6364 69333 6404
rect 69291 6355 69333 6364
rect 69483 6404 69525 6413
rect 69483 6364 69484 6404
rect 69524 6364 69525 6404
rect 69483 6355 69525 6364
rect 69675 6404 69717 6413
rect 69675 6364 69676 6404
rect 69716 6364 69717 6404
rect 69675 6355 69717 6364
rect 71019 6404 71061 6413
rect 71019 6364 71020 6404
rect 71060 6364 71061 6404
rect 71019 6355 71061 6364
rect 71779 6404 71837 6405
rect 71779 6364 71788 6404
rect 71828 6364 71837 6404
rect 71779 6363 71837 6364
rect 71971 6404 72029 6405
rect 71971 6364 71980 6404
rect 72020 6364 72029 6404
rect 71971 6363 72029 6364
rect 72651 6404 72693 6413
rect 72651 6364 72652 6404
rect 72692 6364 72693 6404
rect 72651 6355 72693 6364
rect 72835 6404 72893 6405
rect 72835 6364 72844 6404
rect 72884 6364 72893 6404
rect 72835 6363 72893 6364
rect 73219 6404 73277 6405
rect 73219 6364 73228 6404
rect 73268 6364 73277 6404
rect 73219 6363 73277 6364
rect 73411 6404 73469 6405
rect 73411 6364 73420 6404
rect 73460 6364 73469 6404
rect 73411 6363 73469 6364
rect 73995 6404 74037 6413
rect 73995 6364 73996 6404
rect 74036 6364 74037 6404
rect 73995 6355 74037 6364
rect 74187 6404 74229 6413
rect 74187 6364 74188 6404
rect 74228 6364 74229 6404
rect 74571 6404 74613 6413
rect 74187 6355 74229 6364
rect 74372 6393 74414 6402
rect 52099 6349 52157 6350
rect 74372 6353 74373 6393
rect 74413 6353 74414 6393
rect 74571 6364 74572 6404
rect 74612 6364 74613 6404
rect 74571 6355 74613 6364
rect 74763 6404 74805 6413
rect 74763 6364 74764 6404
rect 74804 6364 74805 6404
rect 74763 6355 74805 6364
rect 74955 6404 74997 6413
rect 74955 6364 74956 6404
rect 74996 6364 74997 6404
rect 74955 6355 74997 6364
rect 75147 6404 75189 6413
rect 75147 6364 75148 6404
rect 75188 6364 75189 6404
rect 75147 6355 75189 6364
rect 75339 6404 75381 6413
rect 75339 6364 75340 6404
rect 75380 6364 75381 6404
rect 75339 6355 75381 6364
rect 76779 6404 76821 6413
rect 77443 6406 77452 6446
rect 77492 6406 77501 6446
rect 78795 6439 78837 6448
rect 79651 6488 79709 6489
rect 79651 6448 79660 6488
rect 79700 6448 79709 6488
rect 79651 6447 79709 6448
rect 80035 6488 80093 6489
rect 80035 6448 80044 6488
rect 80084 6448 80093 6488
rect 80035 6447 80093 6448
rect 80419 6488 80477 6489
rect 80419 6448 80428 6488
rect 80468 6448 80477 6488
rect 80419 6447 80477 6448
rect 81955 6488 82013 6489
rect 81955 6448 81964 6488
rect 82004 6448 82013 6488
rect 81955 6447 82013 6448
rect 83595 6488 83637 6497
rect 83595 6448 83596 6488
rect 83636 6448 83637 6488
rect 83595 6439 83637 6448
rect 98467 6488 98525 6489
rect 98467 6448 98476 6488
rect 98516 6448 98525 6488
rect 98467 6447 98525 6448
rect 77443 6405 77501 6406
rect 76779 6364 76780 6404
rect 76820 6364 76821 6404
rect 76779 6355 76821 6364
rect 77643 6404 77685 6413
rect 77643 6364 77644 6404
rect 77684 6364 77685 6404
rect 77643 6355 77685 6364
rect 77731 6404 77789 6405
rect 77731 6364 77740 6404
rect 77780 6364 77789 6404
rect 77731 6363 77789 6364
rect 78699 6404 78741 6413
rect 78699 6364 78700 6404
rect 78740 6364 78741 6404
rect 78699 6355 78741 6364
rect 78891 6404 78933 6413
rect 78891 6364 78892 6404
rect 78932 6364 78933 6404
rect 78891 6355 78933 6364
rect 79083 6404 79125 6413
rect 79083 6364 79084 6404
rect 79124 6364 79125 6404
rect 79083 6355 79125 6364
rect 79275 6404 79317 6413
rect 79275 6364 79276 6404
rect 79316 6364 79317 6404
rect 79275 6355 79317 6364
rect 82155 6404 82197 6413
rect 82155 6364 82156 6404
rect 82196 6364 82197 6404
rect 82155 6355 82197 6364
rect 82347 6404 82389 6413
rect 82347 6364 82348 6404
rect 82388 6364 82389 6404
rect 82347 6355 82389 6364
rect 82731 6404 82773 6413
rect 82731 6364 82732 6404
rect 82772 6364 82773 6404
rect 82731 6355 82773 6364
rect 82923 6404 82965 6413
rect 82923 6364 82924 6404
rect 82964 6364 82965 6404
rect 82923 6355 82965 6364
rect 83115 6404 83157 6413
rect 83115 6364 83116 6404
rect 83156 6364 83157 6404
rect 83115 6355 83157 6364
rect 83307 6404 83349 6413
rect 83307 6364 83308 6404
rect 83348 6364 83349 6404
rect 83307 6355 83349 6364
rect 83499 6404 83541 6413
rect 83499 6364 83500 6404
rect 83540 6364 83541 6404
rect 83499 6355 83541 6364
rect 83691 6404 83733 6413
rect 83691 6364 83692 6404
rect 83732 6364 83733 6404
rect 83691 6355 83733 6364
rect 83883 6404 83925 6413
rect 83883 6364 83884 6404
rect 83924 6364 83925 6404
rect 83883 6355 83925 6364
rect 84075 6404 84117 6413
rect 84075 6364 84076 6404
rect 84116 6364 84117 6404
rect 84075 6355 84117 6364
rect 84643 6404 84701 6405
rect 84643 6364 84652 6404
rect 84692 6364 84701 6404
rect 84643 6363 84701 6364
rect 86667 6404 86709 6413
rect 86667 6364 86668 6404
rect 86708 6364 86709 6404
rect 86667 6355 86709 6364
rect 86851 6404 86909 6405
rect 86851 6364 86860 6404
rect 86900 6364 86909 6404
rect 86851 6363 86909 6364
rect 87427 6404 87485 6405
rect 87427 6364 87436 6404
rect 87476 6364 87485 6404
rect 87427 6363 87485 6364
rect 74372 6344 74414 6353
rect 10539 6320 10581 6329
rect 10539 6280 10540 6320
rect 10580 6280 10581 6320
rect 10539 6271 10581 6280
rect 16107 6320 16149 6329
rect 16107 6280 16108 6320
rect 16148 6280 16149 6320
rect 16107 6271 16149 6280
rect 19755 6320 19797 6329
rect 19755 6280 19756 6320
rect 19796 6280 19797 6320
rect 19755 6271 19797 6280
rect 27051 6320 27093 6329
rect 27051 6280 27052 6320
rect 27092 6280 27093 6320
rect 27051 6271 27093 6280
rect 27435 6320 27477 6329
rect 27435 6280 27436 6320
rect 27476 6280 27477 6320
rect 27435 6271 27477 6280
rect 27819 6320 27861 6329
rect 27819 6280 27820 6320
rect 27860 6280 27861 6320
rect 27819 6271 27861 6280
rect 32331 6320 32373 6329
rect 32331 6280 32332 6320
rect 32372 6280 32373 6320
rect 32331 6271 32373 6280
rect 34155 6320 34197 6329
rect 34155 6280 34156 6320
rect 34196 6280 34197 6320
rect 34155 6271 34197 6280
rect 40771 6320 40829 6321
rect 40771 6280 40780 6320
rect 40820 6280 40829 6320
rect 40771 6279 40829 6280
rect 50179 6320 50237 6321
rect 50179 6280 50188 6320
rect 50228 6280 50237 6320
rect 50179 6279 50237 6280
rect 56139 6320 56181 6329
rect 56139 6280 56140 6320
rect 56180 6280 56181 6320
rect 56139 6271 56181 6280
rect 56619 6320 56661 6329
rect 56619 6280 56620 6320
rect 56660 6280 56661 6320
rect 56619 6271 56661 6280
rect 60555 6320 60597 6329
rect 60555 6280 60556 6320
rect 60596 6280 60597 6320
rect 60555 6271 60597 6280
rect 63051 6320 63093 6329
rect 63051 6280 63052 6320
rect 63092 6280 63093 6320
rect 63051 6271 63093 6280
rect 71307 6320 71349 6329
rect 71307 6280 71308 6320
rect 71348 6280 71349 6320
rect 71307 6271 71349 6280
rect 72747 6320 72789 6329
rect 72747 6280 72748 6320
rect 72788 6280 72789 6320
rect 72747 6271 72789 6280
rect 82827 6320 82869 6329
rect 82827 6280 82828 6320
rect 82868 6280 82869 6320
rect 82827 6271 82869 6280
rect 83979 6320 84021 6329
rect 83979 6280 83980 6320
rect 84020 6280 84021 6320
rect 83979 6271 84021 6280
rect 84835 6320 84893 6321
rect 84835 6280 84844 6320
rect 84884 6280 84893 6320
rect 84835 6279 84893 6280
rect 86763 6320 86805 6329
rect 86763 6280 86764 6320
rect 86804 6280 86805 6320
rect 86763 6271 86805 6280
rect 1227 6236 1269 6245
rect 1227 6196 1228 6236
rect 1268 6196 1269 6236
rect 1227 6187 1269 6196
rect 17835 6236 17877 6245
rect 17835 6196 17836 6236
rect 17876 6196 17877 6236
rect 17835 6187 17877 6196
rect 18219 6236 18261 6245
rect 18219 6196 18220 6236
rect 18260 6196 18261 6236
rect 18219 6187 18261 6196
rect 18987 6236 19029 6245
rect 18987 6196 18988 6236
rect 19028 6196 19029 6236
rect 18987 6187 19029 6196
rect 19275 6236 19317 6245
rect 19275 6196 19276 6236
rect 19316 6196 19317 6236
rect 19275 6187 19317 6196
rect 20523 6236 20565 6245
rect 20523 6196 20524 6236
rect 20564 6196 20565 6236
rect 20523 6187 20565 6196
rect 20907 6236 20949 6245
rect 20907 6196 20908 6236
rect 20948 6196 20949 6236
rect 20907 6187 20949 6196
rect 23307 6236 23349 6245
rect 23307 6196 23308 6236
rect 23348 6196 23349 6236
rect 23307 6187 23349 6196
rect 23691 6236 23733 6245
rect 23691 6196 23692 6236
rect 23732 6196 23733 6236
rect 23691 6187 23733 6196
rect 24459 6236 24501 6245
rect 24459 6196 24460 6236
rect 24500 6196 24501 6236
rect 24459 6187 24501 6196
rect 25035 6236 25077 6245
rect 25035 6196 25036 6236
rect 25076 6196 25077 6236
rect 25035 6187 25077 6196
rect 25419 6236 25461 6245
rect 25419 6196 25420 6236
rect 25460 6196 25461 6236
rect 25419 6187 25461 6196
rect 26283 6236 26325 6245
rect 26283 6196 26284 6236
rect 26324 6196 26325 6236
rect 26283 6187 26325 6196
rect 26667 6236 26709 6245
rect 26667 6196 26668 6236
rect 26708 6196 26709 6236
rect 26667 6187 26709 6196
rect 31563 6236 31605 6245
rect 31563 6196 31564 6236
rect 31604 6196 31605 6236
rect 31563 6187 31605 6196
rect 31947 6236 31989 6245
rect 31947 6196 31948 6236
rect 31988 6196 31989 6236
rect 31947 6187 31989 6196
rect 32995 6236 33053 6237
rect 32995 6196 33004 6236
rect 33044 6196 33053 6236
rect 32995 6195 33053 6196
rect 33771 6236 33813 6245
rect 33771 6196 33772 6236
rect 33812 6196 33813 6236
rect 33771 6187 33813 6196
rect 34539 6236 34581 6245
rect 34539 6196 34540 6236
rect 34580 6196 34581 6236
rect 34539 6187 34581 6196
rect 34923 6236 34965 6245
rect 34923 6196 34924 6236
rect 34964 6196 34965 6236
rect 34923 6187 34965 6196
rect 37611 6236 37653 6245
rect 37611 6196 37612 6236
rect 37652 6196 37653 6236
rect 37611 6187 37653 6196
rect 38187 6236 38229 6245
rect 38187 6196 38188 6236
rect 38228 6196 38229 6236
rect 38187 6187 38229 6196
rect 46827 6236 46869 6245
rect 46827 6196 46828 6236
rect 46868 6196 46869 6236
rect 46827 6187 46869 6196
rect 47019 6236 47061 6245
rect 47019 6196 47020 6236
rect 47060 6196 47061 6236
rect 47019 6187 47061 6196
rect 47403 6236 47445 6245
rect 47403 6196 47404 6236
rect 47444 6196 47445 6236
rect 47403 6187 47445 6196
rect 47883 6236 47925 6245
rect 47883 6196 47884 6236
rect 47924 6196 47925 6236
rect 47883 6187 47925 6196
rect 50467 6236 50525 6237
rect 50467 6196 50476 6236
rect 50516 6196 50525 6236
rect 50467 6195 50525 6196
rect 51435 6236 51477 6245
rect 51435 6196 51436 6236
rect 51476 6196 51477 6236
rect 51435 6187 51477 6196
rect 52587 6236 52629 6245
rect 52587 6196 52588 6236
rect 52628 6196 52629 6236
rect 52587 6187 52629 6196
rect 54603 6236 54645 6245
rect 54603 6196 54604 6236
rect 54644 6196 54645 6236
rect 54603 6187 54645 6196
rect 54795 6236 54837 6245
rect 54795 6196 54796 6236
rect 54836 6196 54837 6236
rect 54795 6187 54837 6196
rect 57195 6236 57237 6245
rect 57195 6196 57196 6236
rect 57236 6196 57237 6236
rect 57195 6187 57237 6196
rect 57771 6236 57813 6245
rect 57771 6196 57772 6236
rect 57812 6196 57813 6236
rect 57771 6187 57813 6196
rect 58635 6236 58677 6245
rect 58635 6196 58636 6236
rect 58676 6196 58677 6236
rect 58635 6187 58677 6196
rect 60739 6236 60797 6237
rect 60739 6196 60748 6236
rect 60788 6196 60797 6236
rect 60739 6195 60797 6196
rect 62755 6236 62813 6237
rect 62755 6196 62764 6236
rect 62804 6196 62813 6236
rect 62755 6195 62813 6196
rect 68139 6236 68181 6245
rect 68139 6196 68140 6236
rect 68180 6196 68181 6236
rect 68139 6187 68181 6196
rect 69195 6236 69237 6245
rect 69195 6196 69196 6236
rect 69236 6196 69237 6236
rect 69195 6187 69237 6196
rect 69579 6236 69621 6245
rect 69579 6196 69580 6236
rect 69620 6196 69621 6236
rect 69579 6187 69621 6196
rect 71491 6236 71549 6237
rect 71491 6196 71500 6236
rect 71540 6196 71549 6236
rect 71491 6195 71549 6196
rect 74475 6236 74517 6245
rect 74475 6196 74476 6236
rect 74516 6196 74517 6236
rect 74475 6187 74517 6196
rect 74859 6236 74901 6245
rect 74859 6196 74860 6236
rect 74900 6196 74901 6236
rect 74859 6187 74901 6196
rect 75243 6236 75285 6245
rect 75243 6196 75244 6236
rect 75284 6196 75285 6236
rect 75243 6187 75285 6196
rect 75531 6236 75573 6245
rect 75531 6196 75532 6236
rect 75572 6196 75573 6236
rect 75531 6187 75573 6196
rect 77059 6236 77117 6237
rect 77059 6196 77068 6236
rect 77108 6196 77117 6236
rect 77059 6195 77117 6196
rect 77251 6236 77309 6237
rect 77251 6196 77260 6236
rect 77300 6196 77309 6236
rect 77251 6195 77309 6196
rect 81771 6236 81813 6245
rect 81771 6196 81772 6236
rect 81812 6196 81813 6236
rect 81771 6187 81813 6196
rect 84547 6236 84605 6237
rect 84547 6196 84556 6236
rect 84596 6196 84605 6236
rect 84547 6195 84605 6196
rect 98667 6236 98709 6245
rect 98667 6196 98668 6236
rect 98708 6196 98709 6236
rect 98667 6187 98709 6196
rect 1152 6068 98784 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 65408 6068
rect 65448 6028 65490 6068
rect 65530 6028 65572 6068
rect 65612 6028 65654 6068
rect 65694 6028 65736 6068
rect 65776 6028 80528 6068
rect 80568 6028 80610 6068
rect 80650 6028 80692 6068
rect 80732 6028 80774 6068
rect 80814 6028 80856 6068
rect 80896 6028 95648 6068
rect 95688 6028 95730 6068
rect 95770 6028 95812 6068
rect 95852 6028 95894 6068
rect 95934 6028 95976 6068
rect 96016 6028 98784 6068
rect 1152 6004 98784 6028
rect 16971 5900 17013 5909
rect 16971 5860 16972 5900
rect 17012 5860 17013 5900
rect 16971 5851 17013 5860
rect 23019 5900 23061 5909
rect 23019 5860 23020 5900
rect 23060 5860 23061 5900
rect 23019 5851 23061 5860
rect 45387 5900 45429 5909
rect 45387 5860 45388 5900
rect 45428 5860 45429 5900
rect 45387 5851 45429 5860
rect 53355 5900 53397 5909
rect 53355 5860 53356 5900
rect 53396 5860 53397 5900
rect 53355 5851 53397 5860
rect 56811 5900 56853 5909
rect 56811 5860 56812 5900
rect 56852 5860 56853 5900
rect 56811 5851 56853 5860
rect 61315 5900 61373 5901
rect 61315 5860 61324 5900
rect 61364 5860 61373 5900
rect 61315 5859 61373 5860
rect 65067 5900 65109 5909
rect 65067 5860 65068 5900
rect 65108 5860 65109 5900
rect 65067 5851 65109 5860
rect 72075 5900 72117 5909
rect 72075 5860 72076 5900
rect 72116 5860 72117 5900
rect 72075 5851 72117 5860
rect 79371 5900 79413 5909
rect 79371 5860 79372 5900
rect 79412 5860 79413 5900
rect 79371 5851 79413 5860
rect 41731 5816 41789 5817
rect 41731 5776 41740 5816
rect 41780 5776 41789 5816
rect 41731 5775 41789 5776
rect 37035 5743 37077 5752
rect 15339 5732 15381 5741
rect 15339 5692 15340 5732
rect 15380 5692 15381 5732
rect 15339 5683 15381 5692
rect 15531 5732 15573 5741
rect 15531 5692 15532 5732
rect 15572 5692 15573 5732
rect 15531 5683 15573 5692
rect 15723 5732 15765 5741
rect 15723 5692 15724 5732
rect 15764 5692 15765 5732
rect 15723 5683 15765 5692
rect 15915 5732 15957 5741
rect 15915 5692 15916 5732
rect 15956 5692 15957 5732
rect 15915 5683 15957 5692
rect 16107 5732 16149 5741
rect 16107 5692 16108 5732
rect 16148 5692 16149 5732
rect 16107 5683 16149 5692
rect 16299 5732 16341 5741
rect 16299 5692 16300 5732
rect 16340 5692 16341 5732
rect 16299 5683 16341 5692
rect 16491 5732 16533 5741
rect 16491 5692 16492 5732
rect 16532 5692 16533 5732
rect 16491 5683 16533 5692
rect 16683 5732 16725 5741
rect 16683 5692 16684 5732
rect 16724 5692 16725 5732
rect 16683 5683 16725 5692
rect 16875 5732 16917 5741
rect 16875 5692 16876 5732
rect 16916 5692 16917 5732
rect 16875 5683 16917 5692
rect 17067 5732 17109 5741
rect 17067 5692 17068 5732
rect 17108 5692 17109 5732
rect 17067 5683 17109 5692
rect 17259 5732 17301 5741
rect 17259 5692 17260 5732
rect 17300 5692 17301 5732
rect 17259 5683 17301 5692
rect 17451 5732 17493 5741
rect 17451 5692 17452 5732
rect 17492 5692 17493 5732
rect 17451 5683 17493 5692
rect 18123 5732 18165 5741
rect 18123 5692 18124 5732
rect 18164 5692 18165 5732
rect 18123 5683 18165 5692
rect 18315 5732 18357 5741
rect 18315 5692 18316 5732
rect 18356 5692 18357 5732
rect 18315 5683 18357 5692
rect 18603 5732 18645 5741
rect 18603 5692 18604 5732
rect 18644 5692 18645 5732
rect 18603 5683 18645 5692
rect 18795 5732 18837 5741
rect 18795 5692 18796 5732
rect 18836 5692 18837 5732
rect 18795 5683 18837 5692
rect 18987 5732 19029 5741
rect 18987 5692 18988 5732
rect 19028 5692 19029 5732
rect 18987 5683 19029 5692
rect 19179 5732 19221 5741
rect 19179 5692 19180 5732
rect 19220 5692 19221 5732
rect 19179 5683 19221 5692
rect 19371 5732 19413 5741
rect 19371 5692 19372 5732
rect 19412 5692 19413 5732
rect 19371 5683 19413 5692
rect 19563 5732 19605 5741
rect 19563 5692 19564 5732
rect 19604 5692 19605 5732
rect 19563 5683 19605 5692
rect 19755 5732 19797 5741
rect 19755 5692 19756 5732
rect 19796 5692 19797 5732
rect 19755 5683 19797 5692
rect 19947 5732 19989 5741
rect 19947 5692 19948 5732
rect 19988 5692 19989 5732
rect 19947 5683 19989 5692
rect 20139 5732 20181 5741
rect 20139 5692 20140 5732
rect 20180 5692 20181 5732
rect 20139 5683 20181 5692
rect 20331 5732 20373 5741
rect 20331 5692 20332 5732
rect 20372 5692 20373 5732
rect 20331 5683 20373 5692
rect 20523 5732 20565 5741
rect 20523 5692 20524 5732
rect 20564 5692 20565 5732
rect 20523 5683 20565 5692
rect 20715 5732 20757 5741
rect 20715 5692 20716 5732
rect 20756 5692 20757 5732
rect 20715 5683 20757 5692
rect 22723 5732 22781 5733
rect 22723 5692 22732 5732
rect 22772 5692 22781 5732
rect 22723 5691 22781 5692
rect 23011 5732 23069 5733
rect 23011 5692 23020 5732
rect 23060 5692 23069 5732
rect 23011 5691 23069 5692
rect 23211 5732 23253 5741
rect 23211 5692 23212 5732
rect 23252 5692 23253 5732
rect 23211 5683 23253 5692
rect 23299 5732 23357 5733
rect 23299 5692 23308 5732
rect 23348 5692 23357 5732
rect 23299 5691 23357 5692
rect 23787 5732 23829 5741
rect 23787 5692 23788 5732
rect 23828 5692 23829 5732
rect 23787 5683 23829 5692
rect 23979 5732 24021 5741
rect 23979 5692 23980 5732
rect 24020 5692 24021 5732
rect 23979 5683 24021 5692
rect 24171 5732 24213 5741
rect 24171 5692 24172 5732
rect 24212 5692 24213 5732
rect 24171 5683 24213 5692
rect 24363 5732 24405 5741
rect 24363 5692 24364 5732
rect 24404 5692 24405 5732
rect 24363 5683 24405 5692
rect 24739 5732 24797 5733
rect 24739 5692 24748 5732
rect 24788 5692 24797 5732
rect 24739 5691 24797 5692
rect 24931 5732 24989 5733
rect 24931 5692 24940 5732
rect 24980 5692 24989 5732
rect 24931 5691 24989 5692
rect 26571 5732 26613 5741
rect 26571 5692 26572 5732
rect 26612 5692 26613 5732
rect 26571 5683 26613 5692
rect 26763 5732 26805 5741
rect 26763 5692 26764 5732
rect 26804 5692 26805 5732
rect 26763 5683 26805 5692
rect 26955 5732 26997 5741
rect 26955 5692 26956 5732
rect 26996 5692 26997 5732
rect 26955 5683 26997 5692
rect 27147 5732 27189 5741
rect 27147 5692 27148 5732
rect 27188 5692 27189 5732
rect 27147 5683 27189 5692
rect 28491 5732 28533 5741
rect 28491 5692 28492 5732
rect 28532 5692 28533 5732
rect 28491 5683 28533 5692
rect 28683 5732 28725 5741
rect 28683 5692 28684 5732
rect 28724 5692 28725 5732
rect 28683 5683 28725 5692
rect 28963 5732 29021 5733
rect 28963 5692 28972 5732
rect 29012 5692 29021 5732
rect 28963 5691 29021 5692
rect 29155 5732 29213 5733
rect 29155 5692 29164 5732
rect 29204 5692 29213 5732
rect 29155 5691 29213 5692
rect 30115 5732 30173 5733
rect 30115 5692 30124 5732
rect 30164 5692 30173 5732
rect 30115 5691 30173 5692
rect 30307 5732 30365 5733
rect 30307 5692 30316 5732
rect 30356 5692 30365 5732
rect 30307 5691 30365 5692
rect 30595 5732 30653 5733
rect 30595 5692 30604 5732
rect 30644 5692 30653 5732
rect 30595 5691 30653 5692
rect 30787 5732 30845 5733
rect 30787 5692 30796 5732
rect 30836 5692 30845 5732
rect 30787 5691 30845 5692
rect 31083 5732 31125 5741
rect 31083 5692 31084 5732
rect 31124 5692 31125 5732
rect 31083 5683 31125 5692
rect 31275 5732 31317 5741
rect 31275 5692 31276 5732
rect 31316 5692 31317 5732
rect 31275 5683 31317 5692
rect 31467 5732 31509 5741
rect 31467 5692 31468 5732
rect 31508 5692 31509 5732
rect 31467 5683 31509 5692
rect 31659 5732 31701 5741
rect 31659 5692 31660 5732
rect 31700 5692 31701 5732
rect 31659 5683 31701 5692
rect 31851 5732 31893 5741
rect 31851 5692 31852 5732
rect 31892 5692 31893 5732
rect 31851 5683 31893 5692
rect 32043 5732 32085 5741
rect 32043 5692 32044 5732
rect 32084 5692 32085 5732
rect 32043 5683 32085 5692
rect 32235 5732 32277 5741
rect 32235 5692 32236 5732
rect 32276 5692 32277 5732
rect 32235 5683 32277 5692
rect 32427 5732 32469 5741
rect 32427 5692 32428 5732
rect 32468 5692 32469 5732
rect 32427 5683 32469 5692
rect 32619 5732 32661 5741
rect 32619 5692 32620 5732
rect 32660 5692 32661 5732
rect 32619 5683 32661 5692
rect 32811 5732 32853 5741
rect 32811 5692 32812 5732
rect 32852 5692 32853 5732
rect 32811 5683 32853 5692
rect 34155 5732 34197 5741
rect 34155 5692 34156 5732
rect 34196 5692 34197 5732
rect 34155 5683 34197 5692
rect 34347 5732 34389 5741
rect 34347 5692 34348 5732
rect 34388 5692 34389 5732
rect 34347 5683 34389 5692
rect 34539 5732 34581 5741
rect 34539 5692 34540 5732
rect 34580 5692 34581 5732
rect 34539 5683 34581 5692
rect 34731 5732 34773 5741
rect 34731 5692 34732 5732
rect 34772 5692 34773 5732
rect 34731 5683 34773 5692
rect 34923 5732 34965 5741
rect 34923 5692 34924 5732
rect 34964 5692 34965 5732
rect 34923 5683 34965 5692
rect 35115 5732 35157 5741
rect 35115 5692 35116 5732
rect 35156 5692 35157 5732
rect 35115 5683 35157 5692
rect 35395 5732 35453 5733
rect 35395 5692 35404 5732
rect 35444 5692 35453 5732
rect 35395 5691 35453 5692
rect 35587 5732 35645 5733
rect 35587 5692 35596 5732
rect 35636 5692 35645 5732
rect 35587 5691 35645 5692
rect 36075 5732 36117 5741
rect 36075 5692 36076 5732
rect 36116 5692 36117 5732
rect 36075 5683 36117 5692
rect 36267 5732 36309 5741
rect 36267 5692 36268 5732
rect 36308 5692 36309 5732
rect 36267 5683 36309 5692
rect 36459 5732 36501 5741
rect 36459 5692 36460 5732
rect 36500 5692 36501 5732
rect 36459 5683 36501 5692
rect 36651 5732 36693 5741
rect 36651 5692 36652 5732
rect 36692 5692 36693 5732
rect 36651 5683 36693 5692
rect 36843 5732 36885 5741
rect 36843 5692 36844 5732
rect 36884 5692 36885 5732
rect 37035 5703 37036 5743
rect 37076 5703 37077 5743
rect 37035 5694 37077 5703
rect 37219 5732 37277 5733
rect 36843 5683 36885 5692
rect 37219 5692 37228 5732
rect 37268 5692 37277 5732
rect 37219 5691 37277 5692
rect 37515 5732 37557 5741
rect 37515 5692 37516 5732
rect 37556 5692 37557 5732
rect 37515 5683 37557 5692
rect 37707 5732 37749 5741
rect 37707 5692 37708 5732
rect 37748 5692 37749 5732
rect 37707 5683 37749 5692
rect 37899 5732 37941 5741
rect 37899 5692 37900 5732
rect 37940 5692 37941 5732
rect 37899 5683 37941 5692
rect 38091 5732 38133 5741
rect 38091 5692 38092 5732
rect 38132 5692 38133 5732
rect 38091 5683 38133 5692
rect 38563 5732 38621 5733
rect 38563 5692 38572 5732
rect 38612 5692 38621 5732
rect 38563 5691 38621 5692
rect 38755 5732 38813 5733
rect 38755 5692 38764 5732
rect 38804 5692 38813 5732
rect 38755 5691 38813 5692
rect 39147 5732 39189 5741
rect 39147 5692 39148 5732
rect 39188 5692 39189 5732
rect 39147 5683 39189 5692
rect 39339 5732 39381 5741
rect 39339 5692 39340 5732
rect 39380 5692 39381 5732
rect 39339 5683 39381 5692
rect 42595 5732 42653 5733
rect 42595 5692 42604 5732
rect 42644 5692 42653 5732
rect 42595 5691 42653 5692
rect 44035 5732 44093 5733
rect 44035 5692 44044 5732
rect 44084 5692 44093 5732
rect 44035 5691 44093 5692
rect 44235 5732 44277 5741
rect 44235 5692 44236 5732
rect 44276 5692 44277 5732
rect 44235 5683 44277 5692
rect 44323 5732 44381 5733
rect 44323 5692 44332 5732
rect 44372 5692 44381 5732
rect 44323 5691 44381 5692
rect 44515 5732 44573 5733
rect 44515 5692 44524 5732
rect 44564 5692 44573 5732
rect 44515 5691 44573 5692
rect 44715 5732 44757 5741
rect 44715 5692 44716 5732
rect 44756 5692 44757 5732
rect 44715 5683 44757 5692
rect 44803 5732 44861 5733
rect 44803 5692 44812 5732
rect 44852 5692 44861 5732
rect 44803 5691 44861 5692
rect 45091 5732 45149 5733
rect 45091 5692 45100 5732
rect 45140 5692 45149 5732
rect 45091 5691 45149 5692
rect 45195 5732 45237 5741
rect 45195 5692 45196 5732
rect 45236 5692 45237 5732
rect 45195 5683 45237 5692
rect 45379 5732 45437 5733
rect 45379 5692 45388 5732
rect 45428 5692 45437 5732
rect 45379 5691 45437 5692
rect 45667 5732 45725 5733
rect 45667 5692 45676 5732
rect 45716 5692 45725 5732
rect 45667 5691 45725 5692
rect 46627 5732 46685 5733
rect 46627 5692 46636 5732
rect 46676 5692 46685 5732
rect 46627 5691 46685 5692
rect 48643 5732 48701 5733
rect 48643 5692 48652 5732
rect 48692 5692 48701 5732
rect 48643 5691 48701 5692
rect 49603 5732 49661 5733
rect 49603 5692 49612 5732
rect 49652 5692 49661 5732
rect 49603 5691 49661 5692
rect 52195 5732 52253 5733
rect 52195 5692 52204 5732
rect 52244 5692 52253 5732
rect 52195 5691 52253 5692
rect 52395 5732 52437 5741
rect 52395 5692 52396 5732
rect 52436 5692 52437 5732
rect 52395 5683 52437 5692
rect 52483 5732 52541 5733
rect 52483 5692 52492 5732
rect 52532 5692 52541 5732
rect 52483 5691 52541 5692
rect 53739 5732 53781 5741
rect 53739 5692 53740 5732
rect 53780 5692 53781 5732
rect 53739 5683 53781 5692
rect 53931 5732 53973 5741
rect 53931 5692 53932 5732
rect 53972 5692 53973 5732
rect 53931 5683 53973 5692
rect 54315 5732 54357 5741
rect 54315 5692 54316 5732
rect 54356 5692 54357 5732
rect 54315 5683 54357 5692
rect 54507 5732 54549 5741
rect 54507 5692 54508 5732
rect 54548 5692 54549 5732
rect 54507 5683 54549 5692
rect 55659 5732 55701 5741
rect 55659 5692 55660 5732
rect 55700 5692 55701 5732
rect 55659 5683 55701 5692
rect 55755 5732 55797 5741
rect 55755 5692 55756 5732
rect 55796 5692 55797 5732
rect 55755 5683 55797 5692
rect 55843 5732 55901 5733
rect 55843 5692 55852 5732
rect 55892 5692 55901 5732
rect 55843 5691 55901 5692
rect 56331 5732 56373 5741
rect 56331 5692 56332 5732
rect 56372 5692 56373 5732
rect 56331 5683 56373 5692
rect 56523 5732 56565 5741
rect 56523 5692 56524 5732
rect 56564 5692 56565 5732
rect 56523 5683 56565 5692
rect 56715 5732 56757 5741
rect 56715 5692 56716 5732
rect 56756 5692 56757 5732
rect 56715 5683 56757 5692
rect 56907 5732 56949 5741
rect 56907 5692 56908 5732
rect 56948 5692 56949 5732
rect 56907 5683 56949 5692
rect 57291 5732 57333 5741
rect 57291 5692 57292 5732
rect 57332 5692 57333 5732
rect 57291 5683 57333 5692
rect 57675 5740 57717 5749
rect 57675 5700 57676 5740
rect 57716 5700 57717 5740
rect 57675 5691 57717 5700
rect 58251 5732 58293 5741
rect 58251 5692 58252 5732
rect 58292 5692 58293 5732
rect 58251 5683 58293 5692
rect 61227 5732 61269 5741
rect 61227 5692 61228 5732
rect 61268 5692 61269 5732
rect 61227 5683 61269 5692
rect 61323 5732 61365 5741
rect 61323 5692 61324 5732
rect 61364 5692 61365 5732
rect 61323 5683 61365 5692
rect 61995 5732 62037 5741
rect 61995 5692 61996 5732
rect 62036 5692 62037 5732
rect 61995 5683 62037 5692
rect 64579 5732 64637 5733
rect 64579 5692 64588 5732
rect 64628 5692 64637 5732
rect 64579 5691 64637 5692
rect 67267 5732 67325 5733
rect 67267 5692 67276 5732
rect 67316 5692 67325 5732
rect 67267 5691 67325 5692
rect 67459 5732 67517 5733
rect 67459 5692 67468 5732
rect 67508 5692 67517 5732
rect 67459 5691 67517 5692
rect 68331 5732 68373 5741
rect 68331 5692 68332 5732
rect 68372 5692 68373 5732
rect 68331 5683 68373 5692
rect 68523 5732 68565 5741
rect 68523 5692 68524 5732
rect 68564 5692 68565 5732
rect 68523 5683 68565 5692
rect 68715 5732 68757 5741
rect 68715 5692 68716 5732
rect 68756 5692 68757 5732
rect 68715 5683 68757 5692
rect 68907 5732 68949 5741
rect 68907 5692 68908 5732
rect 68948 5692 68949 5732
rect 68907 5683 68949 5692
rect 69579 5732 69621 5741
rect 69579 5692 69580 5732
rect 69620 5692 69621 5732
rect 69579 5683 69621 5692
rect 69771 5732 69813 5741
rect 69771 5692 69772 5732
rect 69812 5692 69813 5732
rect 69771 5683 69813 5692
rect 71299 5732 71357 5733
rect 71299 5692 71308 5732
rect 71348 5692 71357 5732
rect 71299 5691 71357 5692
rect 71491 5732 71549 5733
rect 71491 5692 71500 5732
rect 71540 5692 71549 5732
rect 71491 5691 71549 5692
rect 71979 5732 72021 5741
rect 71979 5692 71980 5732
rect 72020 5692 72021 5732
rect 71979 5683 72021 5692
rect 72171 5732 72213 5741
rect 72171 5692 72172 5732
rect 72212 5692 72213 5732
rect 72171 5683 72213 5692
rect 72363 5732 72405 5741
rect 72363 5692 72364 5732
rect 72404 5692 72405 5732
rect 72363 5683 72405 5692
rect 72555 5732 72597 5741
rect 72555 5692 72556 5732
rect 72596 5692 72597 5732
rect 72555 5683 72597 5692
rect 72747 5732 72789 5741
rect 72747 5692 72748 5732
rect 72788 5692 72789 5732
rect 72747 5683 72789 5692
rect 72939 5732 72981 5741
rect 72939 5692 72940 5732
rect 72980 5692 72981 5732
rect 72939 5683 72981 5692
rect 73419 5732 73461 5741
rect 73419 5692 73420 5732
rect 73460 5692 73461 5732
rect 73419 5683 73461 5692
rect 73611 5732 73653 5741
rect 73611 5692 73612 5732
rect 73652 5692 73653 5732
rect 73611 5683 73653 5692
rect 73803 5732 73845 5741
rect 73803 5692 73804 5732
rect 73844 5692 73845 5732
rect 73803 5683 73845 5692
rect 73995 5732 74037 5741
rect 73995 5692 73996 5732
rect 74036 5692 74037 5732
rect 73995 5683 74037 5692
rect 74275 5732 74333 5733
rect 74275 5692 74284 5732
rect 74324 5692 74333 5732
rect 74275 5691 74333 5692
rect 74467 5732 74525 5733
rect 74467 5692 74476 5732
rect 74516 5692 74525 5732
rect 74467 5691 74525 5692
rect 74955 5732 74997 5741
rect 74955 5692 74956 5732
rect 74996 5692 74997 5732
rect 74955 5683 74997 5692
rect 75051 5732 75093 5741
rect 75051 5692 75052 5732
rect 75092 5692 75093 5732
rect 75051 5683 75093 5692
rect 75723 5732 75765 5741
rect 75723 5692 75724 5732
rect 75764 5692 75765 5732
rect 75723 5683 75765 5692
rect 75915 5732 75957 5741
rect 75915 5692 75916 5732
rect 75956 5692 75957 5732
rect 75915 5683 75957 5692
rect 77259 5732 77301 5741
rect 77259 5692 77260 5732
rect 77300 5692 77301 5732
rect 77259 5683 77301 5692
rect 77451 5732 77493 5741
rect 77451 5692 77452 5732
rect 77492 5692 77493 5732
rect 77451 5683 77493 5692
rect 78027 5732 78069 5741
rect 78027 5692 78028 5732
rect 78068 5692 78069 5732
rect 78027 5683 78069 5692
rect 78507 5732 78549 5741
rect 78507 5692 78508 5732
rect 78548 5692 78549 5732
rect 78507 5683 78549 5692
rect 78699 5732 78741 5741
rect 78699 5692 78700 5732
rect 78740 5692 78741 5732
rect 78699 5683 78741 5692
rect 78891 5732 78933 5741
rect 78891 5692 78892 5732
rect 78932 5692 78933 5732
rect 78891 5683 78933 5692
rect 79083 5732 79125 5741
rect 79083 5692 79084 5732
rect 79124 5692 79125 5732
rect 79083 5683 79125 5692
rect 79275 5732 79317 5741
rect 79275 5692 79276 5732
rect 79316 5692 79317 5732
rect 79275 5683 79317 5692
rect 79467 5732 79509 5741
rect 79467 5692 79468 5732
rect 79508 5692 79509 5732
rect 79467 5683 79509 5692
rect 79659 5732 79701 5741
rect 79659 5692 79660 5732
rect 79700 5692 79701 5732
rect 79659 5683 79701 5692
rect 79851 5732 79893 5741
rect 79851 5692 79852 5732
rect 79892 5692 79893 5732
rect 79851 5683 79893 5692
rect 80043 5732 80085 5741
rect 80043 5692 80044 5732
rect 80084 5692 80085 5732
rect 80043 5683 80085 5692
rect 80235 5732 80277 5741
rect 80235 5692 80236 5732
rect 80276 5692 80277 5732
rect 80235 5683 80277 5692
rect 80427 5732 80469 5741
rect 80427 5692 80428 5732
rect 80468 5692 80469 5732
rect 80427 5683 80469 5692
rect 80619 5732 80661 5741
rect 80619 5692 80620 5732
rect 80660 5692 80661 5732
rect 80619 5683 80661 5692
rect 80907 5732 80949 5741
rect 80907 5692 80908 5732
rect 80948 5692 80949 5732
rect 80907 5683 80949 5692
rect 81099 5732 81141 5741
rect 81099 5692 81100 5732
rect 81140 5692 81141 5732
rect 81099 5683 81141 5692
rect 81291 5732 81333 5741
rect 81291 5692 81292 5732
rect 81332 5692 81333 5732
rect 81291 5683 81333 5692
rect 81483 5732 81525 5741
rect 81483 5692 81484 5732
rect 81524 5692 81525 5732
rect 81483 5683 81525 5692
rect 81675 5732 81717 5741
rect 81675 5692 81676 5732
rect 81716 5692 81717 5732
rect 81675 5683 81717 5692
rect 81867 5732 81909 5741
rect 81867 5692 81868 5732
rect 81908 5692 81909 5732
rect 81867 5683 81909 5692
rect 82155 5732 82197 5741
rect 82155 5692 82156 5732
rect 82196 5692 82197 5732
rect 82155 5683 82197 5692
rect 82347 5732 82389 5741
rect 82347 5692 82348 5732
rect 82388 5692 82389 5732
rect 82347 5683 82389 5692
rect 82539 5732 82581 5741
rect 82539 5692 82540 5732
rect 82580 5692 82581 5732
rect 82539 5683 82581 5692
rect 82731 5732 82773 5741
rect 82731 5692 82732 5732
rect 82772 5692 82773 5732
rect 82731 5683 82773 5692
rect 82923 5732 82965 5741
rect 82923 5692 82924 5732
rect 82964 5692 82965 5732
rect 82923 5683 82965 5692
rect 83115 5732 83157 5741
rect 83115 5692 83116 5732
rect 83156 5692 83157 5732
rect 83115 5683 83157 5692
rect 83307 5732 83349 5741
rect 83307 5692 83308 5732
rect 83348 5692 83349 5732
rect 83307 5683 83349 5692
rect 83499 5732 83541 5741
rect 83499 5692 83500 5732
rect 83540 5692 83541 5732
rect 83499 5683 83541 5692
rect 83691 5732 83733 5741
rect 83691 5692 83692 5732
rect 83732 5692 83733 5732
rect 83691 5683 83733 5692
rect 83883 5732 83925 5741
rect 83883 5692 83884 5732
rect 83924 5692 83925 5732
rect 83883 5683 83925 5692
rect 84555 5732 84597 5741
rect 84555 5692 84556 5732
rect 84596 5692 84597 5732
rect 84555 5683 84597 5692
rect 70147 5661 70205 5662
rect 1699 5648 1757 5649
rect 1699 5608 1708 5648
rect 1748 5608 1757 5648
rect 1699 5607 1757 5608
rect 2083 5648 2141 5649
rect 2083 5608 2092 5648
rect 2132 5608 2141 5648
rect 2083 5607 2141 5608
rect 17731 5648 17789 5649
rect 17731 5608 17740 5648
rect 17780 5608 17789 5648
rect 17731 5607 17789 5608
rect 19083 5648 19125 5657
rect 19083 5608 19084 5648
rect 19124 5608 19125 5648
rect 19083 5599 19125 5608
rect 20235 5648 20277 5657
rect 20235 5608 20236 5648
rect 20276 5608 20277 5648
rect 20235 5599 20277 5608
rect 20995 5648 21053 5649
rect 20995 5608 21004 5648
rect 21044 5608 21053 5648
rect 20995 5607 21053 5608
rect 21379 5648 21437 5649
rect 21379 5608 21388 5648
rect 21428 5608 21437 5648
rect 21379 5607 21437 5608
rect 28099 5648 28157 5649
rect 28099 5608 28108 5648
rect 28148 5608 28157 5648
rect 28099 5607 28157 5608
rect 29539 5648 29597 5649
rect 29539 5608 29548 5648
rect 29588 5608 29597 5648
rect 29539 5607 29597 5608
rect 29923 5648 29981 5649
rect 29923 5608 29932 5648
rect 29972 5608 29981 5648
rect 29923 5607 29981 5608
rect 33763 5648 33821 5649
rect 33763 5608 33772 5648
rect 33812 5608 33821 5648
rect 33763 5607 33821 5608
rect 39243 5648 39285 5657
rect 39243 5608 39244 5648
rect 39284 5608 39285 5648
rect 39243 5599 39285 5608
rect 39715 5648 39773 5649
rect 39715 5608 39724 5648
rect 39764 5608 39773 5648
rect 39715 5607 39773 5608
rect 40099 5648 40157 5649
rect 40099 5608 40108 5648
rect 40148 5608 40157 5648
rect 40099 5607 40157 5608
rect 41251 5648 41309 5649
rect 41251 5608 41260 5648
rect 41300 5608 41309 5648
rect 41251 5607 41309 5608
rect 42883 5648 42941 5649
rect 42883 5608 42892 5648
rect 42932 5608 42941 5648
rect 42883 5607 42941 5608
rect 43267 5648 43325 5649
rect 43267 5608 43276 5648
rect 43316 5608 43325 5648
rect 43267 5607 43325 5608
rect 43651 5648 43709 5649
rect 43651 5608 43660 5648
rect 43700 5608 43709 5648
rect 43651 5607 43709 5608
rect 47107 5648 47165 5649
rect 47107 5608 47116 5648
rect 47156 5608 47165 5648
rect 47107 5607 47165 5608
rect 47491 5648 47549 5649
rect 47491 5608 47500 5648
rect 47540 5608 47549 5648
rect 47491 5607 47549 5608
rect 47875 5648 47933 5649
rect 47875 5608 47884 5648
rect 47924 5608 47933 5648
rect 47875 5607 47933 5608
rect 48259 5648 48317 5649
rect 48259 5608 48268 5648
rect 48308 5608 48317 5648
rect 48259 5607 48317 5608
rect 50083 5648 50141 5649
rect 50083 5608 50092 5648
rect 50132 5608 50141 5648
rect 50083 5607 50141 5608
rect 53155 5648 53213 5649
rect 53155 5608 53164 5648
rect 53204 5608 53213 5648
rect 53155 5607 53213 5608
rect 54883 5648 54941 5649
rect 54883 5608 54892 5648
rect 54932 5608 54941 5648
rect 54883 5607 54941 5608
rect 55267 5648 55325 5649
rect 55267 5608 55276 5648
rect 55316 5608 55325 5648
rect 55267 5607 55325 5608
rect 58723 5648 58781 5649
rect 58723 5608 58732 5648
rect 58772 5608 58781 5648
rect 58723 5607 58781 5608
rect 59107 5648 59165 5649
rect 59107 5608 59116 5648
rect 59156 5608 59165 5648
rect 59107 5607 59165 5608
rect 59491 5648 59549 5649
rect 59491 5608 59500 5648
rect 59540 5608 59549 5648
rect 59491 5607 59549 5608
rect 59875 5648 59933 5649
rect 59875 5608 59884 5648
rect 59924 5608 59933 5648
rect 59875 5607 59933 5608
rect 60259 5648 60317 5649
rect 60259 5608 60268 5648
rect 60308 5608 60317 5648
rect 60259 5607 60317 5608
rect 60643 5648 60701 5649
rect 60643 5608 60652 5648
rect 60692 5608 60701 5648
rect 60643 5607 60701 5608
rect 61803 5648 61845 5657
rect 61803 5608 61804 5648
rect 61844 5608 61845 5648
rect 61803 5599 61845 5608
rect 62467 5648 62525 5649
rect 62467 5608 62476 5648
rect 62516 5608 62525 5648
rect 62467 5607 62525 5608
rect 62851 5648 62909 5649
rect 62851 5608 62860 5648
rect 62900 5608 62909 5648
rect 62851 5607 62909 5608
rect 63235 5648 63293 5649
rect 63235 5608 63244 5648
rect 63284 5608 63293 5648
rect 63235 5607 63293 5608
rect 63619 5648 63677 5649
rect 63619 5608 63628 5648
rect 63668 5608 63677 5648
rect 63619 5607 63677 5608
rect 64003 5648 64061 5649
rect 64003 5608 64012 5648
rect 64052 5608 64061 5648
rect 64003 5607 64061 5608
rect 66979 5648 67037 5649
rect 66979 5608 66988 5648
rect 67028 5608 67037 5648
rect 66979 5607 67037 5608
rect 67843 5648 67901 5649
rect 67843 5608 67852 5648
rect 67892 5608 67901 5648
rect 67843 5607 67901 5608
rect 68811 5648 68853 5657
rect 68811 5608 68812 5648
rect 68852 5608 68853 5648
rect 68811 5599 68853 5608
rect 69283 5648 69341 5649
rect 69283 5608 69292 5648
rect 69332 5608 69341 5648
rect 70147 5621 70156 5661
rect 70196 5621 70205 5661
rect 86589 5661 86631 5670
rect 70147 5620 70205 5621
rect 70531 5648 70589 5649
rect 69283 5607 69341 5608
rect 70531 5608 70540 5648
rect 70580 5608 70589 5648
rect 70531 5607 70589 5608
rect 70915 5648 70973 5649
rect 70915 5608 70924 5648
rect 70964 5608 70973 5648
rect 70915 5607 70973 5608
rect 73515 5648 73557 5657
rect 73515 5608 73516 5648
rect 73556 5608 73557 5648
rect 73515 5599 73557 5608
rect 74859 5648 74901 5657
rect 74859 5608 74860 5648
rect 74900 5608 74901 5648
rect 74859 5599 74901 5608
rect 75523 5648 75581 5649
rect 75523 5608 75532 5648
rect 75572 5608 75581 5648
rect 75523 5607 75581 5608
rect 76291 5648 76349 5649
rect 76291 5608 76300 5648
rect 76340 5608 76349 5648
rect 76291 5607 76349 5608
rect 76675 5648 76733 5649
rect 76675 5608 76684 5648
rect 76724 5608 76733 5648
rect 76675 5607 76733 5608
rect 77059 5648 77117 5649
rect 77059 5608 77068 5648
rect 77108 5608 77117 5648
rect 77059 5607 77117 5608
rect 77835 5648 77877 5657
rect 77835 5608 77836 5648
rect 77876 5608 77877 5648
rect 77835 5599 77877 5608
rect 82635 5648 82677 5657
rect 82635 5608 82636 5648
rect 82676 5608 82677 5648
rect 82635 5599 82677 5608
rect 84363 5648 84405 5657
rect 84363 5608 84364 5648
rect 84404 5608 84405 5648
rect 84363 5599 84405 5608
rect 85027 5648 85085 5649
rect 85027 5608 85036 5648
rect 85076 5608 85085 5648
rect 85027 5607 85085 5608
rect 85411 5648 85469 5649
rect 85411 5608 85420 5648
rect 85460 5608 85469 5648
rect 85411 5607 85469 5608
rect 85795 5648 85853 5649
rect 85795 5608 85804 5648
rect 85844 5608 85853 5648
rect 85795 5607 85853 5608
rect 86179 5648 86237 5649
rect 86179 5608 86188 5648
rect 86228 5608 86237 5648
rect 86589 5621 86590 5661
rect 86630 5621 86631 5661
rect 86589 5612 86631 5621
rect 97507 5648 97565 5649
rect 86179 5607 86237 5608
rect 97507 5608 97516 5648
rect 97556 5608 97565 5648
rect 97507 5607 97565 5608
rect 97891 5648 97949 5649
rect 97891 5608 97900 5648
rect 97940 5608 97949 5648
rect 97891 5607 97949 5608
rect 98467 5648 98525 5649
rect 98467 5608 98476 5648
rect 98516 5608 98525 5648
rect 98467 5607 98525 5608
rect 57291 5590 57333 5599
rect 17259 5564 17301 5573
rect 17259 5524 17260 5564
rect 17300 5524 17301 5564
rect 17259 5515 17301 5524
rect 19755 5564 19797 5573
rect 19755 5524 19756 5564
rect 19796 5524 19797 5564
rect 19755 5515 19797 5524
rect 56523 5564 56565 5573
rect 56523 5524 56524 5564
rect 56564 5524 56565 5564
rect 57291 5550 57292 5590
rect 57332 5550 57333 5590
rect 57291 5541 57333 5550
rect 57675 5564 57717 5573
rect 56523 5515 56565 5524
rect 57675 5524 57676 5564
rect 57716 5524 57717 5564
rect 57675 5515 57717 5524
rect 57867 5564 57909 5573
rect 57867 5524 57868 5564
rect 57908 5524 57909 5564
rect 57867 5515 57909 5524
rect 58251 5564 58293 5573
rect 58251 5524 58252 5564
rect 58292 5524 58293 5564
rect 58251 5515 58293 5524
rect 61899 5564 61941 5573
rect 61899 5524 61900 5564
rect 61940 5524 61941 5564
rect 61899 5515 61941 5524
rect 63819 5564 63861 5573
rect 63819 5524 63820 5564
rect 63860 5524 63861 5564
rect 63819 5515 63861 5524
rect 74475 5564 74517 5573
rect 74475 5524 74476 5564
rect 74516 5524 74517 5564
rect 74475 5515 74517 5524
rect 75915 5564 75957 5573
rect 75915 5524 75916 5564
rect 75956 5524 75957 5564
rect 75915 5515 75957 5524
rect 79083 5564 79125 5573
rect 79083 5524 79084 5564
rect 79124 5524 79125 5564
rect 79083 5515 79125 5524
rect 83883 5564 83925 5573
rect 83883 5524 83884 5564
rect 83924 5524 83925 5564
rect 83883 5515 83925 5524
rect 1515 5480 1557 5489
rect 1515 5440 1516 5480
rect 1556 5440 1557 5480
rect 1515 5431 1557 5440
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 15339 5480 15381 5489
rect 15339 5440 15340 5480
rect 15380 5440 15381 5480
rect 15339 5431 15381 5440
rect 15723 5480 15765 5489
rect 15723 5440 15724 5480
rect 15764 5440 15765 5480
rect 15723 5431 15765 5440
rect 16107 5480 16149 5489
rect 16107 5440 16108 5480
rect 16148 5440 16149 5480
rect 16107 5431 16149 5440
rect 16491 5480 16533 5489
rect 16491 5440 16492 5480
rect 16532 5440 16533 5480
rect 16491 5431 16533 5440
rect 17931 5480 17973 5489
rect 17931 5440 17932 5480
rect 17972 5440 17973 5480
rect 17931 5431 17973 5440
rect 18123 5480 18165 5489
rect 18123 5440 18124 5480
rect 18164 5440 18165 5480
rect 18123 5431 18165 5440
rect 18603 5480 18645 5489
rect 18603 5440 18604 5480
rect 18644 5440 18645 5480
rect 18603 5431 18645 5440
rect 19371 5480 19413 5489
rect 19371 5440 19372 5480
rect 19412 5440 19413 5480
rect 19371 5431 19413 5440
rect 20523 5480 20565 5489
rect 20523 5440 20524 5480
rect 20564 5440 20565 5480
rect 20523 5431 20565 5440
rect 21195 5480 21237 5489
rect 21195 5440 21196 5480
rect 21236 5440 21237 5480
rect 21195 5431 21237 5440
rect 21579 5480 21621 5489
rect 21579 5440 21580 5480
rect 21620 5440 21621 5480
rect 21579 5431 21621 5440
rect 22443 5480 22485 5489
rect 22443 5440 22444 5480
rect 22484 5440 22485 5480
rect 22443 5431 22485 5440
rect 23787 5480 23829 5489
rect 23787 5440 23788 5480
rect 23828 5440 23829 5480
rect 23787 5431 23829 5440
rect 24171 5480 24213 5489
rect 24171 5440 24172 5480
rect 24212 5440 24213 5480
rect 24171 5431 24213 5440
rect 26763 5480 26805 5489
rect 26763 5440 26764 5480
rect 26804 5440 26805 5480
rect 26763 5431 26805 5440
rect 27147 5480 27189 5489
rect 27147 5440 27148 5480
rect 27188 5440 27189 5480
rect 27147 5431 27189 5440
rect 28299 5480 28341 5489
rect 28299 5440 28300 5480
rect 28340 5440 28341 5480
rect 28299 5431 28341 5440
rect 28491 5480 28533 5489
rect 28491 5440 28492 5480
rect 28532 5440 28533 5480
rect 28491 5431 28533 5440
rect 29355 5480 29397 5489
rect 29355 5440 29356 5480
rect 29396 5440 29397 5480
rect 29355 5431 29397 5440
rect 29739 5480 29781 5489
rect 29739 5440 29740 5480
rect 29780 5440 29781 5480
rect 29739 5431 29781 5440
rect 31083 5480 31125 5489
rect 31083 5440 31084 5480
rect 31124 5440 31125 5480
rect 31083 5431 31125 5440
rect 31659 5480 31701 5489
rect 31659 5440 31660 5480
rect 31700 5440 31701 5480
rect 31659 5431 31701 5440
rect 32043 5480 32085 5489
rect 32043 5440 32044 5480
rect 32084 5440 32085 5480
rect 32043 5431 32085 5440
rect 32427 5480 32469 5489
rect 32427 5440 32428 5480
rect 32468 5440 32469 5480
rect 32427 5431 32469 5440
rect 32811 5480 32853 5489
rect 32811 5440 32812 5480
rect 32852 5440 32853 5480
rect 32811 5431 32853 5440
rect 33963 5480 34005 5489
rect 33963 5440 33964 5480
rect 34004 5440 34005 5480
rect 33963 5431 34005 5440
rect 34347 5480 34389 5489
rect 34347 5440 34348 5480
rect 34388 5440 34389 5480
rect 34347 5431 34389 5440
rect 34731 5480 34773 5489
rect 34731 5440 34732 5480
rect 34772 5440 34773 5480
rect 34731 5431 34773 5440
rect 35115 5480 35157 5489
rect 35115 5440 35116 5480
rect 35156 5440 35157 5480
rect 35115 5431 35157 5440
rect 36267 5480 36309 5489
rect 36267 5440 36268 5480
rect 36308 5440 36309 5480
rect 36267 5431 36309 5440
rect 36651 5480 36693 5489
rect 36651 5440 36652 5480
rect 36692 5440 36693 5480
rect 36651 5431 36693 5440
rect 37035 5480 37077 5489
rect 37035 5440 37036 5480
rect 37076 5440 37077 5480
rect 37035 5431 37077 5440
rect 37323 5480 37365 5489
rect 37323 5440 37324 5480
rect 37364 5440 37365 5480
rect 37323 5431 37365 5440
rect 37707 5480 37749 5489
rect 37707 5440 37708 5480
rect 37748 5440 37749 5480
rect 37707 5431 37749 5440
rect 38091 5480 38133 5489
rect 38091 5440 38092 5480
rect 38132 5440 38133 5480
rect 38091 5431 38133 5440
rect 39531 5480 39573 5489
rect 39531 5440 39532 5480
rect 39572 5440 39573 5480
rect 39531 5431 39573 5440
rect 39915 5480 39957 5489
rect 39915 5440 39916 5480
rect 39956 5440 39957 5480
rect 39915 5431 39957 5440
rect 41067 5480 41109 5489
rect 41067 5440 41068 5480
rect 41108 5440 41109 5480
rect 41067 5431 41109 5440
rect 43083 5480 43125 5489
rect 43083 5440 43084 5480
rect 43124 5440 43125 5480
rect 43083 5431 43125 5440
rect 43467 5480 43509 5489
rect 43467 5440 43468 5480
rect 43508 5440 43509 5480
rect 43467 5431 43509 5440
rect 43851 5480 43893 5489
rect 43851 5440 43852 5480
rect 43892 5440 43893 5480
rect 43851 5431 43893 5440
rect 44235 5480 44277 5489
rect 44235 5440 44236 5480
rect 44276 5440 44277 5480
rect 44235 5431 44277 5440
rect 44523 5480 44565 5489
rect 44523 5440 44524 5480
rect 44564 5440 44565 5480
rect 44523 5431 44565 5440
rect 47307 5480 47349 5489
rect 47307 5440 47308 5480
rect 47348 5440 47349 5480
rect 47307 5431 47349 5440
rect 47691 5480 47733 5489
rect 47691 5440 47692 5480
rect 47732 5440 47733 5480
rect 47691 5431 47733 5440
rect 48075 5480 48117 5489
rect 48075 5440 48076 5480
rect 48116 5440 48117 5480
rect 48075 5431 48117 5440
rect 48459 5480 48501 5489
rect 48459 5440 48460 5480
rect 48500 5440 48501 5480
rect 48459 5431 48501 5440
rect 49899 5480 49941 5489
rect 49899 5440 49900 5480
rect 49940 5440 49941 5480
rect 49899 5431 49941 5440
rect 52203 5480 52245 5489
rect 52203 5440 52204 5480
rect 52244 5440 52245 5480
rect 52203 5431 52245 5440
rect 53931 5480 53973 5489
rect 53931 5440 53932 5480
rect 53972 5440 53973 5480
rect 53931 5431 53973 5440
rect 54315 5480 54357 5489
rect 54315 5440 54316 5480
rect 54356 5440 54357 5480
rect 54315 5431 54357 5440
rect 54699 5480 54741 5489
rect 54699 5440 54700 5480
rect 54740 5440 54741 5480
rect 54699 5431 54741 5440
rect 55083 5480 55125 5489
rect 55083 5440 55084 5480
rect 55124 5440 55125 5480
rect 55083 5431 55125 5440
rect 57099 5480 57141 5489
rect 57099 5440 57100 5480
rect 57140 5440 57141 5480
rect 57099 5431 57141 5440
rect 58059 5480 58101 5489
rect 58059 5440 58060 5480
rect 58100 5440 58101 5480
rect 58059 5431 58101 5440
rect 58539 5480 58581 5489
rect 58539 5440 58540 5480
rect 58580 5440 58581 5480
rect 58539 5431 58581 5440
rect 58923 5480 58965 5489
rect 58923 5440 58924 5480
rect 58964 5440 58965 5480
rect 58923 5431 58965 5440
rect 59307 5480 59349 5489
rect 59307 5440 59308 5480
rect 59348 5440 59349 5480
rect 59307 5431 59349 5440
rect 59691 5480 59733 5489
rect 59691 5440 59692 5480
rect 59732 5440 59733 5480
rect 59691 5431 59733 5440
rect 60075 5480 60117 5489
rect 60075 5440 60076 5480
rect 60116 5440 60117 5480
rect 60075 5431 60117 5440
rect 60459 5480 60501 5489
rect 60459 5440 60460 5480
rect 60500 5440 60501 5480
rect 60459 5431 60501 5440
rect 61035 5480 61077 5489
rect 61035 5440 61036 5480
rect 61076 5440 61077 5480
rect 61035 5431 61077 5440
rect 62283 5480 62325 5489
rect 62283 5440 62284 5480
rect 62324 5440 62325 5480
rect 62283 5431 62325 5440
rect 62667 5480 62709 5489
rect 62667 5440 62668 5480
rect 62708 5440 62709 5480
rect 62667 5431 62709 5440
rect 63051 5480 63093 5489
rect 63051 5440 63052 5480
rect 63092 5440 63093 5480
rect 63051 5431 63093 5440
rect 63435 5480 63477 5489
rect 63435 5440 63436 5480
rect 63476 5440 63477 5480
rect 63435 5431 63477 5440
rect 66795 5480 66837 5489
rect 66795 5440 66796 5480
rect 66836 5440 66837 5480
rect 66795 5431 66837 5440
rect 67659 5480 67701 5489
rect 67659 5440 67660 5480
rect 67700 5440 67701 5480
rect 67659 5431 67701 5440
rect 68331 5480 68373 5489
rect 68331 5440 68332 5480
rect 68372 5440 68373 5480
rect 68331 5431 68373 5440
rect 69099 5480 69141 5489
rect 69099 5440 69100 5480
rect 69140 5440 69141 5480
rect 69099 5431 69141 5440
rect 69771 5480 69813 5489
rect 69771 5440 69772 5480
rect 69812 5440 69813 5480
rect 69771 5431 69813 5440
rect 69963 5480 70005 5489
rect 69963 5440 69964 5480
rect 70004 5440 70005 5480
rect 69963 5431 70005 5440
rect 70347 5480 70389 5489
rect 70347 5440 70348 5480
rect 70388 5440 70389 5480
rect 70347 5431 70389 5440
rect 70731 5480 70773 5489
rect 70731 5440 70732 5480
rect 70772 5440 70773 5480
rect 70731 5431 70773 5440
rect 72555 5480 72597 5489
rect 72555 5440 72556 5480
rect 72596 5440 72597 5480
rect 72555 5431 72597 5440
rect 72939 5480 72981 5489
rect 72939 5440 72940 5480
rect 72980 5440 72981 5480
rect 72939 5431 72981 5440
rect 73995 5480 74037 5489
rect 73995 5440 73996 5480
rect 74036 5440 74037 5480
rect 73995 5431 74037 5440
rect 75339 5480 75381 5489
rect 75339 5440 75340 5480
rect 75380 5440 75381 5480
rect 75339 5431 75381 5440
rect 76107 5480 76149 5489
rect 76107 5440 76108 5480
rect 76148 5440 76149 5480
rect 76107 5431 76149 5440
rect 76491 5480 76533 5489
rect 76491 5440 76492 5480
rect 76532 5440 76533 5480
rect 76491 5431 76533 5440
rect 76875 5480 76917 5489
rect 76875 5440 76876 5480
rect 76916 5440 76917 5480
rect 76875 5431 76917 5440
rect 77451 5480 77493 5489
rect 77451 5440 77452 5480
rect 77492 5440 77493 5480
rect 77451 5431 77493 5440
rect 78027 5480 78069 5489
rect 78027 5440 78028 5480
rect 78068 5440 78069 5480
rect 78027 5431 78069 5440
rect 78699 5480 78741 5489
rect 78699 5440 78700 5480
rect 78740 5440 78741 5480
rect 78699 5431 78741 5440
rect 79851 5480 79893 5489
rect 79851 5440 79852 5480
rect 79892 5440 79893 5480
rect 79851 5431 79893 5440
rect 80043 5480 80085 5489
rect 80043 5440 80044 5480
rect 80084 5440 80085 5480
rect 80043 5431 80085 5440
rect 80619 5480 80661 5489
rect 80619 5440 80620 5480
rect 80660 5440 80661 5480
rect 80619 5431 80661 5440
rect 81099 5480 81141 5489
rect 81099 5440 81100 5480
rect 81140 5440 81141 5480
rect 81099 5431 81141 5440
rect 81483 5480 81525 5489
rect 81483 5440 81484 5480
rect 81524 5440 81525 5480
rect 81483 5431 81525 5440
rect 81867 5480 81909 5489
rect 81867 5440 81868 5480
rect 81908 5440 81909 5480
rect 81867 5431 81909 5440
rect 82347 5480 82389 5489
rect 82347 5440 82348 5480
rect 82388 5440 82389 5480
rect 82347 5431 82389 5440
rect 83115 5480 83157 5489
rect 83115 5440 83116 5480
rect 83156 5440 83157 5480
rect 83115 5431 83157 5440
rect 83499 5480 83541 5489
rect 83499 5440 83500 5480
rect 83540 5440 83541 5480
rect 83499 5431 83541 5440
rect 84555 5480 84597 5489
rect 84555 5440 84556 5480
rect 84596 5440 84597 5480
rect 84555 5431 84597 5440
rect 84843 5480 84885 5489
rect 84843 5440 84844 5480
rect 84884 5440 84885 5480
rect 84843 5431 84885 5440
rect 85227 5480 85269 5489
rect 85227 5440 85228 5480
rect 85268 5440 85269 5480
rect 85227 5431 85269 5440
rect 85611 5480 85653 5489
rect 85611 5440 85612 5480
rect 85652 5440 85653 5480
rect 85611 5431 85653 5440
rect 85995 5480 86037 5489
rect 85995 5440 85996 5480
rect 86036 5440 86037 5480
rect 85995 5431 86037 5440
rect 86379 5480 86421 5489
rect 86379 5440 86380 5480
rect 86420 5440 86421 5480
rect 86379 5431 86421 5440
rect 97707 5480 97749 5489
rect 97707 5440 97708 5480
rect 97748 5440 97749 5480
rect 97707 5431 97749 5440
rect 98091 5480 98133 5489
rect 98091 5440 98092 5480
rect 98132 5440 98133 5480
rect 98091 5431 98133 5440
rect 98283 5480 98325 5489
rect 98283 5440 98284 5480
rect 98324 5440 98325 5480
rect 98283 5431 98325 5440
rect 1152 5312 98784 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 64168 5312
rect 64208 5272 64250 5312
rect 64290 5272 64332 5312
rect 64372 5272 64414 5312
rect 64454 5272 64496 5312
rect 64536 5272 79288 5312
rect 79328 5272 79370 5312
rect 79410 5272 79452 5312
rect 79492 5272 79534 5312
rect 79574 5272 79616 5312
rect 79656 5272 94408 5312
rect 94448 5272 94490 5312
rect 94530 5272 94572 5312
rect 94612 5272 94654 5312
rect 94694 5272 94736 5312
rect 94776 5272 98784 5312
rect 1152 5248 98784 5272
rect 22827 5144 22869 5153
rect 22827 5104 22828 5144
rect 22868 5104 22869 5144
rect 22827 5095 22869 5104
rect 27819 5144 27861 5153
rect 27819 5104 27820 5144
rect 27860 5104 27861 5144
rect 27819 5095 27861 5104
rect 30507 5144 30549 5153
rect 30507 5104 30508 5144
rect 30548 5104 30549 5144
rect 30507 5095 30549 5104
rect 57867 5144 57909 5153
rect 57867 5104 57868 5144
rect 57908 5104 57909 5144
rect 57867 5095 57909 5104
rect 61803 5144 61845 5153
rect 61803 5104 61804 5144
rect 61844 5104 61845 5144
rect 61803 5095 61845 5104
rect 67563 5144 67605 5153
rect 67563 5104 67564 5144
rect 67604 5104 67605 5144
rect 67563 5095 67605 5104
rect 67947 5144 67989 5153
rect 67947 5104 67948 5144
rect 67988 5104 67989 5144
rect 67947 5095 67989 5104
rect 70539 5144 70581 5153
rect 70539 5104 70540 5144
rect 70580 5104 70581 5144
rect 70539 5095 70581 5104
rect 73323 5144 73365 5153
rect 73323 5104 73324 5144
rect 73364 5104 73365 5144
rect 73323 5095 73365 5104
rect 19947 5060 19989 5069
rect 19947 5020 19948 5060
rect 19988 5020 19989 5060
rect 19947 5011 19989 5020
rect 28395 5060 28437 5069
rect 28395 5020 28396 5060
rect 28436 5020 28437 5060
rect 28395 5011 28437 5020
rect 31179 5060 31221 5069
rect 31179 5020 31180 5060
rect 31220 5020 31221 5060
rect 31179 5011 31221 5020
rect 31659 5060 31701 5069
rect 31659 5020 31660 5060
rect 31700 5020 31701 5060
rect 31659 5011 31701 5020
rect 41547 5060 41589 5069
rect 41547 5020 41548 5060
rect 41588 5020 41589 5060
rect 41547 5011 41589 5020
rect 56715 5060 56757 5069
rect 56715 5020 56716 5060
rect 56756 5020 56757 5060
rect 56715 5011 56757 5020
rect 65451 5060 65493 5069
rect 65451 5020 65452 5060
rect 65492 5020 65493 5060
rect 65451 5011 65493 5020
rect 71691 5060 71733 5069
rect 71691 5020 71692 5060
rect 71732 5020 71733 5060
rect 71691 5011 71733 5020
rect 79467 5060 79509 5069
rect 79467 5020 79468 5060
rect 79508 5020 79509 5060
rect 79467 5011 79509 5020
rect 1699 4976 1757 4977
rect 1699 4936 1708 4976
rect 1748 4936 1757 4976
rect 1699 4935 1757 4936
rect 2083 4976 2141 4977
rect 2083 4936 2092 4976
rect 2132 4936 2141 4976
rect 2083 4935 2141 4936
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 2851 4976 2909 4977
rect 2851 4936 2860 4976
rect 2900 4936 2909 4976
rect 2851 4935 2909 4936
rect 13699 4976 13757 4977
rect 13699 4936 13708 4976
rect 13748 4936 13757 4976
rect 13699 4935 13757 4936
rect 13891 4976 13949 4977
rect 13891 4936 13900 4976
rect 13940 4936 13949 4976
rect 13891 4935 13949 4936
rect 14275 4976 14333 4977
rect 14275 4936 14284 4976
rect 14324 4936 14333 4976
rect 14275 4935 14333 4936
rect 14659 4976 14717 4977
rect 14659 4936 14668 4976
rect 14708 4936 14717 4976
rect 14659 4935 14717 4936
rect 15043 4976 15101 4977
rect 15043 4936 15052 4976
rect 15092 4936 15101 4976
rect 15043 4935 15101 4936
rect 15427 4976 15485 4977
rect 15427 4936 15436 4976
rect 15476 4936 15485 4976
rect 15427 4935 15485 4936
rect 16387 4976 16445 4977
rect 16387 4936 16396 4976
rect 16436 4936 16445 4976
rect 16387 4935 16445 4936
rect 16771 4976 16829 4977
rect 16771 4936 16780 4976
rect 16820 4936 16829 4976
rect 16771 4935 16829 4936
rect 20323 4976 20381 4977
rect 20323 4936 20332 4976
rect 20372 4936 20381 4976
rect 20323 4935 20381 4936
rect 21475 4976 21533 4977
rect 21475 4936 21484 4976
rect 21524 4936 21533 4976
rect 24651 4976 24693 4985
rect 21475 4935 21533 4936
rect 23779 4963 23837 4964
rect 23779 4923 23788 4963
rect 23828 4923 23837 4963
rect 24651 4936 24652 4976
rect 24692 4936 24693 4976
rect 24651 4927 24693 4936
rect 25891 4976 25949 4977
rect 25891 4936 25900 4976
rect 25940 4936 25949 4976
rect 25891 4935 25949 4936
rect 26083 4976 26141 4977
rect 26083 4936 26092 4976
rect 26132 4936 26141 4976
rect 26083 4935 26141 4936
rect 26467 4976 26525 4977
rect 26467 4936 26476 4976
rect 26516 4936 26525 4976
rect 26467 4935 26525 4936
rect 26851 4976 26909 4977
rect 26851 4936 26860 4976
rect 26900 4936 26909 4976
rect 26851 4935 26909 4936
rect 27235 4976 27293 4977
rect 27235 4936 27244 4976
rect 27284 4936 27293 4976
rect 27235 4935 27293 4936
rect 29155 4976 29213 4977
rect 29155 4936 29164 4976
rect 29204 4936 29213 4976
rect 29155 4935 29213 4936
rect 29539 4976 29597 4977
rect 29539 4936 29548 4976
rect 29588 4936 29597 4976
rect 29539 4935 29597 4936
rect 29923 4976 29981 4977
rect 29923 4936 29932 4976
rect 29972 4936 29981 4976
rect 29923 4935 29981 4936
rect 32227 4976 32285 4977
rect 32227 4936 32236 4976
rect 32276 4936 32285 4976
rect 32227 4935 32285 4936
rect 32611 4976 32669 4977
rect 32611 4936 32620 4976
rect 32660 4936 32669 4976
rect 32611 4935 32669 4936
rect 32995 4976 33053 4977
rect 32995 4936 33004 4976
rect 33044 4936 33053 4976
rect 32995 4935 33053 4936
rect 33379 4976 33437 4977
rect 33379 4936 33388 4976
rect 33428 4936 33437 4976
rect 33379 4935 33437 4936
rect 33763 4976 33821 4977
rect 33763 4936 33772 4976
rect 33812 4936 33821 4976
rect 33763 4935 33821 4936
rect 34147 4976 34205 4977
rect 34147 4936 34156 4976
rect 34196 4936 34205 4976
rect 34147 4935 34205 4936
rect 36651 4976 36693 4985
rect 36651 4936 36652 4976
rect 36692 4936 36693 4976
rect 36651 4927 36693 4936
rect 37123 4976 37181 4977
rect 37123 4936 37132 4976
rect 37172 4936 37181 4976
rect 37123 4935 37181 4936
rect 37507 4976 37565 4977
rect 37507 4936 37516 4976
rect 37556 4936 37565 4976
rect 37507 4935 37565 4936
rect 37891 4976 37949 4977
rect 37891 4936 37900 4976
rect 37940 4936 37949 4976
rect 37891 4935 37949 4936
rect 40195 4976 40253 4977
rect 40195 4936 40204 4976
rect 40244 4936 40253 4976
rect 40195 4935 40253 4936
rect 40579 4976 40637 4977
rect 40579 4936 40588 4976
rect 40628 4936 40637 4976
rect 40579 4935 40637 4936
rect 40963 4976 41021 4977
rect 40963 4936 40972 4976
rect 41012 4936 41021 4976
rect 40963 4935 41021 4936
rect 41347 4976 41405 4977
rect 41347 4936 41356 4976
rect 41396 4936 41405 4976
rect 41347 4935 41405 4936
rect 41731 4976 41789 4977
rect 41731 4936 41740 4976
rect 41780 4936 41789 4976
rect 41731 4935 41789 4936
rect 47971 4976 48029 4977
rect 47971 4936 47980 4976
rect 48020 4936 48029 4976
rect 47971 4935 48029 4936
rect 48355 4976 48413 4977
rect 48355 4936 48364 4976
rect 48404 4936 48413 4976
rect 48355 4935 48413 4936
rect 48739 4976 48797 4977
rect 48739 4936 48748 4976
rect 48788 4936 48797 4976
rect 48739 4935 48797 4936
rect 49123 4976 49181 4977
rect 49123 4936 49132 4976
rect 49172 4936 49181 4976
rect 49123 4935 49181 4936
rect 52387 4976 52445 4977
rect 52387 4936 52396 4976
rect 52436 4936 52445 4976
rect 52387 4935 52445 4936
rect 55747 4976 55805 4977
rect 55747 4936 55756 4976
rect 55796 4936 55805 4976
rect 55747 4935 55805 4936
rect 56427 4976 56469 4985
rect 56427 4936 56428 4976
rect 56468 4936 56469 4976
rect 46819 4934 46877 4935
rect 23779 4922 23837 4923
rect 17163 4905 17205 4914
rect 15819 4892 15861 4901
rect 15819 4852 15820 4892
rect 15860 4852 15861 4892
rect 15819 4843 15861 4852
rect 16011 4892 16053 4901
rect 16011 4852 16012 4892
rect 16052 4852 16053 4892
rect 17163 4865 17164 4905
rect 17204 4865 17205 4905
rect 20715 4905 20757 4914
rect 17163 4856 17205 4865
rect 17355 4892 17397 4901
rect 16011 4843 16053 4852
rect 17355 4852 17356 4892
rect 17396 4852 17397 4892
rect 17355 4843 17397 4852
rect 17547 4892 17589 4901
rect 17547 4852 17548 4892
rect 17588 4852 17589 4892
rect 18019 4892 18077 4893
rect 17547 4843 17589 4852
rect 17739 4881 17781 4890
rect 17739 4841 17740 4881
rect 17780 4841 17781 4881
rect 18019 4852 18028 4892
rect 18068 4852 18077 4892
rect 18019 4851 18077 4852
rect 18211 4892 18269 4893
rect 18211 4852 18220 4892
rect 18260 4852 18269 4892
rect 18211 4851 18269 4852
rect 18603 4892 18645 4901
rect 18603 4852 18604 4892
rect 18644 4852 18645 4892
rect 18603 4843 18645 4852
rect 18795 4892 18837 4901
rect 18795 4852 18796 4892
rect 18836 4852 18837 4892
rect 18795 4843 18837 4852
rect 18987 4892 19029 4901
rect 18987 4852 18988 4892
rect 19028 4852 19029 4892
rect 18987 4843 19029 4852
rect 19179 4892 19221 4901
rect 19179 4852 19180 4892
rect 19220 4852 19221 4892
rect 19179 4843 19221 4852
rect 19371 4892 19413 4901
rect 19371 4852 19372 4892
rect 19412 4852 19413 4892
rect 19371 4843 19413 4852
rect 19563 4892 19605 4901
rect 19563 4852 19564 4892
rect 19604 4852 19605 4892
rect 19563 4843 19605 4852
rect 19947 4892 19989 4901
rect 19947 4852 19948 4892
rect 19988 4852 19989 4892
rect 19947 4843 19989 4852
rect 20120 4892 20162 4901
rect 20120 4852 20121 4892
rect 20161 4852 20162 4892
rect 20715 4865 20716 4905
rect 20756 4865 20757 4905
rect 20715 4856 20757 4865
rect 20907 4892 20949 4901
rect 20120 4843 20162 4852
rect 20907 4852 20908 4892
rect 20948 4852 20949 4892
rect 20907 4843 20949 4852
rect 21099 4892 21141 4901
rect 21099 4852 21100 4892
rect 21140 4852 21141 4892
rect 21099 4843 21141 4852
rect 21291 4892 21333 4901
rect 21291 4852 21292 4892
rect 21332 4852 21333 4892
rect 21291 4843 21333 4852
rect 21867 4892 21909 4901
rect 21867 4852 21868 4892
rect 21908 4852 21909 4892
rect 21867 4843 21909 4852
rect 22059 4892 22101 4901
rect 22059 4852 22060 4892
rect 22100 4852 22101 4892
rect 22059 4843 22101 4852
rect 22251 4892 22293 4901
rect 22251 4852 22252 4892
rect 22292 4852 22293 4892
rect 22251 4843 22293 4852
rect 22443 4892 22485 4901
rect 22443 4852 22444 4892
rect 22484 4852 22485 4892
rect 22443 4843 22485 4852
rect 22627 4892 22685 4893
rect 22627 4852 22636 4892
rect 22676 4852 22685 4892
rect 22627 4851 22685 4852
rect 22827 4892 22869 4901
rect 22827 4852 22828 4892
rect 22868 4852 22869 4892
rect 22827 4843 22869 4852
rect 22915 4892 22973 4893
rect 22915 4852 22924 4892
rect 22964 4852 22973 4892
rect 22915 4851 22973 4852
rect 23403 4892 23445 4901
rect 23403 4852 23404 4892
rect 23444 4852 23445 4892
rect 23403 4843 23445 4852
rect 23595 4892 23637 4901
rect 23595 4852 23596 4892
rect 23636 4852 23637 4892
rect 23595 4843 23637 4852
rect 24171 4892 24213 4901
rect 24171 4852 24172 4892
rect 24212 4852 24213 4892
rect 24171 4843 24213 4852
rect 24363 4892 24405 4901
rect 24363 4852 24364 4892
rect 24404 4852 24405 4892
rect 24363 4843 24405 4852
rect 24555 4892 24597 4901
rect 24555 4852 24556 4892
rect 24596 4852 24597 4892
rect 24555 4843 24597 4852
rect 24747 4892 24789 4901
rect 24747 4852 24748 4892
rect 24788 4852 24789 4892
rect 24747 4843 24789 4852
rect 24939 4892 24981 4901
rect 24939 4852 24940 4892
rect 24980 4852 24981 4892
rect 24939 4843 24981 4852
rect 25131 4892 25173 4901
rect 25131 4852 25132 4892
rect 25172 4852 25173 4892
rect 25131 4843 25173 4852
rect 25323 4892 25365 4901
rect 25323 4852 25324 4892
rect 25364 4852 25365 4892
rect 25323 4843 25365 4852
rect 25515 4892 25557 4901
rect 25515 4852 25516 4892
rect 25556 4852 25557 4892
rect 25515 4843 25557 4852
rect 27627 4892 27669 4901
rect 27627 4852 27628 4892
rect 27668 4852 27669 4892
rect 27627 4843 27669 4852
rect 27819 4892 27861 4901
rect 27819 4852 27820 4892
rect 27860 4852 27861 4892
rect 27819 4843 27861 4852
rect 28011 4892 28053 4901
rect 28011 4852 28012 4892
rect 28052 4852 28053 4892
rect 28011 4843 28053 4852
rect 28203 4892 28245 4901
rect 28203 4852 28204 4892
rect 28244 4852 28245 4892
rect 28203 4843 28245 4852
rect 28395 4892 28437 4901
rect 28395 4852 28396 4892
rect 28436 4852 28437 4892
rect 28395 4843 28437 4852
rect 28587 4892 28629 4901
rect 28587 4852 28588 4892
rect 28628 4852 28629 4892
rect 28587 4843 28629 4852
rect 28779 4892 28821 4901
rect 28779 4852 28780 4892
rect 28820 4852 28821 4892
rect 28779 4843 28821 4852
rect 28971 4892 29013 4901
rect 28971 4852 28972 4892
rect 29012 4852 29013 4892
rect 28971 4843 29013 4852
rect 30315 4892 30357 4901
rect 30315 4852 30316 4892
rect 30356 4852 30357 4892
rect 30315 4843 30357 4852
rect 30507 4892 30549 4901
rect 30507 4852 30508 4892
rect 30548 4852 30549 4892
rect 30507 4843 30549 4852
rect 30699 4892 30741 4901
rect 30699 4852 30700 4892
rect 30740 4852 30741 4892
rect 30699 4843 30741 4852
rect 30891 4892 30933 4901
rect 30891 4852 30892 4892
rect 30932 4852 30933 4892
rect 30891 4843 30933 4852
rect 31171 4892 31229 4893
rect 31171 4852 31180 4892
rect 31220 4852 31229 4892
rect 31171 4851 31229 4852
rect 31363 4892 31421 4893
rect 31363 4852 31372 4892
rect 31412 4852 31421 4892
rect 31851 4892 31893 4901
rect 31363 4851 31421 4852
rect 31659 4881 31701 4890
rect 17739 4832 17781 4841
rect 31659 4841 31660 4881
rect 31700 4841 31701 4881
rect 31851 4852 31852 4892
rect 31892 4852 31893 4892
rect 31851 4843 31893 4852
rect 34539 4892 34581 4901
rect 34539 4852 34540 4892
rect 34580 4852 34581 4892
rect 34539 4843 34581 4852
rect 34731 4892 34773 4901
rect 34731 4852 34732 4892
rect 34772 4852 34773 4892
rect 34731 4843 34773 4852
rect 34923 4892 34965 4901
rect 34923 4852 34924 4892
rect 34964 4852 34965 4892
rect 34923 4843 34965 4852
rect 35115 4892 35157 4901
rect 35115 4852 35116 4892
rect 35156 4852 35157 4892
rect 35691 4892 35733 4901
rect 35115 4843 35157 4852
rect 35307 4881 35349 4890
rect 31659 4832 31701 4841
rect 35307 4841 35308 4881
rect 35348 4841 35349 4881
rect 35307 4832 35349 4841
rect 35499 4881 35541 4890
rect 35499 4841 35500 4881
rect 35540 4841 35541 4881
rect 35691 4852 35692 4892
rect 35732 4852 35733 4892
rect 35691 4843 35733 4852
rect 35883 4892 35925 4901
rect 35883 4852 35884 4892
rect 35924 4852 35925 4892
rect 35883 4843 35925 4852
rect 36067 4892 36125 4893
rect 36067 4852 36076 4892
rect 36116 4852 36125 4892
rect 36067 4851 36125 4852
rect 36259 4892 36317 4893
rect 36259 4852 36268 4892
rect 36308 4852 36317 4892
rect 36259 4851 36317 4852
rect 36555 4892 36597 4901
rect 36555 4852 36556 4892
rect 36596 4852 36597 4892
rect 36555 4843 36597 4852
rect 36747 4892 36789 4901
rect 36747 4852 36748 4892
rect 36788 4852 36789 4892
rect 36747 4843 36789 4852
rect 38283 4892 38325 4901
rect 38283 4852 38284 4892
rect 38324 4852 38325 4892
rect 38283 4843 38325 4852
rect 38475 4892 38517 4901
rect 38475 4852 38476 4892
rect 38516 4852 38517 4892
rect 38475 4843 38517 4852
rect 38667 4892 38709 4901
rect 38667 4852 38668 4892
rect 38708 4852 38709 4892
rect 38667 4843 38709 4852
rect 38859 4892 38901 4901
rect 38859 4852 38860 4892
rect 38900 4852 38901 4892
rect 38859 4843 38901 4852
rect 39043 4892 39101 4893
rect 39043 4852 39052 4892
rect 39092 4852 39101 4892
rect 39043 4851 39101 4852
rect 39235 4892 39293 4893
rect 39235 4852 39244 4892
rect 39284 4852 39293 4892
rect 39235 4851 39293 4852
rect 39627 4892 39669 4901
rect 39627 4852 39628 4892
rect 39668 4852 39669 4892
rect 39627 4843 39669 4852
rect 39819 4892 39861 4901
rect 39819 4852 39820 4892
rect 39860 4852 39861 4892
rect 39819 4843 39861 4852
rect 42987 4892 43029 4901
rect 42987 4852 42988 4892
rect 43028 4852 43029 4892
rect 42987 4843 43029 4852
rect 44323 4892 44381 4893
rect 44323 4852 44332 4892
rect 44372 4852 44381 4892
rect 44323 4851 44381 4852
rect 45571 4892 45629 4893
rect 45571 4852 45580 4892
rect 45620 4852 45629 4892
rect 45571 4851 45629 4852
rect 45859 4892 45917 4893
rect 45859 4852 45868 4892
rect 45908 4852 45917 4892
rect 45859 4851 45917 4852
rect 46059 4892 46101 4901
rect 46059 4852 46060 4892
rect 46100 4852 46101 4892
rect 46059 4843 46101 4852
rect 46147 4892 46205 4893
rect 46147 4852 46156 4892
rect 46196 4852 46205 4892
rect 46147 4851 46205 4852
rect 46531 4892 46589 4893
rect 46531 4852 46540 4892
rect 46580 4852 46589 4892
rect 46531 4851 46589 4852
rect 46635 4892 46677 4901
rect 46819 4894 46828 4934
rect 46868 4894 46877 4934
rect 56427 4927 56469 4936
rect 56899 4976 56957 4977
rect 56899 4936 56908 4976
rect 56948 4936 56957 4976
rect 56899 4935 56957 4936
rect 58819 4976 58877 4977
rect 58819 4936 58828 4976
rect 58868 4936 58877 4976
rect 58819 4935 58877 4936
rect 59203 4976 59261 4977
rect 59203 4936 59212 4976
rect 59252 4936 59261 4976
rect 59203 4935 59261 4936
rect 60355 4976 60413 4977
rect 60355 4936 60364 4976
rect 60404 4936 60413 4976
rect 60355 4935 60413 4936
rect 60739 4976 60797 4977
rect 60739 4936 60748 4976
rect 60788 4936 60797 4976
rect 60739 4935 60797 4936
rect 62755 4976 62813 4977
rect 62755 4936 62764 4976
rect 62804 4936 62813 4976
rect 62755 4935 62813 4936
rect 63907 4976 63965 4977
rect 63907 4936 63916 4976
rect 63956 4936 63965 4976
rect 63907 4935 63965 4936
rect 64291 4976 64349 4977
rect 64291 4936 64300 4976
rect 64340 4936 64349 4976
rect 64291 4935 64349 4936
rect 66115 4976 66173 4977
rect 66115 4936 66124 4976
rect 66164 4936 66173 4976
rect 66115 4935 66173 4936
rect 66499 4976 66557 4977
rect 66499 4936 66508 4976
rect 66548 4936 66557 4976
rect 66499 4935 66557 4936
rect 66883 4976 66941 4977
rect 66883 4936 66892 4976
rect 66932 4936 66941 4976
rect 66883 4935 66941 4936
rect 68899 4976 68957 4977
rect 68899 4936 68908 4976
rect 68948 4936 68957 4976
rect 68899 4935 68957 4936
rect 69283 4976 69341 4977
rect 69283 4936 69292 4976
rect 69332 4936 69341 4976
rect 69283 4935 69341 4936
rect 69675 4976 69717 4985
rect 69675 4936 69676 4976
rect 69716 4936 69717 4976
rect 69675 4927 69717 4936
rect 70915 4976 70973 4977
rect 70915 4936 70924 4976
rect 70964 4936 70973 4976
rect 70915 4935 70973 4936
rect 73699 4976 73757 4977
rect 73699 4936 73708 4976
rect 73748 4936 73757 4976
rect 73699 4935 73757 4936
rect 75915 4976 75957 4985
rect 75915 4936 75916 4976
rect 75956 4936 75957 4976
rect 75915 4927 75957 4936
rect 77539 4976 77597 4977
rect 77539 4936 77548 4976
rect 77588 4936 77597 4976
rect 77539 4935 77597 4936
rect 78499 4976 78557 4977
rect 78499 4936 78508 4976
rect 78548 4936 78557 4976
rect 78499 4935 78557 4936
rect 78883 4976 78941 4977
rect 78883 4936 78892 4976
rect 78932 4936 78941 4976
rect 78883 4935 78941 4936
rect 79843 4976 79901 4977
rect 79843 4936 79852 4976
rect 79892 4936 79901 4976
rect 79843 4935 79901 4936
rect 80227 4976 80285 4977
rect 80227 4936 80236 4976
rect 80276 4936 80285 4976
rect 80227 4935 80285 4936
rect 80611 4976 80669 4977
rect 80611 4936 80620 4976
rect 80660 4936 80669 4976
rect 80611 4935 80669 4936
rect 80907 4976 80949 4985
rect 80907 4936 80908 4976
rect 80948 4936 80949 4976
rect 80907 4927 80949 4936
rect 82147 4976 82205 4977
rect 82147 4936 82156 4976
rect 82196 4936 82205 4976
rect 82147 4935 82205 4936
rect 82531 4976 82589 4977
rect 82531 4936 82540 4976
rect 82580 4936 82589 4976
rect 82531 4935 82589 4936
rect 85795 4976 85853 4977
rect 85795 4936 85804 4976
rect 85844 4936 85853 4976
rect 85795 4935 85853 4936
rect 86179 4976 86237 4977
rect 86179 4936 86188 4976
rect 86228 4936 86237 4976
rect 86179 4935 86237 4936
rect 86563 4976 86621 4977
rect 86563 4936 86572 4976
rect 86612 4936 86621 4976
rect 86563 4935 86621 4936
rect 86947 4976 87005 4977
rect 86947 4936 86956 4976
rect 86996 4936 87005 4976
rect 86947 4935 87005 4936
rect 87331 4976 87389 4977
rect 87331 4936 87340 4976
rect 87380 4936 87389 4976
rect 87331 4935 87389 4936
rect 87715 4976 87773 4977
rect 87715 4936 87724 4976
rect 87764 4936 87773 4976
rect 87715 4935 87773 4936
rect 88099 4976 88157 4977
rect 88099 4936 88108 4976
rect 88148 4936 88157 4976
rect 88099 4935 88157 4936
rect 88483 4976 88541 4977
rect 88483 4936 88492 4976
rect 88532 4936 88541 4976
rect 88483 4935 88541 4936
rect 97123 4976 97181 4977
rect 97123 4936 97132 4976
rect 97172 4936 97181 4976
rect 97123 4935 97181 4936
rect 97699 4976 97757 4977
rect 97699 4936 97708 4976
rect 97748 4936 97757 4976
rect 97699 4935 97757 4936
rect 98083 4976 98141 4977
rect 98083 4936 98092 4976
rect 98132 4936 98141 4976
rect 98083 4935 98141 4936
rect 98467 4976 98525 4977
rect 98467 4936 98476 4976
rect 98516 4936 98525 4976
rect 98467 4935 98525 4936
rect 50864 4905 50906 4914
rect 46819 4893 46877 4894
rect 46635 4852 46636 4892
rect 46676 4852 46677 4892
rect 46635 4843 46677 4852
rect 47011 4892 47069 4893
rect 47011 4852 47020 4892
rect 47060 4852 47069 4892
rect 47011 4851 47069 4852
rect 47115 4892 47157 4901
rect 47115 4852 47116 4892
rect 47156 4852 47157 4892
rect 47115 4843 47157 4852
rect 47299 4892 47357 4893
rect 47299 4852 47308 4892
rect 47348 4852 47357 4892
rect 47299 4851 47357 4852
rect 47491 4892 47549 4893
rect 47491 4852 47500 4892
rect 47540 4852 47549 4892
rect 47491 4851 47549 4852
rect 47595 4892 47637 4901
rect 47595 4852 47596 4892
rect 47636 4852 47637 4892
rect 47595 4843 47637 4852
rect 47779 4892 47837 4893
rect 47779 4852 47788 4892
rect 47828 4852 47837 4892
rect 47779 4851 47837 4852
rect 49515 4892 49557 4901
rect 49515 4852 49516 4892
rect 49556 4852 49557 4892
rect 49515 4843 49557 4852
rect 49699 4892 49757 4893
rect 49699 4852 49708 4892
rect 49748 4852 49757 4892
rect 49699 4851 49757 4852
rect 49891 4892 49949 4893
rect 49891 4852 49900 4892
rect 49940 4852 49949 4892
rect 49891 4851 49949 4852
rect 50091 4892 50133 4901
rect 50091 4852 50092 4892
rect 50132 4852 50133 4892
rect 50091 4843 50133 4852
rect 50283 4892 50325 4901
rect 50283 4852 50284 4892
rect 50324 4852 50325 4892
rect 50283 4843 50325 4852
rect 50475 4892 50517 4901
rect 50475 4852 50476 4892
rect 50516 4852 50517 4892
rect 50475 4843 50517 4852
rect 50667 4892 50709 4901
rect 50667 4852 50668 4892
rect 50708 4852 50709 4892
rect 50864 4865 50865 4905
rect 50905 4865 50906 4905
rect 68139 4905 68181 4914
rect 50864 4856 50906 4865
rect 52771 4892 52829 4893
rect 50667 4843 50709 4852
rect 52771 4852 52780 4892
rect 52820 4852 52829 4892
rect 52771 4851 52829 4852
rect 54019 4892 54077 4893
rect 54019 4852 54028 4892
rect 54068 4852 54077 4892
rect 54019 4851 54077 4852
rect 54979 4892 55037 4893
rect 54979 4852 54988 4892
rect 55028 4852 55037 4892
rect 54979 4851 55037 4852
rect 55179 4892 55221 4901
rect 55179 4852 55180 4892
rect 55220 4852 55221 4892
rect 55179 4843 55221 4852
rect 55371 4892 55413 4901
rect 55371 4852 55372 4892
rect 55412 4852 55413 4892
rect 55371 4843 55413 4852
rect 55947 4892 55989 4901
rect 55947 4852 55948 4892
rect 55988 4852 55989 4892
rect 55947 4843 55989 4852
rect 56131 4892 56189 4893
rect 56131 4852 56140 4892
rect 56180 4852 56189 4892
rect 56131 4851 56189 4852
rect 56331 4892 56373 4901
rect 56331 4852 56332 4892
rect 56372 4852 56373 4892
rect 57099 4892 57141 4901
rect 56331 4843 56373 4852
rect 56515 4871 56573 4872
rect 35499 4832 35541 4841
rect 56515 4831 56524 4871
rect 56564 4831 56573 4871
rect 57099 4852 57100 4892
rect 57140 4852 57141 4892
rect 57099 4843 57141 4852
rect 57291 4892 57333 4901
rect 57291 4852 57292 4892
rect 57332 4852 57333 4892
rect 57291 4843 57333 4852
rect 57483 4892 57525 4901
rect 57483 4852 57484 4892
rect 57524 4852 57525 4892
rect 57483 4843 57525 4852
rect 57675 4892 57717 4901
rect 57675 4852 57676 4892
rect 57716 4852 57717 4892
rect 57675 4843 57717 4852
rect 57867 4892 57909 4901
rect 57867 4852 57868 4892
rect 57908 4852 57909 4892
rect 57867 4843 57909 4852
rect 58059 4892 58101 4901
rect 58059 4852 58060 4892
rect 58100 4852 58101 4892
rect 58059 4843 58101 4852
rect 58251 4892 58293 4901
rect 58251 4852 58252 4892
rect 58292 4852 58293 4892
rect 58251 4843 58293 4852
rect 58443 4892 58485 4901
rect 58443 4852 58444 4892
rect 58484 4852 58485 4892
rect 58443 4843 58485 4852
rect 59683 4892 59741 4893
rect 59683 4852 59692 4892
rect 59732 4852 59741 4892
rect 59683 4851 59741 4852
rect 59875 4892 59933 4893
rect 59875 4852 59884 4892
rect 59924 4852 59933 4892
rect 59875 4851 59933 4852
rect 61315 4892 61373 4893
rect 61315 4852 61324 4892
rect 61364 4852 61373 4892
rect 61315 4851 61373 4852
rect 61707 4892 61749 4901
rect 61707 4852 61708 4892
rect 61748 4852 61749 4892
rect 62083 4892 62141 4893
rect 61707 4843 61749 4852
rect 61891 4871 61949 4872
rect 56515 4830 56573 4831
rect 61891 4831 61900 4871
rect 61940 4831 61949 4871
rect 62083 4852 62092 4892
rect 62132 4852 62141 4892
rect 62083 4851 62141 4852
rect 62275 4892 62333 4893
rect 62275 4852 62284 4892
rect 62324 4852 62333 4892
rect 62275 4851 62333 4852
rect 63235 4892 63293 4893
rect 63235 4852 63244 4892
rect 63284 4852 63293 4892
rect 63235 4851 63293 4852
rect 63427 4892 63485 4893
rect 63427 4852 63436 4892
rect 63476 4852 63485 4892
rect 63427 4851 63485 4852
rect 64771 4892 64829 4893
rect 64771 4852 64780 4892
rect 64820 4852 64829 4892
rect 64771 4851 64829 4852
rect 67179 4892 67221 4901
rect 67179 4852 67180 4892
rect 67220 4852 67221 4892
rect 67179 4843 67221 4852
rect 67371 4892 67413 4901
rect 67371 4852 67372 4892
rect 67412 4852 67413 4892
rect 67371 4843 67413 4852
rect 67563 4892 67605 4901
rect 67563 4852 67564 4892
rect 67604 4852 67605 4892
rect 67563 4843 67605 4852
rect 67755 4892 67797 4901
rect 67755 4852 67756 4892
rect 67796 4852 67797 4892
rect 67755 4843 67797 4852
rect 67947 4892 67989 4901
rect 67947 4852 67948 4892
rect 67988 4852 67989 4892
rect 68139 4865 68140 4905
rect 68180 4865 68181 4905
rect 73126 4905 73168 4914
rect 68139 4856 68181 4865
rect 68331 4892 68373 4901
rect 67947 4843 67989 4852
rect 68331 4852 68332 4892
rect 68372 4852 68373 4892
rect 68331 4843 68373 4852
rect 68523 4892 68565 4901
rect 68523 4852 68524 4892
rect 68564 4852 68565 4892
rect 68523 4843 68565 4852
rect 69579 4892 69621 4901
rect 69579 4852 69580 4892
rect 69620 4852 69621 4892
rect 69579 4843 69621 4852
rect 69771 4892 69813 4901
rect 69771 4852 69772 4892
rect 69812 4852 69813 4892
rect 69771 4843 69813 4852
rect 69963 4892 70005 4901
rect 69963 4852 69964 4892
rect 70004 4852 70005 4892
rect 69963 4843 70005 4852
rect 70155 4892 70197 4901
rect 70155 4852 70156 4892
rect 70196 4852 70197 4892
rect 70155 4843 70197 4852
rect 70347 4892 70389 4901
rect 70347 4852 70348 4892
rect 70388 4852 70389 4892
rect 70347 4843 70389 4852
rect 70539 4892 70581 4901
rect 70539 4852 70540 4892
rect 70580 4852 70581 4892
rect 70539 4843 70581 4852
rect 71115 4892 71157 4901
rect 71115 4852 71116 4892
rect 71156 4852 71157 4892
rect 71115 4843 71157 4852
rect 71307 4892 71349 4901
rect 71307 4852 71308 4892
rect 71348 4852 71349 4892
rect 71307 4843 71349 4852
rect 71499 4892 71541 4901
rect 71499 4852 71500 4892
rect 71540 4852 71541 4892
rect 71499 4843 71541 4852
rect 71691 4892 71733 4901
rect 71691 4852 71692 4892
rect 71732 4852 71733 4892
rect 71691 4843 71733 4852
rect 71979 4892 72021 4901
rect 71979 4852 71980 4892
rect 72020 4852 72021 4892
rect 71979 4843 72021 4852
rect 72171 4892 72213 4901
rect 72171 4852 72172 4892
rect 72212 4852 72213 4892
rect 72171 4843 72213 4852
rect 72363 4892 72405 4901
rect 72363 4852 72364 4892
rect 72404 4852 72405 4892
rect 72363 4843 72405 4852
rect 72555 4892 72597 4901
rect 72555 4852 72556 4892
rect 72596 4852 72597 4892
rect 72939 4892 72981 4901
rect 72555 4843 72597 4852
rect 72742 4881 72800 4882
rect 72742 4841 72751 4881
rect 72791 4841 72800 4881
rect 72939 4852 72940 4892
rect 72980 4852 72981 4892
rect 73126 4865 73127 4905
rect 73167 4865 73168 4905
rect 81387 4905 81429 4914
rect 73126 4856 73168 4865
rect 73323 4892 73365 4901
rect 72939 4843 72981 4852
rect 73323 4852 73324 4892
rect 73364 4852 73365 4892
rect 73323 4843 73365 4852
rect 74187 4892 74229 4901
rect 74187 4852 74188 4892
rect 74228 4852 74229 4892
rect 74187 4843 74229 4852
rect 74379 4892 74421 4901
rect 74379 4852 74380 4892
rect 74420 4852 74421 4892
rect 74379 4843 74421 4852
rect 74659 4892 74717 4893
rect 74659 4852 74668 4892
rect 74708 4852 74717 4892
rect 74659 4851 74717 4852
rect 75819 4892 75861 4901
rect 75819 4852 75820 4892
rect 75860 4852 75861 4892
rect 75819 4843 75861 4852
rect 76011 4892 76053 4901
rect 76011 4852 76012 4892
rect 76052 4852 76053 4892
rect 76395 4892 76437 4901
rect 76011 4843 76053 4852
rect 76198 4881 76256 4882
rect 72742 4840 72800 4841
rect 76198 4841 76207 4881
rect 76247 4841 76256 4881
rect 76395 4852 76396 4892
rect 76436 4852 76437 4892
rect 76395 4843 76437 4852
rect 76587 4892 76629 4901
rect 76587 4852 76588 4892
rect 76628 4852 76629 4892
rect 76587 4843 76629 4852
rect 76779 4892 76821 4901
rect 76779 4852 76780 4892
rect 76820 4852 76821 4892
rect 76779 4843 76821 4852
rect 76971 4892 77013 4901
rect 76971 4852 76972 4892
rect 77012 4852 77013 4892
rect 76971 4843 77013 4852
rect 77163 4892 77205 4901
rect 77163 4852 77164 4892
rect 77204 4852 77205 4892
rect 77163 4843 77205 4852
rect 77827 4892 77885 4893
rect 77827 4852 77836 4892
rect 77876 4852 77885 4892
rect 77827 4851 77885 4852
rect 78019 4892 78077 4893
rect 78019 4852 78028 4892
rect 78068 4852 78077 4892
rect 78019 4851 78077 4852
rect 79275 4892 79317 4901
rect 79275 4852 79276 4892
rect 79316 4852 79317 4892
rect 79275 4843 79317 4852
rect 79467 4892 79509 4901
rect 79467 4852 79468 4892
rect 79508 4852 79509 4892
rect 79467 4843 79509 4852
rect 80811 4892 80853 4901
rect 80811 4852 80812 4892
rect 80852 4852 80853 4892
rect 80811 4843 80853 4852
rect 81003 4892 81045 4901
rect 81003 4852 81004 4892
rect 81044 4852 81045 4892
rect 81003 4843 81045 4852
rect 81195 4892 81237 4901
rect 81195 4852 81196 4892
rect 81236 4852 81237 4892
rect 81387 4865 81388 4905
rect 81428 4865 81429 4905
rect 81387 4856 81429 4865
rect 81579 4892 81621 4901
rect 81195 4843 81237 4852
rect 81579 4852 81580 4892
rect 81620 4852 81621 4892
rect 81579 4843 81621 4852
rect 81771 4892 81813 4901
rect 81771 4852 81772 4892
rect 81812 4852 81813 4892
rect 81771 4843 81813 4852
rect 82731 4892 82773 4901
rect 82731 4852 82732 4892
rect 82772 4852 82773 4892
rect 82731 4843 82773 4852
rect 82923 4892 82965 4901
rect 82923 4852 82924 4892
rect 82964 4852 82965 4892
rect 82923 4843 82965 4852
rect 83307 4892 83349 4901
rect 83307 4852 83308 4892
rect 83348 4852 83349 4892
rect 83307 4843 83349 4852
rect 83499 4892 83541 4901
rect 83499 4852 83500 4892
rect 83540 4852 83541 4892
rect 83499 4843 83541 4852
rect 83691 4892 83733 4901
rect 83691 4852 83692 4892
rect 83732 4852 83733 4892
rect 83691 4843 83733 4852
rect 83883 4892 83925 4901
rect 83883 4852 83884 4892
rect 83924 4852 83925 4892
rect 83883 4843 83925 4852
rect 84555 4892 84597 4901
rect 84555 4852 84556 4892
rect 84596 4852 84597 4892
rect 84555 4843 84597 4852
rect 76198 4840 76256 4841
rect 61891 4830 61949 4831
rect 19083 4808 19125 4817
rect 19083 4768 19084 4808
rect 19124 4768 19125 4808
rect 19083 4759 19125 4768
rect 20811 4808 20853 4817
rect 20811 4768 20812 4808
rect 20852 4768 20853 4808
rect 20811 4759 20853 4768
rect 35403 4808 35445 4817
rect 35403 4768 35404 4808
rect 35444 4768 35445 4808
rect 35403 4759 35445 4768
rect 42211 4808 42269 4809
rect 42211 4768 42220 4808
rect 42260 4768 42269 4808
rect 42211 4767 42269 4768
rect 43459 4808 43517 4809
rect 43459 4768 43468 4808
rect 43508 4768 43517 4808
rect 43459 4767 43517 4768
rect 44707 4808 44765 4809
rect 44707 4768 44716 4808
rect 44756 4768 44765 4808
rect 44707 4767 44765 4768
rect 49611 4808 49653 4817
rect 49611 4768 49612 4808
rect 49652 4768 49653 4808
rect 49611 4759 49653 4768
rect 49995 4808 50037 4817
rect 49995 4768 49996 4808
rect 50036 4768 50037 4808
rect 49995 4759 50037 4768
rect 53635 4808 53693 4809
rect 53635 4768 53644 4808
rect 53684 4768 53693 4808
rect 53635 4767 53693 4768
rect 56043 4808 56085 4817
rect 56043 4768 56044 4808
rect 56084 4768 56085 4808
rect 56043 4759 56085 4768
rect 72075 4808 72117 4817
rect 72075 4768 72076 4808
rect 72116 4768 72117 4808
rect 72075 4759 72117 4768
rect 1515 4724 1557 4733
rect 1515 4684 1516 4724
rect 1556 4684 1557 4724
rect 1515 4675 1557 4684
rect 1899 4724 1941 4733
rect 1899 4684 1900 4724
rect 1940 4684 1941 4724
rect 1899 4675 1941 4684
rect 2283 4724 2325 4733
rect 2283 4684 2284 4724
rect 2324 4684 2325 4724
rect 2283 4675 2325 4684
rect 2667 4724 2709 4733
rect 2667 4684 2668 4724
rect 2708 4684 2709 4724
rect 2667 4675 2709 4684
rect 13515 4724 13557 4733
rect 13515 4684 13516 4724
rect 13556 4684 13557 4724
rect 13515 4675 13557 4684
rect 14091 4724 14133 4733
rect 14091 4684 14092 4724
rect 14132 4684 14133 4724
rect 14091 4675 14133 4684
rect 14475 4724 14517 4733
rect 14475 4684 14476 4724
rect 14516 4684 14517 4724
rect 14475 4675 14517 4684
rect 14859 4724 14901 4733
rect 14859 4684 14860 4724
rect 14900 4684 14901 4724
rect 14859 4675 14901 4684
rect 15243 4724 15285 4733
rect 15243 4684 15244 4724
rect 15284 4684 15285 4724
rect 15243 4675 15285 4684
rect 15627 4724 15669 4733
rect 15627 4684 15628 4724
rect 15668 4684 15669 4724
rect 15627 4675 15669 4684
rect 15915 4724 15957 4733
rect 15915 4684 15916 4724
rect 15956 4684 15957 4724
rect 15915 4675 15957 4684
rect 16587 4724 16629 4733
rect 16587 4684 16588 4724
rect 16628 4684 16629 4724
rect 16587 4675 16629 4684
rect 16971 4724 17013 4733
rect 16971 4684 16972 4724
rect 17012 4684 17013 4724
rect 16971 4675 17013 4684
rect 17259 4724 17301 4733
rect 17259 4684 17260 4724
rect 17300 4684 17301 4724
rect 17259 4675 17301 4684
rect 17643 4724 17685 4733
rect 17643 4684 17644 4724
rect 17684 4684 17685 4724
rect 17643 4675 17685 4684
rect 18699 4724 18741 4733
rect 18699 4684 18700 4724
rect 18740 4684 18741 4724
rect 18699 4675 18741 4684
rect 19467 4724 19509 4733
rect 19467 4684 19468 4724
rect 19508 4684 19509 4724
rect 19467 4675 19509 4684
rect 20523 4724 20565 4733
rect 20523 4684 20524 4724
rect 20564 4684 20565 4724
rect 20523 4675 20565 4684
rect 21195 4724 21237 4733
rect 21195 4684 21196 4724
rect 21236 4684 21237 4724
rect 21195 4675 21237 4684
rect 21675 4724 21717 4733
rect 21675 4684 21676 4724
rect 21716 4684 21717 4724
rect 21675 4675 21717 4684
rect 21963 4724 22005 4733
rect 21963 4684 21964 4724
rect 22004 4684 22005 4724
rect 21963 4675 22005 4684
rect 22347 4724 22389 4733
rect 22347 4684 22348 4724
rect 22388 4684 22389 4724
rect 22347 4675 22389 4684
rect 23499 4724 23541 4733
rect 23499 4684 23500 4724
rect 23540 4684 23541 4724
rect 23499 4675 23541 4684
rect 23979 4724 24021 4733
rect 23979 4684 23980 4724
rect 24020 4684 24021 4724
rect 23979 4675 24021 4684
rect 24267 4724 24309 4733
rect 24267 4684 24268 4724
rect 24308 4684 24309 4724
rect 24267 4675 24309 4684
rect 25035 4724 25077 4733
rect 25035 4684 25036 4724
rect 25076 4684 25077 4724
rect 25035 4675 25077 4684
rect 25419 4724 25461 4733
rect 25419 4684 25420 4724
rect 25460 4684 25461 4724
rect 25419 4675 25461 4684
rect 25707 4724 25749 4733
rect 25707 4684 25708 4724
rect 25748 4684 25749 4724
rect 25707 4675 25749 4684
rect 26283 4724 26325 4733
rect 26283 4684 26284 4724
rect 26324 4684 26325 4724
rect 26283 4675 26325 4684
rect 26667 4724 26709 4733
rect 26667 4684 26668 4724
rect 26708 4684 26709 4724
rect 26667 4675 26709 4684
rect 27051 4724 27093 4733
rect 27051 4684 27052 4724
rect 27092 4684 27093 4724
rect 27051 4675 27093 4684
rect 27435 4724 27477 4733
rect 27435 4684 27436 4724
rect 27476 4684 27477 4724
rect 27435 4675 27477 4684
rect 28107 4724 28149 4733
rect 28107 4684 28108 4724
rect 28148 4684 28149 4724
rect 28107 4675 28149 4684
rect 28875 4724 28917 4733
rect 28875 4684 28876 4724
rect 28916 4684 28917 4724
rect 28875 4675 28917 4684
rect 29355 4724 29397 4733
rect 29355 4684 29356 4724
rect 29396 4684 29397 4724
rect 29355 4675 29397 4684
rect 29739 4724 29781 4733
rect 29739 4684 29740 4724
rect 29780 4684 29781 4724
rect 29739 4675 29781 4684
rect 30123 4724 30165 4733
rect 30123 4684 30124 4724
rect 30164 4684 30165 4724
rect 30123 4675 30165 4684
rect 30795 4724 30837 4733
rect 30795 4684 30796 4724
rect 30836 4684 30837 4724
rect 30795 4675 30837 4684
rect 32427 4724 32469 4733
rect 32427 4684 32428 4724
rect 32468 4684 32469 4724
rect 32427 4675 32469 4684
rect 32811 4724 32853 4733
rect 32811 4684 32812 4724
rect 32852 4684 32853 4724
rect 32811 4675 32853 4684
rect 33195 4724 33237 4733
rect 33195 4684 33196 4724
rect 33236 4684 33237 4724
rect 33195 4675 33237 4684
rect 33579 4724 33621 4733
rect 33579 4684 33580 4724
rect 33620 4684 33621 4724
rect 33579 4675 33621 4684
rect 33963 4724 34005 4733
rect 33963 4684 33964 4724
rect 34004 4684 34005 4724
rect 33963 4675 34005 4684
rect 34347 4724 34389 4733
rect 34347 4684 34348 4724
rect 34388 4684 34389 4724
rect 34347 4675 34389 4684
rect 34635 4724 34677 4733
rect 34635 4684 34636 4724
rect 34676 4684 34677 4724
rect 34635 4675 34677 4684
rect 35019 4724 35061 4733
rect 35019 4684 35020 4724
rect 35060 4684 35061 4724
rect 35019 4675 35061 4684
rect 35787 4724 35829 4733
rect 35787 4684 35788 4724
rect 35828 4684 35829 4724
rect 35787 4675 35829 4684
rect 37323 4724 37365 4733
rect 37323 4684 37324 4724
rect 37364 4684 37365 4724
rect 37323 4675 37365 4684
rect 37707 4724 37749 4733
rect 37707 4684 37708 4724
rect 37748 4684 37749 4724
rect 37707 4675 37749 4684
rect 38091 4724 38133 4733
rect 38091 4684 38092 4724
rect 38132 4684 38133 4724
rect 38091 4675 38133 4684
rect 38379 4724 38421 4733
rect 38379 4684 38380 4724
rect 38420 4684 38421 4724
rect 38379 4675 38421 4684
rect 38763 4724 38805 4733
rect 38763 4684 38764 4724
rect 38804 4684 38805 4724
rect 38763 4675 38805 4684
rect 39723 4724 39765 4733
rect 39723 4684 39724 4724
rect 39764 4684 39765 4724
rect 39723 4675 39765 4684
rect 40395 4724 40437 4733
rect 40395 4684 40396 4724
rect 40436 4684 40437 4724
rect 40395 4675 40437 4684
rect 40779 4724 40821 4733
rect 40779 4684 40780 4724
rect 40820 4684 40821 4724
rect 40779 4675 40821 4684
rect 41163 4724 41205 4733
rect 41163 4684 41164 4724
rect 41204 4684 41205 4724
rect 41163 4675 41205 4684
rect 41931 4724 41973 4733
rect 41931 4684 41932 4724
rect 41972 4684 41973 4724
rect 41931 4675 41973 4684
rect 45867 4724 45909 4733
rect 45867 4684 45868 4724
rect 45908 4684 45909 4724
rect 45867 4675 45909 4684
rect 46827 4724 46869 4733
rect 46827 4684 46828 4724
rect 46868 4684 46869 4724
rect 46827 4675 46869 4684
rect 47307 4724 47349 4733
rect 47307 4684 47308 4724
rect 47348 4684 47349 4724
rect 47307 4675 47349 4684
rect 47787 4724 47829 4733
rect 47787 4684 47788 4724
rect 47828 4684 47829 4724
rect 47787 4675 47829 4684
rect 48171 4724 48213 4733
rect 48171 4684 48172 4724
rect 48212 4684 48213 4724
rect 48171 4675 48213 4684
rect 48555 4724 48597 4733
rect 48555 4684 48556 4724
rect 48596 4684 48597 4724
rect 48555 4675 48597 4684
rect 48939 4724 48981 4733
rect 48939 4684 48940 4724
rect 48980 4684 48981 4724
rect 48939 4675 48981 4684
rect 49323 4724 49365 4733
rect 49323 4684 49324 4724
rect 49364 4684 49365 4724
rect 49323 4675 49365 4684
rect 50379 4724 50421 4733
rect 50379 4684 50380 4724
rect 50420 4684 50421 4724
rect 50379 4675 50421 4684
rect 50763 4724 50805 4733
rect 50763 4684 50764 4724
rect 50804 4684 50805 4724
rect 50763 4675 50805 4684
rect 52203 4724 52245 4733
rect 52203 4684 52204 4724
rect 52244 4684 52245 4724
rect 52203 4675 52245 4684
rect 55275 4724 55317 4733
rect 55275 4684 55276 4724
rect 55316 4684 55317 4724
rect 55275 4675 55317 4684
rect 55563 4724 55605 4733
rect 55563 4684 55564 4724
rect 55604 4684 55605 4724
rect 55563 4675 55605 4684
rect 57195 4724 57237 4733
rect 57195 4684 57196 4724
rect 57236 4684 57237 4724
rect 57195 4675 57237 4684
rect 57579 4724 57621 4733
rect 57579 4684 57580 4724
rect 57620 4684 57621 4724
rect 57579 4675 57621 4684
rect 58347 4724 58389 4733
rect 58347 4684 58348 4724
rect 58388 4684 58389 4724
rect 58347 4675 58389 4684
rect 58635 4724 58677 4733
rect 58635 4684 58636 4724
rect 58676 4684 58677 4724
rect 58635 4675 58677 4684
rect 59019 4724 59061 4733
rect 59019 4684 59020 4724
rect 59060 4684 59061 4724
rect 59019 4675 59061 4684
rect 59691 4724 59733 4733
rect 59691 4684 59692 4724
rect 59732 4684 59733 4724
rect 59691 4675 59733 4684
rect 60171 4724 60213 4733
rect 60171 4684 60172 4724
rect 60212 4684 60213 4724
rect 60171 4675 60213 4684
rect 60555 4724 60597 4733
rect 60555 4684 60556 4724
rect 60596 4684 60597 4724
rect 60555 4675 60597 4684
rect 61219 4724 61277 4725
rect 61219 4684 61228 4724
rect 61268 4684 61277 4724
rect 61219 4683 61277 4684
rect 61507 4724 61565 4725
rect 61507 4684 61516 4724
rect 61556 4684 61565 4724
rect 61507 4683 61565 4684
rect 62571 4724 62613 4733
rect 62571 4684 62572 4724
rect 62612 4684 62613 4724
rect 62571 4675 62613 4684
rect 63723 4724 63765 4733
rect 63723 4684 63724 4724
rect 63764 4684 63765 4724
rect 63723 4675 63765 4684
rect 64107 4724 64149 4733
rect 64107 4684 64108 4724
rect 64148 4684 64149 4724
rect 64107 4675 64149 4684
rect 65931 4724 65973 4733
rect 65931 4684 65932 4724
rect 65972 4684 65973 4724
rect 65931 4675 65973 4684
rect 66315 4724 66357 4733
rect 66315 4684 66316 4724
rect 66356 4684 66357 4724
rect 66315 4675 66357 4684
rect 66699 4724 66741 4733
rect 66699 4684 66700 4724
rect 66740 4684 66741 4724
rect 66699 4675 66741 4684
rect 67275 4724 67317 4733
rect 67275 4684 67276 4724
rect 67316 4684 67317 4724
rect 67275 4675 67317 4684
rect 68427 4724 68469 4733
rect 68427 4684 68428 4724
rect 68468 4684 68469 4724
rect 68427 4675 68469 4684
rect 68715 4724 68757 4733
rect 68715 4684 68716 4724
rect 68756 4684 68757 4724
rect 68715 4675 68757 4684
rect 69099 4724 69141 4733
rect 69099 4684 69100 4724
rect 69140 4684 69141 4724
rect 69099 4675 69141 4684
rect 70059 4724 70101 4733
rect 70059 4684 70060 4724
rect 70100 4684 70101 4724
rect 70059 4675 70101 4684
rect 70731 4724 70773 4733
rect 70731 4684 70732 4724
rect 70772 4684 70773 4724
rect 70731 4675 70773 4684
rect 71211 4724 71253 4733
rect 71211 4684 71212 4724
rect 71252 4684 71253 4724
rect 71211 4675 71253 4684
rect 72459 4724 72501 4733
rect 72459 4684 72460 4724
rect 72500 4684 72501 4724
rect 72459 4675 72501 4684
rect 72843 4724 72885 4733
rect 72843 4684 72844 4724
rect 72884 4684 72885 4724
rect 72843 4675 72885 4684
rect 73515 4724 73557 4733
rect 73515 4684 73516 4724
rect 73556 4684 73557 4724
rect 73515 4675 73557 4684
rect 74283 4724 74325 4733
rect 74283 4684 74284 4724
rect 74324 4684 74325 4724
rect 74283 4675 74325 4684
rect 75147 4724 75189 4733
rect 75147 4684 75148 4724
rect 75188 4684 75189 4724
rect 75147 4675 75189 4684
rect 76299 4724 76341 4733
rect 76299 4684 76300 4724
rect 76340 4684 76341 4724
rect 76299 4675 76341 4684
rect 76683 4724 76725 4733
rect 76683 4684 76684 4724
rect 76724 4684 76725 4724
rect 76683 4675 76725 4684
rect 77067 4724 77109 4733
rect 77067 4684 77068 4724
rect 77108 4684 77109 4724
rect 77067 4675 77109 4684
rect 77355 4724 77397 4733
rect 77355 4684 77356 4724
rect 77396 4684 77397 4724
rect 77355 4675 77397 4684
rect 78315 4724 78357 4733
rect 78315 4684 78316 4724
rect 78356 4684 78357 4724
rect 78315 4675 78357 4684
rect 78699 4724 78741 4733
rect 78699 4684 78700 4724
rect 78740 4684 78741 4724
rect 78699 4675 78741 4684
rect 79659 4724 79701 4733
rect 79659 4684 79660 4724
rect 79700 4684 79701 4724
rect 79659 4675 79701 4684
rect 80043 4724 80085 4733
rect 80043 4684 80044 4724
rect 80084 4684 80085 4724
rect 80043 4675 80085 4684
rect 80427 4724 80469 4733
rect 80427 4684 80428 4724
rect 80468 4684 80469 4724
rect 80427 4675 80469 4684
rect 81291 4724 81333 4733
rect 81291 4684 81292 4724
rect 81332 4684 81333 4724
rect 81291 4675 81333 4684
rect 81675 4724 81717 4733
rect 81675 4684 81676 4724
rect 81716 4684 81717 4724
rect 81675 4675 81717 4684
rect 81963 4724 82005 4733
rect 81963 4684 81964 4724
rect 82004 4684 82005 4724
rect 81963 4675 82005 4684
rect 82347 4724 82389 4733
rect 82347 4684 82348 4724
rect 82388 4684 82389 4724
rect 82347 4675 82389 4684
rect 82827 4724 82869 4733
rect 82827 4684 82828 4724
rect 82868 4684 82869 4724
rect 82827 4675 82869 4684
rect 83403 4724 83445 4733
rect 83403 4684 83404 4724
rect 83444 4684 83445 4724
rect 83403 4675 83445 4684
rect 83787 4724 83829 4733
rect 83787 4684 83788 4724
rect 83828 4684 83829 4724
rect 83787 4675 83829 4684
rect 84939 4724 84981 4733
rect 84939 4684 84940 4724
rect 84980 4684 84981 4724
rect 84939 4675 84981 4684
rect 85611 4724 85653 4733
rect 85611 4684 85612 4724
rect 85652 4684 85653 4724
rect 85611 4675 85653 4684
rect 85995 4724 86037 4733
rect 85995 4684 85996 4724
rect 86036 4684 86037 4724
rect 85995 4675 86037 4684
rect 86379 4724 86421 4733
rect 86379 4684 86380 4724
rect 86420 4684 86421 4724
rect 86379 4675 86421 4684
rect 86763 4724 86805 4733
rect 86763 4684 86764 4724
rect 86804 4684 86805 4724
rect 86763 4675 86805 4684
rect 87147 4724 87189 4733
rect 87147 4684 87148 4724
rect 87188 4684 87189 4724
rect 87147 4675 87189 4684
rect 87531 4724 87573 4733
rect 87531 4684 87532 4724
rect 87572 4684 87573 4724
rect 87531 4675 87573 4684
rect 87915 4724 87957 4733
rect 87915 4684 87916 4724
rect 87956 4684 87957 4724
rect 87915 4675 87957 4684
rect 88299 4724 88341 4733
rect 88299 4684 88300 4724
rect 88340 4684 88341 4724
rect 88299 4675 88341 4684
rect 97323 4724 97365 4733
rect 97323 4684 97324 4724
rect 97364 4684 97365 4724
rect 97323 4675 97365 4684
rect 97515 4724 97557 4733
rect 97515 4684 97516 4724
rect 97556 4684 97557 4724
rect 97515 4675 97557 4684
rect 97899 4724 97941 4733
rect 97899 4684 97900 4724
rect 97940 4684 97941 4724
rect 97899 4675 97941 4684
rect 98283 4724 98325 4733
rect 98283 4684 98284 4724
rect 98324 4684 98325 4724
rect 98283 4675 98325 4684
rect 1152 4556 98784 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 65408 4556
rect 65448 4516 65490 4556
rect 65530 4516 65572 4556
rect 65612 4516 65654 4556
rect 65694 4516 65736 4556
rect 65776 4516 80528 4556
rect 80568 4516 80610 4556
rect 80650 4516 80692 4556
rect 80732 4516 80774 4556
rect 80814 4516 80856 4556
rect 80896 4516 95648 4556
rect 95688 4516 95730 4556
rect 95770 4516 95812 4556
rect 95852 4516 95894 4556
rect 95934 4516 95976 4556
rect 96016 4516 98784 4556
rect 1152 4492 98784 4516
rect 35011 4430 35069 4431
rect 34059 4388 34101 4397
rect 35011 4390 35020 4430
rect 35060 4390 35069 4430
rect 35011 4389 35069 4390
rect 34059 4348 34060 4388
rect 34100 4348 34101 4388
rect 34059 4339 34101 4348
rect 35787 4388 35829 4397
rect 35787 4348 35788 4388
rect 35828 4348 35829 4388
rect 35787 4339 35829 4348
rect 45483 4388 45525 4397
rect 45483 4348 45484 4388
rect 45524 4348 45525 4388
rect 45483 4339 45525 4348
rect 53163 4388 53205 4397
rect 53163 4348 53164 4388
rect 53204 4348 53205 4388
rect 53163 4339 53205 4348
rect 55179 4388 55221 4397
rect 55179 4348 55180 4388
rect 55220 4348 55221 4388
rect 55179 4339 55221 4348
rect 56715 4388 56757 4397
rect 56715 4348 56716 4388
rect 56756 4348 56757 4388
rect 56715 4339 56757 4348
rect 61219 4388 61277 4389
rect 61219 4348 61228 4388
rect 61268 4348 61277 4388
rect 61219 4347 61277 4348
rect 69003 4388 69045 4397
rect 69003 4348 69004 4388
rect 69044 4348 69045 4388
rect 69003 4339 69045 4348
rect 70923 4388 70965 4397
rect 70923 4348 70924 4388
rect 70964 4348 70965 4388
rect 70923 4339 70965 4348
rect 72843 4388 72885 4397
rect 72843 4348 72844 4388
rect 72884 4348 72885 4388
rect 72843 4339 72885 4348
rect 85419 4388 85461 4397
rect 85419 4348 85420 4388
rect 85460 4348 85461 4388
rect 85419 4339 85461 4348
rect 22731 4304 22773 4313
rect 22731 4264 22732 4304
rect 22772 4264 22773 4304
rect 22731 4255 22773 4264
rect 47587 4304 47645 4305
rect 47587 4264 47596 4304
rect 47636 4264 47645 4304
rect 47587 4263 47645 4264
rect 64195 4304 64253 4305
rect 64195 4264 64204 4304
rect 64244 4264 64253 4304
rect 64195 4263 64253 4264
rect 77635 4304 77693 4305
rect 77635 4264 77644 4304
rect 77684 4264 77693 4304
rect 77635 4263 77693 4264
rect 17547 4231 17589 4240
rect 16963 4220 17021 4221
rect 16963 4180 16972 4220
rect 17012 4180 17021 4220
rect 16963 4179 17021 4180
rect 17155 4220 17213 4221
rect 17155 4180 17164 4220
rect 17204 4180 17213 4220
rect 17155 4179 17213 4180
rect 17355 4220 17397 4229
rect 17355 4180 17356 4220
rect 17396 4180 17397 4220
rect 17547 4191 17548 4231
rect 17588 4191 17589 4231
rect 17547 4182 17589 4191
rect 18883 4220 18941 4221
rect 17355 4171 17397 4180
rect 18883 4180 18892 4220
rect 18932 4180 18941 4220
rect 18883 4179 18941 4180
rect 19075 4220 19133 4221
rect 19075 4180 19084 4220
rect 19124 4180 19133 4220
rect 19075 4179 19133 4180
rect 19563 4220 19605 4229
rect 19563 4180 19564 4220
rect 19604 4180 19605 4220
rect 19563 4171 19605 4180
rect 19755 4220 19797 4229
rect 19755 4180 19756 4220
rect 19796 4180 19797 4220
rect 19755 4171 19797 4180
rect 19947 4220 19989 4229
rect 19947 4180 19948 4220
rect 19988 4180 19989 4220
rect 19947 4171 19989 4180
rect 20144 4220 20186 4229
rect 20144 4180 20145 4220
rect 20185 4180 20186 4220
rect 20144 4171 20186 4180
rect 21099 4220 21141 4229
rect 21099 4180 21100 4220
rect 21140 4180 21141 4220
rect 21099 4171 21141 4180
rect 21291 4220 21333 4229
rect 21291 4180 21292 4220
rect 21332 4180 21333 4220
rect 21291 4171 21333 4180
rect 21483 4220 21525 4229
rect 21483 4180 21484 4220
rect 21524 4180 21525 4220
rect 21483 4171 21525 4180
rect 21675 4220 21717 4229
rect 21675 4180 21676 4220
rect 21716 4180 21717 4220
rect 21675 4171 21717 4180
rect 21867 4220 21909 4229
rect 21867 4180 21868 4220
rect 21908 4180 21909 4220
rect 21867 4171 21909 4180
rect 22059 4220 22101 4229
rect 22059 4180 22060 4220
rect 22100 4180 22101 4220
rect 22059 4171 22101 4180
rect 22251 4220 22293 4229
rect 22251 4180 22252 4220
rect 22292 4180 22293 4220
rect 22251 4171 22293 4180
rect 22443 4220 22485 4229
rect 22443 4180 22444 4220
rect 22484 4180 22485 4220
rect 22443 4171 22485 4180
rect 22635 4220 22677 4229
rect 22635 4180 22636 4220
rect 22676 4180 22677 4220
rect 22635 4171 22677 4180
rect 22827 4220 22869 4229
rect 22827 4180 22828 4220
rect 22868 4180 22869 4220
rect 22827 4171 22869 4180
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23829 4220
rect 23787 4171 23829 4180
rect 23979 4220 24021 4229
rect 23979 4180 23980 4220
rect 24020 4180 24021 4220
rect 23979 4171 24021 4180
rect 24171 4220 24213 4229
rect 24171 4180 24172 4220
rect 24212 4180 24213 4220
rect 24171 4171 24213 4180
rect 24363 4220 24405 4229
rect 24363 4180 24364 4220
rect 24404 4180 24405 4220
rect 24363 4171 24405 4180
rect 24555 4220 24597 4229
rect 24555 4180 24556 4220
rect 24596 4180 24597 4220
rect 24555 4171 24597 4180
rect 24747 4220 24789 4229
rect 24747 4180 24748 4220
rect 24788 4180 24789 4220
rect 24747 4171 24789 4180
rect 24939 4220 24981 4229
rect 24939 4180 24940 4220
rect 24980 4180 24981 4220
rect 24939 4171 24981 4180
rect 25131 4220 25173 4229
rect 25131 4180 25132 4220
rect 25172 4180 25173 4220
rect 25131 4171 25173 4180
rect 27243 4220 27285 4229
rect 27243 4180 27244 4220
rect 27284 4180 27285 4220
rect 27243 4171 27285 4180
rect 27435 4220 27477 4229
rect 27435 4180 27436 4220
rect 27476 4180 27477 4220
rect 27435 4171 27477 4180
rect 27627 4220 27669 4229
rect 27627 4180 27628 4220
rect 27668 4180 27669 4220
rect 27627 4171 27669 4180
rect 27819 4220 27861 4229
rect 27819 4180 27820 4220
rect 27860 4180 27861 4220
rect 27819 4171 27861 4180
rect 28011 4220 28053 4229
rect 28011 4180 28012 4220
rect 28052 4180 28053 4220
rect 28011 4171 28053 4180
rect 28203 4220 28245 4229
rect 29443 4220 29501 4221
rect 28203 4180 28204 4220
rect 28244 4180 28245 4220
rect 28203 4171 28245 4180
rect 29251 4219 29309 4220
rect 29251 4179 29260 4219
rect 29300 4179 29309 4219
rect 29443 4180 29452 4220
rect 29492 4180 29501 4220
rect 29443 4179 29501 4180
rect 29931 4220 29973 4229
rect 29931 4180 29932 4220
rect 29972 4180 29973 4220
rect 29251 4178 29309 4179
rect 29931 4171 29973 4180
rect 30123 4220 30165 4229
rect 30123 4180 30124 4220
rect 30164 4180 30165 4220
rect 30123 4171 30165 4180
rect 30315 4220 30357 4229
rect 30315 4180 30316 4220
rect 30356 4180 30357 4220
rect 30315 4171 30357 4180
rect 30507 4220 30549 4229
rect 30507 4180 30508 4220
rect 30548 4180 30549 4220
rect 30507 4171 30549 4180
rect 30699 4220 30741 4229
rect 30699 4180 30700 4220
rect 30740 4180 30741 4220
rect 30699 4171 30741 4180
rect 30891 4220 30933 4229
rect 30891 4180 30892 4220
rect 30932 4180 30933 4220
rect 30891 4171 30933 4180
rect 31083 4220 31125 4229
rect 31083 4180 31084 4220
rect 31124 4180 31125 4220
rect 31083 4171 31125 4180
rect 31275 4220 31317 4229
rect 31275 4180 31276 4220
rect 31316 4180 31317 4220
rect 31275 4171 31317 4180
rect 33859 4220 33917 4221
rect 33859 4180 33868 4220
rect 33908 4180 33917 4220
rect 33859 4179 33917 4180
rect 34051 4220 34109 4221
rect 34051 4180 34060 4220
rect 34100 4180 34109 4220
rect 34051 4179 34109 4180
rect 34435 4220 34493 4221
rect 34435 4180 34444 4220
rect 34484 4180 34493 4220
rect 34435 4179 34493 4180
rect 34627 4220 34685 4221
rect 34627 4180 34636 4220
rect 34676 4180 34685 4220
rect 34627 4179 34685 4180
rect 35011 4220 35069 4221
rect 35011 4180 35020 4220
rect 35060 4180 35069 4220
rect 35011 4179 35069 4180
rect 35203 4220 35261 4221
rect 35779 4220 35837 4221
rect 35203 4180 35212 4220
rect 35252 4180 35261 4220
rect 35203 4179 35261 4180
rect 35579 4219 35637 4220
rect 35579 4179 35588 4219
rect 35628 4179 35637 4219
rect 35779 4180 35788 4220
rect 35828 4180 35837 4220
rect 35779 4179 35837 4180
rect 37611 4220 37653 4229
rect 37611 4180 37612 4220
rect 37652 4180 37653 4220
rect 35579 4178 35637 4179
rect 37611 4171 37653 4180
rect 37803 4220 37845 4229
rect 37803 4180 37804 4220
rect 37844 4180 37845 4220
rect 37803 4171 37845 4180
rect 37995 4220 38037 4229
rect 37995 4180 37996 4220
rect 38036 4180 38037 4220
rect 37995 4171 38037 4180
rect 38187 4220 38229 4229
rect 38187 4180 38188 4220
rect 38228 4180 38229 4220
rect 38187 4171 38229 4180
rect 38379 4220 38421 4229
rect 38379 4180 38380 4220
rect 38420 4180 38421 4220
rect 38379 4171 38421 4180
rect 38571 4220 38613 4229
rect 38571 4180 38572 4220
rect 38612 4180 38613 4220
rect 38571 4171 38613 4180
rect 38763 4220 38805 4229
rect 38763 4180 38764 4220
rect 38804 4180 38805 4220
rect 38763 4171 38805 4180
rect 38955 4220 38997 4229
rect 38955 4180 38956 4220
rect 38996 4180 38997 4220
rect 38955 4171 38997 4180
rect 39147 4220 39189 4229
rect 39147 4180 39148 4220
rect 39188 4180 39189 4220
rect 39147 4171 39189 4180
rect 39339 4220 39381 4229
rect 39339 4180 39340 4220
rect 39380 4180 39381 4220
rect 39339 4171 39381 4180
rect 44619 4220 44661 4229
rect 44619 4180 44620 4220
rect 44660 4180 44661 4220
rect 44619 4171 44661 4180
rect 45955 4220 46013 4221
rect 45955 4180 45964 4220
rect 46004 4180 46013 4220
rect 45955 4179 46013 4180
rect 47115 4220 47157 4229
rect 47115 4180 47116 4220
rect 47156 4180 47157 4220
rect 47115 4171 47157 4180
rect 48451 4220 48509 4221
rect 48451 4180 48460 4220
rect 48500 4180 48509 4220
rect 48451 4179 48509 4180
rect 49035 4220 49077 4229
rect 49035 4180 49036 4220
rect 49076 4180 49077 4220
rect 49035 4171 49077 4180
rect 49227 4220 49269 4229
rect 49227 4180 49228 4220
rect 49268 4180 49269 4220
rect 49227 4171 49269 4180
rect 49515 4217 49557 4226
rect 49515 4177 49516 4217
rect 49556 4177 49557 4217
rect 49515 4168 49557 4177
rect 49995 4220 50037 4229
rect 49995 4180 49996 4220
rect 50036 4180 50037 4220
rect 49995 4171 50037 4180
rect 51531 4220 51573 4229
rect 51531 4180 51532 4220
rect 51572 4180 51573 4220
rect 51531 4171 51573 4180
rect 52011 4220 52053 4229
rect 52011 4180 52012 4220
rect 52052 4180 52053 4220
rect 52011 4171 52053 4180
rect 52107 4220 52149 4229
rect 52107 4180 52108 4220
rect 52148 4180 52149 4220
rect 52107 4171 52149 4180
rect 52195 4220 52253 4221
rect 52195 4180 52204 4220
rect 52244 4180 52253 4220
rect 52195 4179 52253 4180
rect 52395 4220 52437 4229
rect 52395 4180 52396 4220
rect 52436 4180 52437 4220
rect 52395 4171 52437 4180
rect 52587 4220 52629 4229
rect 52587 4180 52588 4220
rect 52628 4180 52629 4220
rect 52587 4171 52629 4180
rect 52971 4220 53013 4229
rect 52971 4180 52972 4220
rect 53012 4180 53013 4220
rect 52971 4171 53013 4180
rect 53355 4220 53397 4229
rect 53355 4180 53356 4220
rect 53396 4180 53397 4220
rect 53355 4171 53397 4180
rect 53547 4220 53589 4229
rect 53547 4180 53548 4220
rect 53588 4180 53589 4220
rect 53547 4171 53589 4180
rect 54595 4220 54653 4221
rect 54595 4180 54604 4220
rect 54644 4180 54653 4220
rect 54595 4179 54653 4180
rect 54787 4220 54845 4221
rect 54787 4180 54796 4220
rect 54836 4180 54845 4220
rect 54787 4179 54845 4180
rect 55083 4220 55125 4229
rect 55083 4180 55084 4220
rect 55124 4180 55125 4220
rect 55083 4171 55125 4180
rect 55275 4220 55317 4229
rect 55275 4180 55276 4220
rect 55316 4180 55317 4220
rect 55275 4171 55317 4180
rect 56523 4220 56565 4229
rect 56523 4180 56524 4220
rect 56564 4180 56565 4220
rect 56523 4171 56565 4180
rect 57003 4220 57045 4229
rect 57003 4180 57004 4220
rect 57044 4180 57045 4220
rect 57003 4171 57045 4180
rect 57579 4220 57621 4229
rect 57579 4180 57580 4220
rect 57620 4180 57621 4220
rect 57579 4171 57621 4180
rect 57955 4220 58013 4221
rect 57955 4180 57964 4220
rect 58004 4180 58013 4220
rect 57955 4179 58013 4180
rect 58827 4220 58869 4229
rect 58827 4180 58828 4220
rect 58868 4180 58869 4220
rect 58827 4171 58869 4180
rect 59203 4220 59261 4221
rect 59203 4180 59212 4220
rect 59252 4180 59261 4220
rect 59203 4179 59261 4180
rect 60163 4220 60221 4221
rect 60163 4180 60172 4220
rect 60212 4180 60221 4220
rect 60643 4220 60701 4221
rect 60163 4179 60221 4180
rect 60451 4209 60509 4210
rect 60451 4169 60460 4209
rect 60500 4169 60509 4209
rect 60643 4180 60652 4220
rect 60692 4180 60701 4220
rect 60643 4179 60701 4180
rect 60939 4220 60981 4229
rect 60939 4180 60940 4220
rect 60980 4180 60981 4220
rect 60939 4171 60981 4180
rect 61035 4220 61077 4229
rect 61035 4180 61036 4220
rect 61076 4180 61077 4220
rect 61035 4171 61077 4180
rect 63435 4220 63477 4229
rect 63435 4180 63436 4220
rect 63476 4180 63477 4220
rect 63435 4171 63477 4180
rect 64579 4220 64637 4221
rect 64579 4180 64588 4220
rect 64628 4180 64637 4220
rect 64579 4179 64637 4180
rect 64771 4220 64829 4221
rect 64771 4180 64780 4220
rect 64820 4180 64829 4220
rect 64771 4179 64829 4180
rect 66883 4220 66941 4221
rect 66883 4180 66892 4220
rect 66932 4180 66941 4220
rect 66883 4179 66941 4180
rect 67075 4220 67133 4221
rect 67075 4180 67084 4220
rect 67124 4180 67133 4220
rect 67075 4179 67133 4180
rect 67755 4220 67797 4229
rect 67755 4180 67756 4220
rect 67796 4180 67797 4220
rect 67755 4171 67797 4180
rect 67947 4220 67989 4229
rect 67947 4180 67948 4220
rect 67988 4180 67989 4220
rect 67947 4171 67989 4180
rect 68139 4220 68181 4229
rect 68139 4180 68140 4220
rect 68180 4180 68181 4220
rect 68139 4171 68181 4180
rect 68331 4220 68373 4229
rect 68331 4180 68332 4220
rect 68372 4180 68373 4220
rect 68331 4171 68373 4180
rect 68523 4220 68565 4229
rect 68523 4180 68524 4220
rect 68564 4180 68565 4220
rect 68523 4171 68565 4180
rect 68715 4220 68757 4229
rect 68715 4180 68716 4220
rect 68756 4180 68757 4220
rect 68715 4171 68757 4180
rect 68907 4220 68949 4229
rect 68907 4180 68908 4220
rect 68948 4180 68949 4220
rect 68907 4171 68949 4180
rect 69099 4220 69141 4229
rect 69099 4180 69100 4220
rect 69140 4180 69141 4220
rect 69099 4171 69141 4180
rect 70059 4220 70101 4229
rect 70059 4180 70060 4220
rect 70100 4180 70101 4220
rect 70059 4171 70101 4180
rect 70251 4220 70293 4229
rect 70251 4180 70252 4220
rect 70292 4180 70293 4220
rect 70251 4171 70293 4180
rect 70443 4220 70485 4229
rect 70443 4180 70444 4220
rect 70484 4180 70485 4220
rect 70443 4171 70485 4180
rect 70635 4220 70677 4229
rect 70635 4180 70636 4220
rect 70676 4180 70677 4220
rect 70635 4171 70677 4180
rect 70827 4220 70869 4229
rect 70827 4180 70828 4220
rect 70868 4180 70869 4220
rect 70827 4171 70869 4180
rect 71019 4220 71061 4229
rect 71019 4180 71020 4220
rect 71060 4180 71061 4220
rect 71019 4171 71061 4180
rect 71211 4220 71253 4229
rect 71211 4180 71212 4220
rect 71252 4180 71253 4220
rect 71211 4171 71253 4180
rect 71403 4220 71445 4229
rect 71403 4180 71404 4220
rect 71444 4180 71445 4220
rect 71403 4171 71445 4180
rect 71595 4220 71637 4229
rect 71595 4180 71596 4220
rect 71636 4180 71637 4220
rect 71595 4171 71637 4180
rect 71787 4220 71829 4229
rect 71787 4180 71788 4220
rect 71828 4180 71829 4220
rect 71787 4171 71829 4180
rect 71979 4220 72021 4229
rect 71979 4180 71980 4220
rect 72020 4180 72021 4220
rect 71979 4171 72021 4180
rect 72171 4220 72213 4229
rect 72171 4180 72172 4220
rect 72212 4180 72213 4220
rect 72171 4171 72213 4180
rect 72747 4220 72789 4229
rect 72747 4180 72748 4220
rect 72788 4180 72789 4220
rect 72747 4171 72789 4180
rect 72939 4220 72981 4229
rect 72939 4180 72940 4220
rect 72980 4180 72981 4220
rect 72939 4171 72981 4180
rect 73131 4220 73173 4229
rect 73131 4180 73132 4220
rect 73172 4180 73173 4220
rect 73131 4171 73173 4180
rect 73323 4220 73365 4229
rect 73323 4180 73324 4220
rect 73364 4180 73365 4220
rect 73323 4171 73365 4180
rect 73515 4220 73557 4229
rect 73515 4180 73516 4220
rect 73556 4180 73557 4220
rect 73515 4171 73557 4180
rect 73707 4220 73749 4229
rect 73707 4180 73708 4220
rect 73748 4180 73749 4220
rect 73707 4171 73749 4180
rect 74667 4220 74709 4229
rect 74667 4180 74668 4220
rect 74708 4180 74709 4220
rect 74667 4171 74709 4180
rect 74859 4220 74901 4229
rect 74859 4180 74860 4220
rect 74900 4180 74901 4220
rect 74859 4171 74901 4180
rect 75819 4220 75861 4229
rect 75819 4180 75820 4220
rect 75860 4180 75861 4220
rect 75819 4171 75861 4180
rect 76011 4220 76053 4229
rect 76011 4180 76012 4220
rect 76052 4180 76053 4220
rect 76011 4171 76053 4180
rect 76587 4220 76629 4229
rect 76587 4180 76588 4220
rect 76628 4180 76629 4220
rect 76587 4171 76629 4180
rect 76779 4220 76821 4229
rect 76779 4180 76780 4220
rect 76820 4180 76821 4220
rect 76779 4171 76821 4180
rect 77155 4220 77213 4221
rect 77155 4180 77164 4220
rect 77204 4180 77213 4220
rect 77155 4179 77213 4180
rect 77347 4220 77405 4221
rect 77347 4180 77356 4220
rect 77396 4180 77405 4220
rect 77347 4179 77405 4180
rect 78411 4220 78453 4229
rect 78411 4180 78412 4220
rect 78452 4180 78453 4220
rect 78411 4171 78453 4180
rect 78795 4220 78837 4229
rect 78795 4180 78796 4220
rect 78836 4180 78837 4220
rect 78795 4171 78837 4180
rect 78987 4220 79029 4229
rect 78987 4180 78988 4220
rect 79028 4180 79029 4220
rect 78987 4171 79029 4180
rect 80715 4220 80757 4229
rect 80715 4180 80716 4220
rect 80756 4180 80757 4220
rect 80715 4171 80757 4180
rect 80907 4220 80949 4229
rect 80907 4180 80908 4220
rect 80948 4180 80949 4220
rect 80907 4171 80949 4180
rect 81283 4220 81341 4221
rect 81283 4180 81292 4220
rect 81332 4180 81341 4220
rect 81283 4179 81341 4180
rect 83211 4220 83253 4229
rect 83211 4180 83212 4220
rect 83252 4180 83253 4220
rect 83211 4171 83253 4180
rect 83403 4220 83445 4229
rect 83403 4180 83404 4220
rect 83444 4180 83445 4220
rect 83403 4171 83445 4180
rect 84267 4220 84309 4229
rect 84267 4180 84268 4220
rect 84308 4180 84309 4220
rect 84267 4171 84309 4180
rect 85323 4220 85365 4229
rect 85323 4180 85324 4220
rect 85364 4180 85365 4220
rect 85323 4171 85365 4180
rect 85515 4220 85557 4229
rect 85515 4180 85516 4220
rect 85556 4180 85557 4220
rect 85515 4171 85557 4180
rect 60451 4168 60509 4169
rect 36451 4149 36509 4150
rect 1507 4136 1565 4137
rect 1507 4096 1516 4136
rect 1556 4096 1565 4136
rect 1507 4095 1565 4096
rect 1891 4136 1949 4137
rect 1891 4096 1900 4136
rect 1940 4096 1949 4136
rect 1891 4095 1949 4096
rect 2275 4136 2333 4137
rect 2275 4096 2284 4136
rect 2324 4096 2333 4136
rect 2275 4095 2333 4096
rect 2659 4136 2717 4137
rect 2659 4096 2668 4136
rect 2708 4096 2717 4136
rect 2659 4095 2717 4096
rect 3043 4136 3101 4137
rect 3043 4096 3052 4136
rect 3092 4096 3101 4136
rect 3043 4095 3101 4096
rect 3427 4136 3485 4137
rect 3427 4096 3436 4136
rect 3476 4096 3485 4136
rect 3427 4095 3485 4096
rect 3811 4136 3869 4137
rect 3811 4096 3820 4136
rect 3860 4096 3869 4136
rect 3811 4095 3869 4096
rect 4195 4136 4253 4137
rect 4195 4096 4204 4136
rect 4244 4096 4253 4136
rect 4195 4095 4253 4096
rect 4579 4136 4637 4137
rect 4579 4096 4588 4136
rect 4628 4096 4637 4136
rect 4579 4095 4637 4096
rect 4963 4136 5021 4137
rect 4963 4096 4972 4136
rect 5012 4096 5021 4136
rect 4963 4095 5021 4096
rect 5347 4136 5405 4137
rect 5347 4096 5356 4136
rect 5396 4096 5405 4136
rect 5347 4095 5405 4096
rect 5731 4136 5789 4137
rect 5731 4096 5740 4136
rect 5780 4096 5789 4136
rect 5731 4095 5789 4096
rect 6115 4136 6173 4137
rect 6115 4096 6124 4136
rect 6164 4096 6173 4136
rect 6115 4095 6173 4096
rect 6499 4136 6557 4137
rect 6499 4096 6508 4136
rect 6548 4096 6557 4136
rect 6499 4095 6557 4096
rect 6883 4136 6941 4137
rect 6883 4096 6892 4136
rect 6932 4096 6941 4136
rect 6883 4095 6941 4096
rect 7267 4136 7325 4137
rect 7267 4096 7276 4136
rect 7316 4096 7325 4136
rect 7267 4095 7325 4096
rect 7651 4136 7709 4137
rect 7651 4096 7660 4136
rect 7700 4096 7709 4136
rect 7651 4095 7709 4096
rect 8035 4136 8093 4137
rect 8035 4096 8044 4136
rect 8084 4096 8093 4136
rect 8035 4095 8093 4096
rect 8419 4136 8477 4137
rect 8419 4096 8428 4136
rect 8468 4096 8477 4136
rect 8419 4095 8477 4096
rect 8803 4136 8861 4137
rect 8803 4096 8812 4136
rect 8852 4096 8861 4136
rect 8803 4095 8861 4096
rect 9187 4136 9245 4137
rect 9187 4096 9196 4136
rect 9236 4096 9245 4136
rect 9187 4095 9245 4096
rect 9571 4136 9629 4137
rect 9571 4096 9580 4136
rect 9620 4096 9629 4136
rect 9571 4095 9629 4096
rect 9955 4136 10013 4137
rect 9955 4096 9964 4136
rect 10004 4096 10013 4136
rect 9955 4095 10013 4096
rect 10339 4136 10397 4137
rect 10339 4096 10348 4136
rect 10388 4096 10397 4136
rect 10339 4095 10397 4096
rect 10723 4136 10781 4137
rect 10723 4096 10732 4136
rect 10772 4096 10781 4136
rect 10723 4095 10781 4096
rect 11107 4136 11165 4137
rect 11107 4096 11116 4136
rect 11156 4096 11165 4136
rect 11107 4095 11165 4096
rect 11491 4136 11549 4137
rect 11491 4096 11500 4136
rect 11540 4096 11549 4136
rect 11491 4095 11549 4096
rect 11875 4136 11933 4137
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 11875 4095 11933 4096
rect 12259 4136 12317 4137
rect 12259 4096 12268 4136
rect 12308 4096 12317 4136
rect 12259 4095 12317 4096
rect 12643 4136 12701 4137
rect 12643 4096 12652 4136
rect 12692 4096 12701 4136
rect 12643 4095 12701 4096
rect 13027 4136 13085 4137
rect 13027 4096 13036 4136
rect 13076 4096 13085 4136
rect 13027 4095 13085 4096
rect 13411 4136 13469 4137
rect 13411 4096 13420 4136
rect 13460 4096 13469 4136
rect 13411 4095 13469 4096
rect 13795 4136 13853 4137
rect 13795 4096 13804 4136
rect 13844 4096 13853 4136
rect 13795 4095 13853 4096
rect 14179 4136 14237 4137
rect 14179 4096 14188 4136
rect 14228 4096 14237 4136
rect 14179 4095 14237 4096
rect 14563 4136 14621 4137
rect 14563 4096 14572 4136
rect 14612 4096 14621 4136
rect 14563 4095 14621 4096
rect 14947 4136 15005 4137
rect 14947 4096 14956 4136
rect 14996 4096 15005 4136
rect 14947 4095 15005 4096
rect 15331 4136 15389 4137
rect 15331 4096 15340 4136
rect 15380 4096 15389 4136
rect 15331 4095 15389 4096
rect 15715 4136 15773 4137
rect 15715 4096 15724 4136
rect 15764 4096 15773 4136
rect 15715 4095 15773 4096
rect 16099 4136 16157 4137
rect 16099 4096 16108 4136
rect 16148 4096 16157 4136
rect 16099 4095 16157 4096
rect 16483 4136 16541 4137
rect 16483 4096 16492 4136
rect 16532 4096 16541 4136
rect 16483 4095 16541 4096
rect 17731 4136 17789 4137
rect 17731 4096 17740 4136
rect 17780 4096 17789 4136
rect 17731 4095 17789 4096
rect 18115 4136 18173 4137
rect 18115 4096 18124 4136
rect 18164 4096 18173 4136
rect 18115 4095 18173 4096
rect 18499 4136 18557 4137
rect 18499 4096 18508 4136
rect 18548 4096 18557 4136
rect 18499 4095 18557 4096
rect 20323 4136 20381 4137
rect 20323 4096 20332 4136
rect 20372 4096 20381 4136
rect 20323 4095 20381 4096
rect 20707 4136 20765 4137
rect 20707 4096 20716 4136
rect 20756 4096 20765 4136
rect 20707 4095 20765 4096
rect 22347 4136 22389 4145
rect 22347 4096 22348 4136
rect 22388 4096 22389 4136
rect 22347 4087 22389 4096
rect 23011 4136 23069 4137
rect 23011 4096 23020 4136
rect 23060 4096 23069 4136
rect 23011 4095 23069 4096
rect 23395 4136 23453 4137
rect 23395 4096 23404 4136
rect 23444 4096 23453 4136
rect 23395 4095 23453 4096
rect 24267 4136 24309 4145
rect 24267 4096 24268 4136
rect 24308 4096 24309 4136
rect 24267 4087 24309 4096
rect 25035 4136 25077 4145
rect 25035 4096 25036 4136
rect 25076 4096 25077 4136
rect 25035 4087 25077 4096
rect 25315 4136 25373 4137
rect 25315 4096 25324 4136
rect 25364 4096 25373 4136
rect 25315 4095 25373 4096
rect 25699 4136 25757 4137
rect 25699 4096 25708 4136
rect 25748 4096 25757 4136
rect 25699 4095 25757 4096
rect 26083 4136 26141 4137
rect 26083 4096 26092 4136
rect 26132 4096 26141 4136
rect 26083 4095 26141 4096
rect 26467 4136 26525 4137
rect 26467 4096 26476 4136
rect 26516 4096 26525 4136
rect 26467 4095 26525 4096
rect 26851 4136 26909 4137
rect 26851 4096 26860 4136
rect 26900 4096 26909 4136
rect 26851 4095 26909 4096
rect 28387 4136 28445 4137
rect 28387 4096 28396 4136
rect 28436 4096 28445 4136
rect 28387 4095 28445 4096
rect 28771 4136 28829 4137
rect 28771 4096 28780 4136
rect 28820 4096 28829 4136
rect 28771 4095 28829 4096
rect 31179 4136 31221 4145
rect 31179 4096 31180 4136
rect 31220 4096 31221 4136
rect 31179 4087 31221 4096
rect 31459 4136 31517 4137
rect 31459 4096 31468 4136
rect 31508 4096 31517 4136
rect 31459 4095 31517 4096
rect 31843 4136 31901 4137
rect 31843 4096 31852 4136
rect 31892 4096 31901 4136
rect 31843 4095 31901 4096
rect 32227 4136 32285 4137
rect 32227 4096 32236 4136
rect 32276 4096 32285 4136
rect 32227 4095 32285 4096
rect 32611 4136 32669 4137
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32611 4095 32669 4096
rect 32995 4136 33053 4137
rect 32995 4096 33004 4136
rect 33044 4096 33053 4136
rect 32995 4095 33053 4096
rect 33379 4136 33437 4137
rect 33379 4096 33388 4136
rect 33428 4096 33437 4136
rect 33379 4095 33437 4096
rect 36067 4136 36125 4137
rect 36067 4096 36076 4136
rect 36116 4096 36125 4136
rect 36451 4109 36460 4149
rect 36500 4109 36509 4149
rect 37219 4149 37277 4150
rect 36451 4108 36509 4109
rect 36835 4136 36893 4137
rect 36067 4095 36125 4096
rect 36835 4096 36844 4136
rect 36884 4096 36893 4136
rect 37219 4109 37228 4149
rect 37268 4109 37277 4149
rect 37219 4108 37277 4109
rect 39523 4149 39581 4150
rect 39523 4109 39532 4149
rect 39572 4109 39581 4149
rect 88963 4149 89021 4150
rect 39523 4108 39581 4109
rect 39907 4136 39965 4137
rect 36835 4095 36893 4096
rect 39907 4096 39916 4136
rect 39956 4096 39965 4136
rect 39907 4095 39965 4096
rect 40291 4136 40349 4137
rect 40291 4096 40300 4136
rect 40340 4096 40349 4136
rect 40291 4095 40349 4096
rect 40675 4136 40733 4137
rect 40675 4096 40684 4136
rect 40724 4096 40733 4136
rect 40675 4095 40733 4096
rect 41059 4136 41117 4137
rect 41059 4096 41068 4136
rect 41108 4096 41117 4136
rect 41059 4095 41117 4096
rect 41443 4136 41501 4137
rect 41443 4096 41452 4136
rect 41492 4096 41501 4136
rect 41443 4095 41501 4096
rect 41827 4136 41885 4137
rect 41827 4096 41836 4136
rect 41876 4096 41885 4136
rect 41827 4095 41885 4096
rect 42211 4136 42269 4137
rect 42211 4096 42220 4136
rect 42260 4096 42269 4136
rect 42211 4095 42269 4096
rect 42595 4136 42653 4137
rect 42595 4096 42604 4136
rect 42644 4096 42653 4136
rect 42595 4095 42653 4096
rect 42979 4136 43037 4137
rect 42979 4096 42988 4136
rect 43028 4096 43037 4136
rect 42979 4095 43037 4096
rect 43363 4136 43421 4137
rect 43363 4096 43372 4136
rect 43412 4096 43421 4136
rect 43363 4095 43421 4096
rect 50851 4136 50909 4137
rect 50851 4096 50860 4136
rect 50900 4096 50909 4136
rect 50851 4095 50909 4096
rect 51235 4136 51293 4137
rect 51235 4096 51244 4136
rect 51284 4096 51293 4136
rect 51235 4095 51293 4096
rect 51723 4136 51765 4145
rect 51723 4096 51724 4136
rect 51764 4096 51765 4136
rect 51723 4087 51765 4096
rect 53923 4136 53981 4137
rect 53923 4096 53932 4136
rect 53972 4096 53981 4136
rect 53923 4095 53981 4096
rect 54307 4136 54365 4137
rect 54307 4096 54316 4136
rect 54356 4096 54365 4136
rect 54307 4095 54365 4096
rect 55651 4136 55709 4137
rect 55651 4096 55660 4136
rect 55700 4096 55709 4136
rect 55651 4095 55709 4096
rect 56035 4136 56093 4137
rect 56035 4096 56044 4136
rect 56084 4096 56093 4136
rect 56035 4095 56093 4096
rect 61603 4136 61661 4137
rect 61603 4096 61612 4136
rect 61652 4096 61661 4136
rect 61603 4095 61661 4096
rect 61987 4136 62045 4137
rect 61987 4096 61996 4136
rect 62036 4096 62045 4136
rect 61987 4095 62045 4096
rect 62371 4136 62429 4137
rect 62371 4096 62380 4136
rect 62420 4096 62429 4136
rect 62371 4095 62429 4096
rect 62755 4136 62813 4137
rect 62755 4096 62764 4136
rect 62804 4096 62813 4136
rect 62755 4095 62813 4096
rect 65251 4136 65309 4137
rect 65251 4096 65260 4136
rect 65300 4096 65309 4136
rect 65251 4095 65309 4096
rect 65635 4136 65693 4137
rect 65635 4096 65644 4136
rect 65684 4096 65693 4136
rect 65635 4095 65693 4096
rect 66019 4136 66077 4137
rect 66019 4096 66028 4136
rect 66068 4096 66077 4136
rect 66019 4095 66077 4096
rect 66403 4136 66461 4137
rect 66403 4096 66412 4136
rect 66452 4096 66461 4136
rect 66403 4095 66461 4096
rect 67555 4136 67613 4137
rect 67555 4096 67564 4136
rect 67604 4096 67613 4136
rect 67555 4095 67613 4096
rect 69475 4136 69533 4137
rect 69475 4096 69484 4136
rect 69524 4096 69533 4136
rect 69475 4095 69533 4096
rect 69859 4136 69917 4137
rect 69859 4096 69868 4136
rect 69908 4096 69917 4136
rect 69859 4095 69917 4096
rect 71307 4136 71349 4145
rect 71307 4096 71308 4136
rect 71348 4096 71349 4136
rect 71307 4087 71349 4096
rect 72547 4136 72605 4137
rect 72547 4096 72556 4136
rect 72596 4096 72605 4136
rect 72547 4095 72605 4096
rect 74083 4136 74141 4137
rect 74083 4096 74092 4136
rect 74132 4096 74141 4136
rect 74083 4095 74141 4096
rect 74467 4136 74525 4137
rect 74467 4096 74476 4136
rect 74516 4096 74525 4136
rect 74467 4095 74525 4096
rect 75235 4136 75293 4137
rect 75235 4096 75244 4136
rect 75284 4096 75293 4136
rect 75235 4095 75293 4096
rect 75619 4136 75677 4137
rect 75619 4096 75628 4136
rect 75668 4096 75677 4136
rect 75619 4095 75677 4096
rect 76387 4136 76445 4137
rect 76387 4096 76396 4136
rect 76436 4096 76445 4136
rect 76387 4095 76445 4096
rect 79363 4136 79421 4137
rect 79363 4096 79372 4136
rect 79412 4096 79421 4136
rect 79363 4095 79421 4096
rect 79747 4136 79805 4137
rect 79747 4096 79756 4136
rect 79796 4096 79805 4136
rect 79747 4095 79805 4096
rect 80131 4136 80189 4137
rect 80131 4096 80140 4136
rect 80180 4096 80189 4136
rect 80131 4095 80189 4096
rect 80515 4136 80573 4137
rect 80515 4096 80524 4136
rect 80564 4096 80573 4136
rect 80515 4095 80573 4096
rect 82627 4136 82685 4137
rect 82627 4096 82636 4136
rect 82676 4096 82685 4136
rect 82627 4095 82685 4096
rect 83011 4136 83069 4137
rect 83011 4096 83020 4136
rect 83060 4096 83069 4136
rect 83011 4095 83069 4096
rect 83779 4136 83837 4137
rect 83779 4096 83788 4136
rect 83828 4096 83837 4136
rect 83779 4095 83837 4096
rect 85891 4136 85949 4137
rect 85891 4096 85900 4136
rect 85940 4096 85949 4136
rect 85891 4095 85949 4096
rect 86275 4136 86333 4137
rect 86275 4096 86284 4136
rect 86324 4096 86333 4136
rect 86275 4095 86333 4096
rect 86659 4136 86717 4137
rect 86659 4096 86668 4136
rect 86708 4096 86717 4136
rect 86659 4095 86717 4096
rect 87043 4136 87101 4137
rect 87043 4096 87052 4136
rect 87092 4096 87101 4136
rect 87043 4095 87101 4096
rect 87427 4136 87485 4137
rect 87427 4096 87436 4136
rect 87476 4096 87485 4136
rect 87427 4095 87485 4096
rect 87811 4136 87869 4137
rect 87811 4096 87820 4136
rect 87860 4096 87869 4136
rect 87811 4095 87869 4096
rect 88195 4136 88253 4137
rect 88195 4096 88204 4136
rect 88244 4096 88253 4136
rect 88195 4095 88253 4096
rect 88579 4136 88637 4137
rect 88579 4096 88588 4136
rect 88628 4096 88637 4136
rect 88963 4109 88972 4149
rect 89012 4109 89021 4149
rect 97411 4149 97469 4150
rect 88963 4108 89021 4109
rect 89347 4136 89405 4137
rect 88579 4095 88637 4096
rect 89347 4096 89356 4136
rect 89396 4096 89405 4136
rect 89347 4095 89405 4096
rect 89731 4136 89789 4137
rect 89731 4096 89740 4136
rect 89780 4096 89789 4136
rect 89731 4095 89789 4096
rect 90115 4136 90173 4137
rect 90115 4096 90124 4136
rect 90164 4096 90173 4136
rect 90115 4095 90173 4096
rect 90499 4136 90557 4137
rect 90499 4096 90508 4136
rect 90548 4096 90557 4136
rect 90499 4095 90557 4096
rect 90883 4136 90941 4137
rect 90883 4096 90892 4136
rect 90932 4096 90941 4136
rect 90883 4095 90941 4096
rect 91267 4136 91325 4137
rect 91267 4096 91276 4136
rect 91316 4096 91325 4136
rect 91267 4095 91325 4096
rect 91651 4136 91709 4137
rect 91651 4096 91660 4136
rect 91700 4096 91709 4136
rect 91651 4095 91709 4096
rect 92035 4136 92093 4137
rect 92035 4096 92044 4136
rect 92084 4096 92093 4136
rect 92035 4095 92093 4096
rect 92419 4136 92477 4137
rect 92419 4096 92428 4136
rect 92468 4096 92477 4136
rect 92419 4095 92477 4096
rect 92803 4136 92861 4137
rect 92803 4096 92812 4136
rect 92852 4096 92861 4136
rect 92803 4095 92861 4096
rect 93187 4136 93245 4137
rect 93187 4096 93196 4136
rect 93236 4096 93245 4136
rect 93187 4095 93245 4096
rect 93571 4136 93629 4137
rect 93571 4096 93580 4136
rect 93620 4096 93629 4136
rect 93571 4095 93629 4096
rect 93955 4136 94013 4137
rect 93955 4096 93964 4136
rect 94004 4096 94013 4136
rect 93955 4095 94013 4096
rect 94339 4136 94397 4137
rect 94339 4096 94348 4136
rect 94388 4096 94397 4136
rect 94339 4095 94397 4096
rect 94723 4136 94781 4137
rect 94723 4096 94732 4136
rect 94772 4096 94781 4136
rect 94723 4095 94781 4096
rect 95107 4136 95165 4137
rect 95107 4096 95116 4136
rect 95156 4096 95165 4136
rect 95107 4095 95165 4096
rect 95491 4136 95549 4137
rect 95491 4096 95500 4136
rect 95540 4096 95549 4136
rect 95491 4095 95549 4096
rect 95875 4136 95933 4137
rect 95875 4096 95884 4136
rect 95924 4096 95933 4136
rect 95875 4095 95933 4096
rect 96259 4136 96317 4137
rect 96259 4096 96268 4136
rect 96308 4096 96317 4136
rect 96259 4095 96317 4096
rect 96643 4136 96701 4137
rect 96643 4096 96652 4136
rect 96692 4096 96701 4136
rect 96643 4095 96701 4096
rect 97027 4136 97085 4137
rect 97027 4096 97036 4136
rect 97076 4096 97085 4136
rect 97411 4109 97420 4149
rect 97460 4109 97469 4149
rect 97411 4108 97469 4109
rect 97795 4136 97853 4137
rect 97027 4095 97085 4096
rect 97795 4096 97804 4136
rect 97844 4096 97853 4136
rect 97795 4095 97853 4096
rect 98179 4136 98237 4137
rect 98179 4096 98188 4136
rect 98228 4096 98237 4136
rect 98179 4095 98237 4096
rect 98563 4136 98621 4137
rect 98563 4096 98572 4136
rect 98612 4096 98621 4136
rect 98563 4095 98621 4096
rect 21099 4052 21141 4061
rect 21099 4012 21100 4052
rect 21140 4012 21141 4052
rect 21099 4003 21141 4012
rect 23979 4052 24021 4061
rect 23979 4012 23980 4052
rect 24020 4012 24021 4052
rect 23979 4003 24021 4012
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 29259 4052 29301 4061
rect 29259 4012 29260 4052
rect 29300 4012 29301 4052
rect 29259 4003 29301 4012
rect 30891 4052 30933 4061
rect 30891 4012 30892 4052
rect 30932 4012 30933 4052
rect 30891 4003 30933 4012
rect 34443 4052 34485 4061
rect 34443 4012 34444 4052
rect 34484 4012 34485 4052
rect 34443 4003 34485 4012
rect 38571 4052 38613 4061
rect 38571 4012 38572 4052
rect 38612 4012 38613 4052
rect 38571 4003 38613 4012
rect 42795 4052 42837 4061
rect 42795 4012 42796 4052
rect 42836 4012 42837 4052
rect 42795 4003 42837 4012
rect 49515 4052 49557 4061
rect 49515 4012 49516 4052
rect 49556 4012 49557 4052
rect 49515 4003 49557 4012
rect 49995 4052 50037 4061
rect 49995 4012 49996 4052
rect 50036 4012 50037 4052
rect 49995 4003 50037 4012
rect 50187 4052 50229 4061
rect 50187 4012 50188 4052
rect 50228 4012 50229 4052
rect 50187 4003 50229 4012
rect 51627 4052 51669 4061
rect 51627 4012 51628 4052
rect 51668 4012 51669 4052
rect 51627 4003 51669 4012
rect 52971 4052 53013 4061
rect 52971 4012 52972 4052
rect 53012 4012 53013 4052
rect 52971 4003 53013 4012
rect 56523 4052 56565 4061
rect 56523 4012 56524 4052
rect 56564 4012 56565 4052
rect 56523 4003 56565 4012
rect 57003 4052 57045 4061
rect 57003 4012 57004 4052
rect 57044 4012 57045 4052
rect 57003 4003 57045 4012
rect 57579 4052 57621 4061
rect 57579 4012 57580 4052
rect 57620 4012 57621 4052
rect 57579 4003 57621 4012
rect 60459 4052 60501 4061
rect 60459 4012 60460 4052
rect 60500 4012 60501 4052
rect 60459 4003 60501 4012
rect 63627 4052 63669 4061
rect 63627 4012 63628 4052
rect 63668 4012 63669 4052
rect 63627 4003 63669 4012
rect 64779 4052 64821 4061
rect 64779 4012 64780 4052
rect 64820 4012 64821 4052
rect 64779 4003 64821 4012
rect 67083 4052 67125 4061
rect 67083 4012 67084 4052
rect 67124 4012 67125 4052
rect 67083 4003 67125 4012
rect 68523 4052 68565 4061
rect 68523 4012 68524 4052
rect 68564 4012 68565 4052
rect 68523 4003 68565 4012
rect 70443 4052 70485 4061
rect 70443 4012 70444 4052
rect 70484 4012 70485 4052
rect 70443 4003 70485 4012
rect 74859 4052 74901 4061
rect 74859 4012 74860 4052
rect 74900 4012 74901 4052
rect 74859 4003 74901 4012
rect 81579 4052 81621 4061
rect 81579 4012 81580 4052
rect 81620 4012 81621 4052
rect 81579 4003 81621 4012
rect 84459 4052 84501 4061
rect 84459 4012 84460 4052
rect 84500 4012 84501 4052
rect 84459 4003 84501 4012
rect 86091 4052 86133 4061
rect 86091 4012 86092 4052
rect 86132 4012 86133 4052
rect 86091 4003 86133 4012
rect 94923 4052 94965 4061
rect 94923 4012 94924 4052
rect 94964 4012 94965 4052
rect 94923 4003 94965 4012
rect 1707 3968 1749 3977
rect 1707 3928 1708 3968
rect 1748 3928 1749 3968
rect 1707 3919 1749 3928
rect 2091 3968 2133 3977
rect 2091 3928 2092 3968
rect 2132 3928 2133 3968
rect 2091 3919 2133 3928
rect 2475 3968 2517 3977
rect 2475 3928 2476 3968
rect 2516 3928 2517 3968
rect 2475 3919 2517 3928
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 3243 3968 3285 3977
rect 3243 3928 3244 3968
rect 3284 3928 3285 3968
rect 3243 3919 3285 3928
rect 3627 3968 3669 3977
rect 3627 3928 3628 3968
rect 3668 3928 3669 3968
rect 3627 3919 3669 3928
rect 4011 3968 4053 3977
rect 4011 3928 4012 3968
rect 4052 3928 4053 3968
rect 4011 3919 4053 3928
rect 4395 3968 4437 3977
rect 4395 3928 4396 3968
rect 4436 3928 4437 3968
rect 4395 3919 4437 3928
rect 4779 3968 4821 3977
rect 4779 3928 4780 3968
rect 4820 3928 4821 3968
rect 4779 3919 4821 3928
rect 5163 3968 5205 3977
rect 5163 3928 5164 3968
rect 5204 3928 5205 3968
rect 5163 3919 5205 3928
rect 5547 3968 5589 3977
rect 5547 3928 5548 3968
rect 5588 3928 5589 3968
rect 5547 3919 5589 3928
rect 5931 3968 5973 3977
rect 5931 3928 5932 3968
rect 5972 3928 5973 3968
rect 5931 3919 5973 3928
rect 6315 3968 6357 3977
rect 6315 3928 6316 3968
rect 6356 3928 6357 3968
rect 6315 3919 6357 3928
rect 6699 3968 6741 3977
rect 6699 3928 6700 3968
rect 6740 3928 6741 3968
rect 6699 3919 6741 3928
rect 7083 3968 7125 3977
rect 7083 3928 7084 3968
rect 7124 3928 7125 3968
rect 7083 3919 7125 3928
rect 7467 3968 7509 3977
rect 7467 3928 7468 3968
rect 7508 3928 7509 3968
rect 7467 3919 7509 3928
rect 7851 3968 7893 3977
rect 7851 3928 7852 3968
rect 7892 3928 7893 3968
rect 7851 3919 7893 3928
rect 8235 3968 8277 3977
rect 8235 3928 8236 3968
rect 8276 3928 8277 3968
rect 8235 3919 8277 3928
rect 8619 3968 8661 3977
rect 8619 3928 8620 3968
rect 8660 3928 8661 3968
rect 8619 3919 8661 3928
rect 9003 3968 9045 3977
rect 9003 3928 9004 3968
rect 9044 3928 9045 3968
rect 9003 3919 9045 3928
rect 9387 3968 9429 3977
rect 9387 3928 9388 3968
rect 9428 3928 9429 3968
rect 9387 3919 9429 3928
rect 9771 3968 9813 3977
rect 9771 3928 9772 3968
rect 9812 3928 9813 3968
rect 9771 3919 9813 3928
rect 10155 3968 10197 3977
rect 10155 3928 10156 3968
rect 10196 3928 10197 3968
rect 10155 3919 10197 3928
rect 10539 3968 10581 3977
rect 10539 3928 10540 3968
rect 10580 3928 10581 3968
rect 10539 3919 10581 3928
rect 10923 3968 10965 3977
rect 10923 3928 10924 3968
rect 10964 3928 10965 3968
rect 10923 3919 10965 3928
rect 11307 3968 11349 3977
rect 11307 3928 11308 3968
rect 11348 3928 11349 3968
rect 11307 3919 11349 3928
rect 11691 3968 11733 3977
rect 11691 3928 11692 3968
rect 11732 3928 11733 3968
rect 11691 3919 11733 3928
rect 12075 3968 12117 3977
rect 12075 3928 12076 3968
rect 12116 3928 12117 3968
rect 12075 3919 12117 3928
rect 12459 3968 12501 3977
rect 12459 3928 12460 3968
rect 12500 3928 12501 3968
rect 12459 3919 12501 3928
rect 12843 3968 12885 3977
rect 12843 3928 12844 3968
rect 12884 3928 12885 3968
rect 12843 3919 12885 3928
rect 13227 3968 13269 3977
rect 13227 3928 13228 3968
rect 13268 3928 13269 3968
rect 13227 3919 13269 3928
rect 13611 3968 13653 3977
rect 13611 3928 13612 3968
rect 13652 3928 13653 3968
rect 13611 3919 13653 3928
rect 13995 3968 14037 3977
rect 13995 3928 13996 3968
rect 14036 3928 14037 3968
rect 13995 3919 14037 3928
rect 14379 3968 14421 3977
rect 14379 3928 14380 3968
rect 14420 3928 14421 3968
rect 14379 3919 14421 3928
rect 14763 3968 14805 3977
rect 14763 3928 14764 3968
rect 14804 3928 14805 3968
rect 14763 3919 14805 3928
rect 15147 3968 15189 3977
rect 15147 3928 15148 3968
rect 15188 3928 15189 3968
rect 15147 3919 15189 3928
rect 15531 3968 15573 3977
rect 15531 3928 15532 3968
rect 15572 3928 15573 3968
rect 15531 3919 15573 3928
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 16299 3968 16341 3977
rect 16299 3928 16300 3968
rect 16340 3928 16341 3968
rect 16299 3919 16341 3928
rect 16683 3968 16725 3977
rect 16683 3928 16684 3968
rect 16724 3928 16725 3968
rect 16683 3919 16725 3928
rect 17355 3968 17397 3977
rect 17355 3928 17356 3968
rect 17396 3928 17397 3968
rect 17355 3919 17397 3928
rect 17931 3968 17973 3977
rect 17931 3928 17932 3968
rect 17972 3928 17973 3968
rect 17931 3919 17973 3928
rect 18315 3968 18357 3977
rect 18315 3928 18316 3968
rect 18356 3928 18357 3968
rect 18315 3919 18357 3928
rect 18699 3968 18741 3977
rect 18699 3928 18700 3968
rect 18740 3928 18741 3968
rect 18699 3919 18741 3928
rect 19755 3968 19797 3977
rect 19755 3928 19756 3968
rect 19796 3928 19797 3968
rect 19755 3919 19797 3928
rect 19947 3968 19989 3977
rect 19947 3928 19948 3968
rect 19988 3928 19989 3968
rect 19947 3919 19989 3928
rect 20523 3968 20565 3977
rect 20523 3928 20524 3968
rect 20564 3928 20565 3968
rect 20523 3919 20565 3928
rect 20907 3968 20949 3977
rect 20907 3928 20908 3968
rect 20948 3928 20949 3968
rect 20907 3919 20949 3928
rect 21483 3968 21525 3977
rect 21483 3928 21484 3968
rect 21524 3928 21525 3968
rect 21483 3919 21525 3928
rect 21867 3968 21909 3977
rect 21867 3928 21868 3968
rect 21908 3928 21909 3968
rect 21867 3919 21909 3928
rect 23211 3968 23253 3977
rect 23211 3928 23212 3968
rect 23252 3928 23253 3968
rect 23211 3919 23253 3928
rect 23595 3968 23637 3977
rect 23595 3928 23596 3968
rect 23636 3928 23637 3968
rect 23595 3919 23637 3928
rect 24555 3968 24597 3977
rect 24555 3928 24556 3968
rect 24596 3928 24597 3968
rect 24555 3919 24597 3928
rect 25515 3968 25557 3977
rect 25515 3928 25516 3968
rect 25556 3928 25557 3968
rect 25515 3919 25557 3928
rect 25899 3968 25941 3977
rect 25899 3928 25900 3968
rect 25940 3928 25941 3968
rect 25899 3919 25941 3928
rect 26283 3968 26325 3977
rect 26283 3928 26284 3968
rect 26324 3928 26325 3968
rect 26283 3919 26325 3928
rect 26667 3968 26709 3977
rect 26667 3928 26668 3968
rect 26708 3928 26709 3968
rect 26667 3919 26709 3928
rect 27051 3968 27093 3977
rect 27051 3928 27052 3968
rect 27092 3928 27093 3968
rect 27051 3919 27093 3928
rect 27435 3968 27477 3977
rect 27435 3928 27436 3968
rect 27476 3928 27477 3968
rect 27435 3919 27477 3928
rect 27627 3968 27669 3977
rect 27627 3928 27628 3968
rect 27668 3928 27669 3968
rect 27627 3919 27669 3928
rect 28587 3968 28629 3977
rect 28587 3928 28588 3968
rect 28628 3928 28629 3968
rect 28587 3919 28629 3928
rect 28971 3968 29013 3977
rect 28971 3928 28972 3968
rect 29012 3928 29013 3968
rect 28971 3919 29013 3928
rect 30123 3968 30165 3977
rect 30123 3928 30124 3968
rect 30164 3928 30165 3968
rect 30123 3919 30165 3928
rect 30315 3968 30357 3977
rect 30315 3928 30316 3968
rect 30356 3928 30357 3968
rect 30315 3919 30357 3928
rect 31659 3968 31701 3977
rect 31659 3928 31660 3968
rect 31700 3928 31701 3968
rect 31659 3919 31701 3928
rect 32043 3968 32085 3977
rect 32043 3928 32044 3968
rect 32084 3928 32085 3968
rect 32043 3919 32085 3928
rect 32427 3968 32469 3977
rect 32427 3928 32428 3968
rect 32468 3928 32469 3968
rect 32427 3919 32469 3928
rect 32811 3968 32853 3977
rect 32811 3928 32812 3968
rect 32852 3928 32853 3968
rect 32811 3919 32853 3928
rect 33195 3968 33237 3977
rect 33195 3928 33196 3968
rect 33236 3928 33237 3968
rect 33195 3919 33237 3928
rect 33579 3968 33621 3977
rect 33579 3928 33580 3968
rect 33620 3928 33621 3968
rect 33579 3919 33621 3928
rect 36267 3968 36309 3977
rect 36267 3928 36268 3968
rect 36308 3928 36309 3968
rect 36267 3919 36309 3928
rect 36651 3968 36693 3977
rect 36651 3928 36652 3968
rect 36692 3928 36693 3968
rect 36651 3919 36693 3928
rect 37035 3968 37077 3977
rect 37035 3928 37036 3968
rect 37076 3928 37077 3968
rect 37035 3919 37077 3928
rect 37419 3968 37461 3977
rect 37419 3928 37420 3968
rect 37460 3928 37461 3968
rect 37419 3919 37461 3928
rect 37803 3968 37845 3977
rect 37803 3928 37804 3968
rect 37844 3928 37845 3968
rect 37803 3919 37845 3928
rect 38187 3968 38229 3977
rect 38187 3928 38188 3968
rect 38228 3928 38229 3968
rect 38187 3919 38229 3928
rect 38955 3968 38997 3977
rect 38955 3928 38956 3968
rect 38996 3928 38997 3968
rect 38955 3919 38997 3928
rect 39339 3968 39381 3977
rect 39339 3928 39340 3968
rect 39380 3928 39381 3968
rect 39339 3919 39381 3928
rect 39723 3968 39765 3977
rect 39723 3928 39724 3968
rect 39764 3928 39765 3968
rect 39723 3919 39765 3928
rect 40107 3968 40149 3977
rect 40107 3928 40108 3968
rect 40148 3928 40149 3968
rect 40107 3919 40149 3928
rect 40491 3968 40533 3977
rect 40491 3928 40492 3968
rect 40532 3928 40533 3968
rect 40491 3919 40533 3928
rect 40875 3968 40917 3977
rect 40875 3928 40876 3968
rect 40916 3928 40917 3968
rect 40875 3919 40917 3928
rect 41259 3968 41301 3977
rect 41259 3928 41260 3968
rect 41300 3928 41301 3968
rect 41259 3919 41301 3928
rect 41643 3968 41685 3977
rect 41643 3928 41644 3968
rect 41684 3928 41685 3968
rect 41643 3919 41685 3928
rect 42027 3968 42069 3977
rect 42027 3928 42028 3968
rect 42068 3928 42069 3968
rect 42027 3919 42069 3928
rect 42411 3968 42453 3977
rect 42411 3928 42412 3968
rect 42452 3928 42453 3968
rect 42411 3919 42453 3928
rect 43179 3968 43221 3977
rect 43179 3928 43180 3968
rect 43220 3928 43221 3968
rect 43179 3919 43221 3928
rect 43563 3968 43605 3977
rect 43563 3928 43564 3968
rect 43604 3928 43605 3968
rect 43563 3919 43605 3928
rect 44235 3968 44277 3977
rect 44235 3928 44236 3968
rect 44276 3928 44277 3968
rect 44235 3919 44277 3928
rect 46731 3968 46773 3977
rect 46731 3928 46732 3968
rect 46772 3928 46773 3968
rect 46731 3919 46773 3928
rect 49227 3968 49269 3977
rect 49227 3928 49228 3968
rect 49268 3928 49269 3968
rect 49227 3919 49269 3928
rect 49707 3968 49749 3977
rect 49707 3928 49708 3968
rect 49748 3928 49749 3968
rect 49707 3919 49749 3928
rect 50667 3968 50709 3977
rect 50667 3928 50668 3968
rect 50708 3928 50709 3968
rect 50667 3919 50709 3928
rect 51051 3968 51093 3977
rect 51051 3928 51052 3968
rect 51092 3928 51093 3968
rect 51051 3919 51093 3928
rect 52395 3968 52437 3977
rect 52395 3928 52396 3968
rect 52436 3928 52437 3968
rect 52395 3919 52437 3928
rect 53355 3968 53397 3977
rect 53355 3928 53356 3968
rect 53396 3928 53397 3968
rect 53355 3919 53397 3928
rect 53739 3968 53781 3977
rect 53739 3928 53740 3968
rect 53780 3928 53781 3968
rect 53739 3919 53781 3928
rect 54123 3968 54165 3977
rect 54123 3928 54124 3968
rect 54164 3928 54165 3968
rect 54123 3919 54165 3928
rect 55467 3968 55509 3977
rect 55467 3928 55468 3968
rect 55508 3928 55509 3968
rect 55467 3919 55509 3928
rect 55851 3968 55893 3977
rect 55851 3928 55852 3968
rect 55892 3928 55893 3968
rect 55851 3919 55893 3928
rect 57195 3968 57237 3977
rect 57195 3928 57196 3968
rect 57236 3928 57237 3968
rect 57195 3919 57237 3928
rect 57387 3968 57429 3977
rect 57387 3928 57388 3968
rect 57428 3928 57429 3968
rect 57387 3919 57429 3928
rect 61419 3968 61461 3977
rect 61419 3928 61420 3968
rect 61460 3928 61461 3968
rect 61419 3919 61461 3928
rect 61803 3968 61845 3977
rect 61803 3928 61804 3968
rect 61844 3928 61845 3968
rect 61803 3919 61845 3928
rect 62187 3968 62229 3977
rect 62187 3928 62188 3968
rect 62228 3928 62229 3968
rect 62187 3919 62229 3928
rect 62571 3968 62613 3977
rect 62571 3928 62572 3968
rect 62612 3928 62613 3968
rect 62571 3919 62613 3928
rect 65067 3968 65109 3977
rect 65067 3928 65068 3968
rect 65108 3928 65109 3968
rect 65067 3919 65109 3928
rect 65451 3968 65493 3977
rect 65451 3928 65452 3968
rect 65492 3928 65493 3968
rect 65451 3919 65493 3928
rect 65835 3968 65877 3977
rect 65835 3928 65836 3968
rect 65876 3928 65877 3968
rect 65835 3919 65877 3928
rect 66219 3968 66261 3977
rect 66219 3928 66220 3968
rect 66260 3928 66261 3968
rect 66219 3919 66261 3928
rect 67371 3968 67413 3977
rect 67371 3928 67372 3968
rect 67412 3928 67413 3968
rect 67371 3919 67413 3928
rect 67755 3968 67797 3977
rect 67755 3928 67756 3968
rect 67796 3928 67797 3968
rect 67755 3919 67797 3928
rect 68139 3968 68181 3977
rect 68139 3928 68140 3968
rect 68180 3928 68181 3968
rect 68139 3919 68181 3928
rect 69291 3968 69333 3977
rect 69291 3928 69292 3968
rect 69332 3928 69333 3968
rect 69291 3919 69333 3928
rect 69675 3968 69717 3977
rect 69675 3928 69676 3968
rect 69716 3928 69717 3968
rect 69675 3919 69717 3928
rect 70251 3968 70293 3977
rect 70251 3928 70252 3968
rect 70292 3928 70293 3968
rect 70251 3919 70293 3928
rect 71787 3968 71829 3977
rect 71787 3928 71788 3968
rect 71828 3928 71829 3968
rect 71787 3919 71829 3928
rect 72171 3968 72213 3977
rect 72171 3928 72172 3968
rect 72212 3928 72213 3968
rect 72171 3919 72213 3928
rect 72363 3968 72405 3977
rect 72363 3928 72364 3968
rect 72404 3928 72405 3968
rect 72363 3919 72405 3928
rect 73323 3968 73365 3977
rect 73323 3928 73324 3968
rect 73364 3928 73365 3968
rect 73323 3919 73365 3928
rect 73707 3968 73749 3977
rect 73707 3928 73708 3968
rect 73748 3928 73749 3968
rect 73707 3919 73749 3928
rect 73899 3968 73941 3977
rect 73899 3928 73900 3968
rect 73940 3928 73941 3968
rect 73899 3919 73941 3928
rect 74283 3968 74325 3977
rect 74283 3928 74284 3968
rect 74324 3928 74325 3968
rect 74283 3919 74325 3928
rect 75051 3968 75093 3977
rect 75051 3928 75052 3968
rect 75092 3928 75093 3968
rect 75051 3919 75093 3928
rect 75435 3968 75477 3977
rect 75435 3928 75436 3968
rect 75476 3928 75477 3968
rect 75435 3919 75477 3928
rect 76011 3968 76053 3977
rect 76011 3928 76012 3968
rect 76052 3928 76053 3968
rect 76011 3919 76053 3928
rect 76203 3968 76245 3977
rect 76203 3928 76204 3968
rect 76244 3928 76245 3968
rect 76203 3919 76245 3928
rect 76779 3968 76821 3977
rect 76779 3928 76780 3968
rect 76820 3928 76821 3968
rect 76779 3919 76821 3928
rect 78795 3968 78837 3977
rect 78795 3928 78796 3968
rect 78836 3928 78837 3968
rect 78795 3919 78837 3928
rect 79179 3968 79221 3977
rect 79179 3928 79180 3968
rect 79220 3928 79221 3968
rect 79179 3919 79221 3928
rect 79563 3968 79605 3977
rect 79563 3928 79564 3968
rect 79604 3928 79605 3968
rect 79563 3919 79605 3928
rect 79947 3968 79989 3977
rect 79947 3928 79948 3968
rect 79988 3928 79989 3968
rect 79947 3919 79989 3928
rect 80331 3968 80373 3977
rect 80331 3928 80332 3968
rect 80372 3928 80373 3968
rect 80331 3919 80373 3928
rect 80907 3968 80949 3977
rect 80907 3928 80908 3968
rect 80948 3928 80949 3968
rect 80907 3919 80949 3928
rect 82443 3968 82485 3977
rect 82443 3928 82444 3968
rect 82484 3928 82485 3968
rect 82443 3919 82485 3928
rect 82827 3968 82869 3977
rect 82827 3928 82828 3968
rect 82868 3928 82869 3968
rect 82827 3919 82869 3928
rect 83403 3968 83445 3977
rect 83403 3928 83404 3968
rect 83444 3928 83445 3968
rect 83403 3919 83445 3928
rect 83595 3968 83637 3977
rect 83595 3928 83596 3968
rect 83636 3928 83637 3968
rect 83595 3919 83637 3928
rect 85707 3968 85749 3977
rect 85707 3928 85708 3968
rect 85748 3928 85749 3968
rect 85707 3919 85749 3928
rect 86475 3968 86517 3977
rect 86475 3928 86476 3968
rect 86516 3928 86517 3968
rect 86475 3919 86517 3928
rect 86859 3968 86901 3977
rect 86859 3928 86860 3968
rect 86900 3928 86901 3968
rect 86859 3919 86901 3928
rect 87243 3968 87285 3977
rect 87243 3928 87244 3968
rect 87284 3928 87285 3968
rect 87243 3919 87285 3928
rect 87627 3968 87669 3977
rect 87627 3928 87628 3968
rect 87668 3928 87669 3968
rect 87627 3919 87669 3928
rect 88011 3968 88053 3977
rect 88011 3928 88012 3968
rect 88052 3928 88053 3968
rect 88011 3919 88053 3928
rect 88395 3968 88437 3977
rect 88395 3928 88396 3968
rect 88436 3928 88437 3968
rect 88395 3919 88437 3928
rect 88779 3968 88821 3977
rect 88779 3928 88780 3968
rect 88820 3928 88821 3968
rect 88779 3919 88821 3928
rect 89163 3968 89205 3977
rect 89163 3928 89164 3968
rect 89204 3928 89205 3968
rect 89163 3919 89205 3928
rect 89547 3968 89589 3977
rect 89547 3928 89548 3968
rect 89588 3928 89589 3968
rect 89547 3919 89589 3928
rect 89931 3968 89973 3977
rect 89931 3928 89932 3968
rect 89972 3928 89973 3968
rect 89931 3919 89973 3928
rect 90315 3968 90357 3977
rect 90315 3928 90316 3968
rect 90356 3928 90357 3968
rect 90315 3919 90357 3928
rect 90699 3968 90741 3977
rect 90699 3928 90700 3968
rect 90740 3928 90741 3968
rect 90699 3919 90741 3928
rect 91083 3968 91125 3977
rect 91083 3928 91084 3968
rect 91124 3928 91125 3968
rect 91083 3919 91125 3928
rect 91467 3968 91509 3977
rect 91467 3928 91468 3968
rect 91508 3928 91509 3968
rect 91467 3919 91509 3928
rect 91851 3968 91893 3977
rect 91851 3928 91852 3968
rect 91892 3928 91893 3968
rect 91851 3919 91893 3928
rect 92235 3968 92277 3977
rect 92235 3928 92236 3968
rect 92276 3928 92277 3968
rect 92235 3919 92277 3928
rect 92619 3968 92661 3977
rect 92619 3928 92620 3968
rect 92660 3928 92661 3968
rect 92619 3919 92661 3928
rect 93003 3968 93045 3977
rect 93003 3928 93004 3968
rect 93044 3928 93045 3968
rect 93003 3919 93045 3928
rect 93387 3968 93429 3977
rect 93387 3928 93388 3968
rect 93428 3928 93429 3968
rect 93387 3919 93429 3928
rect 93771 3968 93813 3977
rect 93771 3928 93772 3968
rect 93812 3928 93813 3968
rect 93771 3919 93813 3928
rect 94155 3968 94197 3977
rect 94155 3928 94156 3968
rect 94196 3928 94197 3968
rect 94155 3919 94197 3928
rect 94539 3968 94581 3977
rect 94539 3928 94540 3968
rect 94580 3928 94581 3968
rect 94539 3919 94581 3928
rect 95307 3968 95349 3977
rect 95307 3928 95308 3968
rect 95348 3928 95349 3968
rect 95307 3919 95349 3928
rect 95691 3968 95733 3977
rect 95691 3928 95692 3968
rect 95732 3928 95733 3968
rect 95691 3919 95733 3928
rect 96075 3968 96117 3977
rect 96075 3928 96076 3968
rect 96116 3928 96117 3968
rect 96075 3919 96117 3928
rect 96459 3968 96501 3977
rect 96459 3928 96460 3968
rect 96500 3928 96501 3968
rect 96459 3919 96501 3928
rect 96843 3968 96885 3977
rect 96843 3928 96844 3968
rect 96884 3928 96885 3968
rect 96843 3919 96885 3928
rect 97227 3968 97269 3977
rect 97227 3928 97228 3968
rect 97268 3928 97269 3968
rect 97227 3919 97269 3928
rect 97611 3968 97653 3977
rect 97611 3928 97612 3968
rect 97652 3928 97653 3968
rect 97611 3919 97653 3928
rect 97995 3968 98037 3977
rect 97995 3928 97996 3968
rect 98036 3928 98037 3968
rect 97995 3919 98037 3928
rect 98379 3968 98421 3977
rect 98379 3928 98380 3968
rect 98420 3928 98421 3968
rect 98379 3919 98421 3928
rect 1152 3800 98784 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 64168 3800
rect 64208 3760 64250 3800
rect 64290 3760 64332 3800
rect 64372 3760 64414 3800
rect 64454 3760 64496 3800
rect 64536 3760 79288 3800
rect 79328 3760 79370 3800
rect 79410 3760 79452 3800
rect 79492 3760 79534 3800
rect 79574 3760 79616 3800
rect 79656 3760 94408 3800
rect 94448 3760 94490 3800
rect 94530 3760 94572 3800
rect 94612 3760 94654 3800
rect 94694 3760 94736 3800
rect 94776 3760 98784 3800
rect 1152 3736 98784 3760
rect 49803 3632 49845 3641
rect 49803 3592 49804 3632
rect 49844 3592 49845 3632
rect 49803 3583 49845 3592
rect 65355 3632 65397 3641
rect 65355 3592 65356 3632
rect 65396 3592 65397 3632
rect 65355 3583 65397 3592
rect 81771 3632 81813 3641
rect 81771 3592 81772 3632
rect 81812 3592 81813 3632
rect 81771 3583 81813 3592
rect 85131 3632 85173 3641
rect 85131 3592 85132 3632
rect 85172 3592 85173 3632
rect 85131 3583 85173 3592
rect 49611 3548 49653 3557
rect 49611 3508 49612 3548
rect 49652 3508 49653 3548
rect 49611 3499 49653 3508
rect 50091 3548 50133 3557
rect 50091 3508 50092 3548
rect 50132 3508 50133 3548
rect 50091 3499 50133 3508
rect 50283 3548 50325 3557
rect 50283 3508 50284 3548
rect 50324 3508 50325 3548
rect 50283 3499 50325 3508
rect 52491 3548 52533 3557
rect 52491 3508 52492 3548
rect 52532 3508 52533 3548
rect 52491 3499 52533 3508
rect 52683 3548 52725 3557
rect 52683 3508 52684 3548
rect 52724 3508 52725 3548
rect 52683 3499 52725 3508
rect 54795 3548 54837 3557
rect 54795 3508 54796 3548
rect 54836 3508 54837 3548
rect 54795 3499 54837 3508
rect 57291 3548 57333 3557
rect 57291 3508 57292 3548
rect 57332 3508 57333 3548
rect 57291 3499 57333 3508
rect 60267 3548 60309 3557
rect 60267 3508 60268 3548
rect 60308 3508 60309 3548
rect 60267 3499 60309 3508
rect 64971 3548 65013 3557
rect 64971 3508 64972 3548
rect 65012 3508 65013 3548
rect 64971 3499 65013 3508
rect 82635 3548 82677 3557
rect 82635 3508 82636 3548
rect 82676 3508 82677 3548
rect 82635 3499 82677 3508
rect 75907 3475 75965 3476
rect 1219 3464 1277 3465
rect 1219 3424 1228 3464
rect 1268 3424 1277 3464
rect 1219 3423 1277 3424
rect 1603 3464 1661 3465
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 1603 3423 1661 3424
rect 1987 3464 2045 3465
rect 1987 3424 1996 3464
rect 2036 3424 2045 3464
rect 1987 3423 2045 3424
rect 2371 3464 2429 3465
rect 2371 3424 2380 3464
rect 2420 3424 2429 3464
rect 2371 3423 2429 3424
rect 2755 3464 2813 3465
rect 2755 3424 2764 3464
rect 2804 3424 2813 3464
rect 2755 3423 2813 3424
rect 3139 3464 3197 3465
rect 3139 3424 3148 3464
rect 3188 3424 3197 3464
rect 3139 3423 3197 3424
rect 3523 3464 3581 3465
rect 3523 3424 3532 3464
rect 3572 3424 3581 3464
rect 3523 3423 3581 3424
rect 3907 3464 3965 3465
rect 3907 3424 3916 3464
rect 3956 3424 3965 3464
rect 3907 3423 3965 3424
rect 4291 3464 4349 3465
rect 4291 3424 4300 3464
rect 4340 3424 4349 3464
rect 4291 3423 4349 3424
rect 4675 3464 4733 3465
rect 4675 3424 4684 3464
rect 4724 3424 4733 3464
rect 4675 3423 4733 3424
rect 5059 3464 5117 3465
rect 5059 3424 5068 3464
rect 5108 3424 5117 3464
rect 5059 3423 5117 3424
rect 5443 3464 5501 3465
rect 5443 3424 5452 3464
rect 5492 3424 5501 3464
rect 5443 3423 5501 3424
rect 5827 3464 5885 3465
rect 5827 3424 5836 3464
rect 5876 3424 5885 3464
rect 5827 3423 5885 3424
rect 6211 3464 6269 3465
rect 6211 3424 6220 3464
rect 6260 3424 6269 3464
rect 6211 3423 6269 3424
rect 6595 3464 6653 3465
rect 6595 3424 6604 3464
rect 6644 3424 6653 3464
rect 6595 3423 6653 3424
rect 6979 3464 7037 3465
rect 6979 3424 6988 3464
rect 7028 3424 7037 3464
rect 6979 3423 7037 3424
rect 7363 3464 7421 3465
rect 7363 3424 7372 3464
rect 7412 3424 7421 3464
rect 7363 3423 7421 3424
rect 7747 3464 7805 3465
rect 7747 3424 7756 3464
rect 7796 3424 7805 3464
rect 7747 3423 7805 3424
rect 8131 3464 8189 3465
rect 8131 3424 8140 3464
rect 8180 3424 8189 3464
rect 8131 3423 8189 3424
rect 8515 3464 8573 3465
rect 8515 3424 8524 3464
rect 8564 3424 8573 3464
rect 8515 3423 8573 3424
rect 8899 3464 8957 3465
rect 8899 3424 8908 3464
rect 8948 3424 8957 3464
rect 8899 3423 8957 3424
rect 9283 3464 9341 3465
rect 9283 3424 9292 3464
rect 9332 3424 9341 3464
rect 9283 3423 9341 3424
rect 9667 3464 9725 3465
rect 9667 3424 9676 3464
rect 9716 3424 9725 3464
rect 9667 3423 9725 3424
rect 10051 3464 10109 3465
rect 10051 3424 10060 3464
rect 10100 3424 10109 3464
rect 10051 3423 10109 3424
rect 10435 3464 10493 3465
rect 10435 3424 10444 3464
rect 10484 3424 10493 3464
rect 10435 3423 10493 3424
rect 10819 3464 10877 3465
rect 10819 3424 10828 3464
rect 10868 3424 10877 3464
rect 10819 3423 10877 3424
rect 11203 3464 11261 3465
rect 11203 3424 11212 3464
rect 11252 3424 11261 3464
rect 11203 3423 11261 3424
rect 11587 3464 11645 3465
rect 11587 3424 11596 3464
rect 11636 3424 11645 3464
rect 11587 3423 11645 3424
rect 11971 3464 12029 3465
rect 11971 3424 11980 3464
rect 12020 3424 12029 3464
rect 11971 3423 12029 3424
rect 12355 3464 12413 3465
rect 12355 3424 12364 3464
rect 12404 3424 12413 3464
rect 12355 3423 12413 3424
rect 12739 3464 12797 3465
rect 12739 3424 12748 3464
rect 12788 3424 12797 3464
rect 12739 3423 12797 3424
rect 13123 3464 13181 3465
rect 13123 3424 13132 3464
rect 13172 3424 13181 3464
rect 13123 3423 13181 3424
rect 13507 3464 13565 3465
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13507 3423 13565 3424
rect 13891 3464 13949 3465
rect 13891 3424 13900 3464
rect 13940 3424 13949 3464
rect 13891 3423 13949 3424
rect 14275 3464 14333 3465
rect 14275 3424 14284 3464
rect 14324 3424 14333 3464
rect 14275 3423 14333 3424
rect 14659 3464 14717 3465
rect 14659 3424 14668 3464
rect 14708 3424 14717 3464
rect 14659 3423 14717 3424
rect 15043 3464 15101 3465
rect 15043 3424 15052 3464
rect 15092 3424 15101 3464
rect 15043 3423 15101 3424
rect 15427 3464 15485 3465
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 15811 3464 15869 3465
rect 15811 3424 15820 3464
rect 15860 3424 15869 3464
rect 15811 3423 15869 3424
rect 16195 3464 16253 3465
rect 16195 3424 16204 3464
rect 16244 3424 16253 3464
rect 16195 3423 16253 3424
rect 16579 3464 16637 3465
rect 16579 3424 16588 3464
rect 16628 3424 16637 3464
rect 16579 3423 16637 3424
rect 16963 3464 17021 3465
rect 16963 3424 16972 3464
rect 17012 3424 17021 3464
rect 16963 3423 17021 3424
rect 17347 3464 17405 3465
rect 17347 3424 17356 3464
rect 17396 3424 17405 3464
rect 17347 3423 17405 3424
rect 18499 3464 18557 3465
rect 18499 3424 18508 3464
rect 18548 3424 18557 3464
rect 18499 3423 18557 3424
rect 18883 3464 18941 3465
rect 18883 3424 18892 3464
rect 18932 3424 18941 3464
rect 18883 3423 18941 3424
rect 19267 3464 19325 3465
rect 19267 3424 19276 3464
rect 19316 3424 19325 3464
rect 19267 3423 19325 3424
rect 19651 3464 19709 3465
rect 19651 3424 19660 3464
rect 19700 3424 19709 3464
rect 19651 3423 19709 3424
rect 20035 3464 20093 3465
rect 20035 3424 20044 3464
rect 20084 3424 20093 3464
rect 20035 3423 20093 3424
rect 20419 3464 20477 3465
rect 20419 3424 20428 3464
rect 20468 3424 20477 3464
rect 20419 3423 20477 3424
rect 20803 3464 20861 3465
rect 20803 3424 20812 3464
rect 20852 3424 20861 3464
rect 20803 3423 20861 3424
rect 21187 3464 21245 3465
rect 21187 3424 21196 3464
rect 21236 3424 21245 3464
rect 21187 3423 21245 3424
rect 21571 3464 21629 3465
rect 21571 3424 21580 3464
rect 21620 3424 21629 3464
rect 21571 3423 21629 3424
rect 21955 3464 22013 3465
rect 21955 3424 21964 3464
rect 22004 3424 22013 3464
rect 21955 3423 22013 3424
rect 22339 3464 22397 3465
rect 22339 3424 22348 3464
rect 22388 3424 22397 3464
rect 22339 3423 22397 3424
rect 22723 3464 22781 3465
rect 22723 3424 22732 3464
rect 22772 3424 22781 3464
rect 22723 3423 22781 3424
rect 23107 3464 23165 3465
rect 23107 3424 23116 3464
rect 23156 3424 23165 3464
rect 23107 3423 23165 3424
rect 23491 3464 23549 3465
rect 23491 3424 23500 3464
rect 23540 3424 23549 3464
rect 23491 3423 23549 3424
rect 23875 3464 23933 3465
rect 23875 3424 23884 3464
rect 23924 3424 23933 3464
rect 23875 3423 23933 3424
rect 24259 3464 24317 3465
rect 24259 3424 24268 3464
rect 24308 3424 24317 3464
rect 24259 3423 24317 3424
rect 24643 3464 24701 3465
rect 24643 3424 24652 3464
rect 24692 3424 24701 3464
rect 24643 3423 24701 3424
rect 25027 3464 25085 3465
rect 25027 3424 25036 3464
rect 25076 3424 25085 3464
rect 25027 3423 25085 3424
rect 25411 3464 25469 3465
rect 25411 3424 25420 3464
rect 25460 3424 25469 3464
rect 25411 3423 25469 3424
rect 25795 3464 25853 3465
rect 25795 3424 25804 3464
rect 25844 3424 25853 3464
rect 25795 3423 25853 3424
rect 26179 3464 26237 3465
rect 26179 3424 26188 3464
rect 26228 3424 26237 3464
rect 26179 3423 26237 3424
rect 26563 3464 26621 3465
rect 26563 3424 26572 3464
rect 26612 3424 26621 3464
rect 26563 3423 26621 3424
rect 26947 3464 27005 3465
rect 26947 3424 26956 3464
rect 26996 3424 27005 3464
rect 26947 3423 27005 3424
rect 27331 3464 27389 3465
rect 27331 3424 27340 3464
rect 27380 3424 27389 3464
rect 27331 3423 27389 3424
rect 27715 3464 27773 3465
rect 27715 3424 27724 3464
rect 27764 3424 27773 3464
rect 27715 3423 27773 3424
rect 28099 3464 28157 3465
rect 28099 3424 28108 3464
rect 28148 3424 28157 3464
rect 28099 3423 28157 3424
rect 28483 3464 28541 3465
rect 28483 3424 28492 3464
rect 28532 3424 28541 3464
rect 28483 3423 28541 3424
rect 28867 3464 28925 3465
rect 28867 3424 28876 3464
rect 28916 3424 28925 3464
rect 28867 3423 28925 3424
rect 29251 3464 29309 3465
rect 29251 3424 29260 3464
rect 29300 3424 29309 3464
rect 29251 3423 29309 3424
rect 29635 3464 29693 3465
rect 29635 3424 29644 3464
rect 29684 3424 29693 3464
rect 29635 3423 29693 3424
rect 30019 3464 30077 3465
rect 30019 3424 30028 3464
rect 30068 3424 30077 3464
rect 30019 3423 30077 3424
rect 30403 3464 30461 3465
rect 30403 3424 30412 3464
rect 30452 3424 30461 3464
rect 30403 3423 30461 3424
rect 30787 3464 30845 3465
rect 30787 3424 30796 3464
rect 30836 3424 30845 3464
rect 30787 3423 30845 3424
rect 31171 3464 31229 3465
rect 31171 3424 31180 3464
rect 31220 3424 31229 3464
rect 31171 3423 31229 3424
rect 31555 3464 31613 3465
rect 31555 3424 31564 3464
rect 31604 3424 31613 3464
rect 31555 3423 31613 3424
rect 31939 3464 31997 3465
rect 31939 3424 31948 3464
rect 31988 3424 31997 3464
rect 31939 3423 31997 3424
rect 32323 3464 32381 3465
rect 32323 3424 32332 3464
rect 32372 3424 32381 3464
rect 32323 3423 32381 3424
rect 32707 3464 32765 3465
rect 32707 3424 32716 3464
rect 32756 3424 32765 3464
rect 32707 3423 32765 3424
rect 33091 3464 33149 3465
rect 33091 3424 33100 3464
rect 33140 3424 33149 3464
rect 33091 3423 33149 3424
rect 33475 3464 33533 3465
rect 33475 3424 33484 3464
rect 33524 3424 33533 3464
rect 33475 3423 33533 3424
rect 33859 3464 33917 3465
rect 33859 3424 33868 3464
rect 33908 3424 33917 3464
rect 33859 3423 33917 3424
rect 34243 3464 34301 3465
rect 34243 3424 34252 3464
rect 34292 3424 34301 3464
rect 34243 3423 34301 3424
rect 35299 3464 35357 3465
rect 35299 3424 35308 3464
rect 35348 3424 35357 3464
rect 35299 3423 35357 3424
rect 35683 3464 35741 3465
rect 35683 3424 35692 3464
rect 35732 3424 35741 3464
rect 35683 3423 35741 3424
rect 36067 3464 36125 3465
rect 36067 3424 36076 3464
rect 36116 3424 36125 3464
rect 36067 3423 36125 3424
rect 36451 3464 36509 3465
rect 36451 3424 36460 3464
rect 36500 3424 36509 3464
rect 36451 3423 36509 3424
rect 36835 3464 36893 3465
rect 36835 3424 36844 3464
rect 36884 3424 36893 3464
rect 36835 3423 36893 3424
rect 37219 3464 37277 3465
rect 37219 3424 37228 3464
rect 37268 3424 37277 3464
rect 37219 3423 37277 3424
rect 37603 3464 37661 3465
rect 37603 3424 37612 3464
rect 37652 3424 37661 3464
rect 37603 3423 37661 3424
rect 37987 3464 38045 3465
rect 37987 3424 37996 3464
rect 38036 3424 38045 3464
rect 37987 3423 38045 3424
rect 38371 3464 38429 3465
rect 38371 3424 38380 3464
rect 38420 3424 38429 3464
rect 38371 3423 38429 3424
rect 38755 3464 38813 3465
rect 38755 3424 38764 3464
rect 38804 3424 38813 3464
rect 38755 3423 38813 3424
rect 39139 3464 39197 3465
rect 39139 3424 39148 3464
rect 39188 3424 39197 3464
rect 39139 3423 39197 3424
rect 39523 3464 39581 3465
rect 39523 3424 39532 3464
rect 39572 3424 39581 3464
rect 39523 3423 39581 3424
rect 39907 3464 39965 3465
rect 39907 3424 39916 3464
rect 39956 3424 39965 3464
rect 39907 3423 39965 3424
rect 40291 3464 40349 3465
rect 40291 3424 40300 3464
rect 40340 3424 40349 3464
rect 40291 3423 40349 3424
rect 40675 3464 40733 3465
rect 40675 3424 40684 3464
rect 40724 3424 40733 3464
rect 40675 3423 40733 3424
rect 41059 3464 41117 3465
rect 41059 3424 41068 3464
rect 41108 3424 41117 3464
rect 41059 3423 41117 3424
rect 41443 3464 41501 3465
rect 41443 3424 41452 3464
rect 41492 3424 41501 3464
rect 41443 3423 41501 3424
rect 41827 3464 41885 3465
rect 41827 3424 41836 3464
rect 41876 3424 41885 3464
rect 41827 3423 41885 3424
rect 42211 3464 42269 3465
rect 42211 3424 42220 3464
rect 42260 3424 42269 3464
rect 42211 3423 42269 3424
rect 42595 3464 42653 3465
rect 42595 3424 42604 3464
rect 42644 3424 42653 3464
rect 42595 3423 42653 3424
rect 42979 3464 43037 3465
rect 42979 3424 42988 3464
rect 43028 3424 43037 3464
rect 42979 3423 43037 3424
rect 43363 3464 43421 3465
rect 43363 3424 43372 3464
rect 43412 3424 43421 3464
rect 43363 3423 43421 3424
rect 43747 3464 43805 3465
rect 43747 3424 43756 3464
rect 43796 3424 43805 3464
rect 43747 3423 43805 3424
rect 44131 3464 44189 3465
rect 44131 3424 44140 3464
rect 44180 3424 44189 3464
rect 44131 3423 44189 3424
rect 44515 3464 44573 3465
rect 44515 3424 44524 3464
rect 44564 3424 44573 3464
rect 44515 3423 44573 3424
rect 44899 3464 44957 3465
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 44899 3423 44957 3424
rect 45283 3464 45341 3465
rect 45283 3424 45292 3464
rect 45332 3424 45341 3464
rect 45283 3423 45341 3424
rect 45667 3464 45725 3465
rect 45667 3424 45676 3464
rect 45716 3424 45725 3464
rect 45667 3423 45725 3424
rect 47971 3464 48029 3465
rect 47971 3424 47980 3464
rect 48020 3424 48029 3464
rect 47971 3423 48029 3424
rect 48355 3464 48413 3465
rect 48355 3424 48364 3464
rect 48404 3424 48413 3464
rect 48355 3423 48413 3424
rect 48739 3464 48797 3465
rect 48739 3424 48748 3464
rect 48788 3424 48797 3464
rect 48739 3423 48797 3424
rect 50467 3464 50525 3465
rect 50467 3424 50476 3464
rect 50516 3424 50525 3464
rect 50467 3423 50525 3424
rect 50851 3464 50909 3465
rect 50851 3424 50860 3464
rect 50900 3424 50909 3464
rect 50851 3423 50909 3424
rect 51427 3464 51485 3465
rect 51427 3424 51436 3464
rect 51476 3424 51485 3464
rect 51427 3423 51485 3424
rect 51811 3464 51869 3465
rect 51811 3424 51820 3464
rect 51860 3424 51869 3464
rect 51811 3423 51869 3424
rect 52195 3464 52253 3465
rect 52195 3424 52204 3464
rect 52244 3424 52253 3464
rect 52195 3423 52253 3424
rect 53155 3464 53213 3465
rect 53155 3424 53164 3464
rect 53204 3424 53213 3464
rect 53155 3423 53213 3424
rect 53539 3464 53597 3465
rect 53539 3424 53548 3464
rect 53588 3424 53597 3464
rect 53539 3423 53597 3424
rect 53923 3464 53981 3465
rect 53923 3424 53932 3464
rect 53972 3424 53981 3464
rect 53923 3423 53981 3424
rect 54307 3464 54365 3465
rect 54307 3424 54316 3464
rect 54356 3424 54365 3464
rect 54307 3423 54365 3424
rect 55267 3464 55325 3465
rect 55267 3424 55276 3464
rect 55316 3424 55325 3464
rect 55267 3423 55325 3424
rect 55651 3464 55709 3465
rect 55651 3424 55660 3464
rect 55700 3424 55709 3464
rect 55651 3423 55709 3424
rect 56035 3464 56093 3465
rect 56035 3424 56044 3464
rect 56084 3424 56093 3464
rect 56035 3423 56093 3424
rect 56419 3464 56477 3465
rect 56419 3424 56428 3464
rect 56468 3424 56477 3464
rect 56419 3423 56477 3424
rect 56803 3464 56861 3465
rect 56803 3424 56812 3464
rect 56852 3424 56861 3464
rect 56803 3423 56861 3424
rect 57763 3464 57821 3465
rect 57763 3424 57772 3464
rect 57812 3424 57821 3464
rect 57763 3423 57821 3424
rect 58147 3464 58205 3465
rect 58147 3424 58156 3464
rect 58196 3424 58205 3464
rect 58147 3423 58205 3424
rect 58531 3464 58589 3465
rect 58531 3424 58540 3464
rect 58580 3424 58589 3464
rect 58531 3423 58589 3424
rect 58915 3464 58973 3465
rect 58915 3424 58924 3464
rect 58964 3424 58973 3464
rect 58915 3423 58973 3424
rect 60739 3464 60797 3465
rect 60739 3424 60748 3464
rect 60788 3424 60797 3464
rect 60739 3423 60797 3424
rect 61123 3464 61181 3465
rect 61123 3424 61132 3464
rect 61172 3424 61181 3464
rect 61123 3423 61181 3424
rect 61507 3464 61565 3465
rect 61507 3424 61516 3464
rect 61556 3424 61565 3464
rect 61507 3423 61565 3424
rect 61891 3464 61949 3465
rect 61891 3424 61900 3464
rect 61940 3424 61949 3464
rect 61891 3423 61949 3424
rect 62275 3464 62333 3465
rect 62275 3424 62284 3464
rect 62324 3424 62333 3464
rect 62275 3423 62333 3424
rect 63235 3464 63293 3465
rect 63235 3424 63244 3464
rect 63284 3424 63293 3464
rect 63235 3423 63293 3424
rect 63619 3464 63677 3465
rect 63619 3424 63628 3464
rect 63668 3424 63677 3464
rect 63619 3423 63677 3424
rect 64003 3464 64061 3465
rect 64003 3424 64012 3464
rect 64052 3424 64061 3464
rect 64003 3423 64061 3424
rect 64387 3464 64445 3465
rect 64387 3424 64396 3464
rect 64436 3424 64445 3464
rect 64387 3423 64445 3424
rect 64771 3464 64829 3465
rect 64771 3424 64780 3464
rect 64820 3424 64829 3464
rect 64771 3423 64829 3424
rect 65155 3464 65213 3465
rect 65155 3424 65164 3464
rect 65204 3424 65213 3464
rect 65155 3423 65213 3424
rect 65539 3464 65597 3465
rect 65539 3424 65548 3464
rect 65588 3424 65597 3464
rect 65539 3423 65597 3424
rect 65923 3464 65981 3465
rect 65923 3424 65932 3464
rect 65972 3424 65981 3464
rect 65923 3423 65981 3424
rect 66307 3464 66365 3465
rect 66307 3424 66316 3464
rect 66356 3424 66365 3464
rect 66307 3423 66365 3424
rect 66691 3464 66749 3465
rect 66691 3424 66700 3464
rect 66740 3424 66749 3464
rect 66691 3423 66749 3424
rect 67075 3464 67133 3465
rect 67075 3424 67084 3464
rect 67124 3424 67133 3464
rect 67075 3423 67133 3424
rect 67459 3464 67517 3465
rect 67459 3424 67468 3464
rect 67508 3424 67517 3464
rect 67459 3423 67517 3424
rect 67843 3464 67901 3465
rect 67843 3424 67852 3464
rect 67892 3424 67901 3464
rect 67843 3423 67901 3424
rect 68227 3464 68285 3465
rect 68227 3424 68236 3464
rect 68276 3424 68285 3464
rect 68227 3423 68285 3424
rect 68611 3464 68669 3465
rect 68611 3424 68620 3464
rect 68660 3424 68669 3464
rect 68611 3423 68669 3424
rect 68995 3464 69053 3465
rect 68995 3424 69004 3464
rect 69044 3424 69053 3464
rect 68995 3423 69053 3424
rect 69379 3464 69437 3465
rect 69379 3424 69388 3464
rect 69428 3424 69437 3464
rect 69379 3423 69437 3424
rect 69763 3464 69821 3465
rect 69763 3424 69772 3464
rect 69812 3424 69821 3464
rect 69763 3423 69821 3424
rect 70147 3464 70205 3465
rect 70147 3424 70156 3464
rect 70196 3424 70205 3464
rect 70915 3464 70973 3465
rect 70147 3423 70205 3424
rect 70541 3451 70599 3452
rect 70541 3411 70550 3451
rect 70590 3411 70599 3451
rect 70915 3424 70924 3464
rect 70964 3424 70973 3464
rect 70915 3423 70973 3424
rect 71299 3464 71357 3465
rect 71299 3424 71308 3464
rect 71348 3424 71357 3464
rect 71299 3423 71357 3424
rect 71683 3464 71741 3465
rect 71683 3424 71692 3464
rect 71732 3424 71741 3464
rect 71683 3423 71741 3424
rect 72067 3464 72125 3465
rect 72067 3424 72076 3464
rect 72116 3424 72125 3464
rect 72067 3423 72125 3424
rect 72451 3464 72509 3465
rect 72451 3424 72460 3464
rect 72500 3424 72509 3464
rect 72451 3423 72509 3424
rect 72835 3464 72893 3465
rect 72835 3424 72844 3464
rect 72884 3424 72893 3464
rect 72835 3423 72893 3424
rect 73219 3464 73277 3465
rect 73219 3424 73228 3464
rect 73268 3424 73277 3464
rect 73219 3423 73277 3424
rect 73603 3464 73661 3465
rect 73603 3424 73612 3464
rect 73652 3424 73661 3464
rect 73603 3423 73661 3424
rect 73987 3464 74045 3465
rect 73987 3424 73996 3464
rect 74036 3424 74045 3464
rect 73987 3423 74045 3424
rect 74371 3464 74429 3465
rect 74371 3424 74380 3464
rect 74420 3424 74429 3464
rect 74371 3423 74429 3424
rect 74755 3464 74813 3465
rect 74755 3424 74764 3464
rect 74804 3424 74813 3464
rect 74755 3423 74813 3424
rect 75139 3464 75197 3465
rect 75139 3424 75148 3464
rect 75188 3424 75197 3464
rect 75139 3423 75197 3424
rect 75523 3464 75581 3465
rect 75523 3424 75532 3464
rect 75572 3424 75581 3464
rect 75907 3435 75916 3475
rect 75956 3435 75965 3475
rect 75907 3434 75965 3435
rect 76291 3464 76349 3465
rect 75523 3423 75581 3424
rect 76291 3424 76300 3464
rect 76340 3424 76349 3464
rect 76291 3423 76349 3424
rect 76675 3464 76733 3465
rect 76675 3424 76684 3464
rect 76724 3424 76733 3464
rect 76675 3423 76733 3424
rect 77059 3464 77117 3465
rect 77059 3424 77068 3464
rect 77108 3424 77117 3464
rect 77059 3423 77117 3424
rect 77443 3464 77501 3465
rect 77443 3424 77452 3464
rect 77492 3424 77501 3464
rect 77443 3423 77501 3424
rect 77827 3464 77885 3465
rect 77827 3424 77836 3464
rect 77876 3424 77885 3464
rect 77827 3423 77885 3424
rect 78211 3464 78269 3465
rect 78211 3424 78220 3464
rect 78260 3424 78269 3464
rect 78211 3423 78269 3424
rect 78595 3464 78653 3465
rect 78595 3424 78604 3464
rect 78644 3424 78653 3464
rect 78595 3423 78653 3424
rect 78979 3464 79037 3465
rect 78979 3424 78988 3464
rect 79028 3424 79037 3464
rect 78979 3423 79037 3424
rect 79363 3464 79421 3465
rect 79363 3424 79372 3464
rect 79412 3424 79421 3464
rect 79363 3423 79421 3424
rect 79747 3464 79805 3465
rect 79747 3424 79756 3464
rect 79796 3424 79805 3464
rect 79747 3423 79805 3424
rect 80131 3464 80189 3465
rect 80131 3424 80140 3464
rect 80180 3424 80189 3464
rect 80131 3423 80189 3424
rect 80515 3464 80573 3465
rect 80515 3424 80524 3464
rect 80564 3424 80573 3464
rect 80515 3423 80573 3424
rect 82435 3464 82493 3465
rect 82435 3424 82444 3464
rect 82484 3424 82493 3464
rect 82435 3423 82493 3424
rect 82819 3464 82877 3465
rect 82819 3424 82828 3464
rect 82868 3424 82877 3464
rect 82819 3423 82877 3424
rect 83203 3464 83261 3465
rect 83203 3424 83212 3464
rect 83252 3424 83261 3464
rect 83203 3423 83261 3424
rect 83587 3464 83645 3465
rect 83587 3424 83596 3464
rect 83636 3424 83645 3464
rect 83587 3423 83645 3424
rect 83971 3464 84029 3465
rect 83971 3424 83980 3464
rect 84020 3424 84029 3464
rect 83971 3423 84029 3424
rect 84355 3464 84413 3465
rect 84355 3424 84364 3464
rect 84404 3424 84413 3464
rect 84355 3423 84413 3424
rect 84739 3464 84797 3465
rect 84739 3424 84748 3464
rect 84788 3424 84797 3464
rect 84739 3423 84797 3424
rect 85507 3464 85565 3465
rect 85507 3424 85516 3464
rect 85556 3424 85565 3464
rect 85507 3423 85565 3424
rect 85891 3464 85949 3465
rect 85891 3424 85900 3464
rect 85940 3424 85949 3464
rect 85891 3423 85949 3424
rect 86275 3464 86333 3465
rect 86275 3424 86284 3464
rect 86324 3424 86333 3464
rect 86275 3423 86333 3424
rect 86659 3464 86717 3465
rect 86659 3424 86668 3464
rect 86708 3424 86717 3464
rect 86659 3423 86717 3424
rect 87043 3464 87101 3465
rect 87043 3424 87052 3464
rect 87092 3424 87101 3464
rect 87043 3423 87101 3424
rect 87427 3464 87485 3465
rect 87427 3424 87436 3464
rect 87476 3424 87485 3464
rect 87427 3423 87485 3424
rect 87811 3464 87869 3465
rect 87811 3424 87820 3464
rect 87860 3424 87869 3464
rect 87811 3423 87869 3424
rect 88195 3464 88253 3465
rect 88195 3424 88204 3464
rect 88244 3424 88253 3464
rect 88195 3423 88253 3424
rect 88579 3464 88637 3465
rect 88579 3424 88588 3464
rect 88628 3424 88637 3464
rect 88579 3423 88637 3424
rect 88963 3464 89021 3465
rect 88963 3424 88972 3464
rect 89012 3424 89021 3464
rect 88963 3423 89021 3424
rect 89347 3464 89405 3465
rect 89347 3424 89356 3464
rect 89396 3424 89405 3464
rect 89347 3423 89405 3424
rect 89731 3464 89789 3465
rect 89731 3424 89740 3464
rect 89780 3424 89789 3464
rect 89731 3423 89789 3424
rect 90115 3464 90173 3465
rect 90115 3424 90124 3464
rect 90164 3424 90173 3464
rect 90115 3423 90173 3424
rect 90499 3464 90557 3465
rect 90499 3424 90508 3464
rect 90548 3424 90557 3464
rect 90499 3423 90557 3424
rect 90883 3464 90941 3465
rect 90883 3424 90892 3464
rect 90932 3424 90941 3464
rect 90883 3423 90941 3424
rect 91267 3464 91325 3465
rect 91267 3424 91276 3464
rect 91316 3424 91325 3464
rect 91267 3423 91325 3424
rect 91651 3464 91709 3465
rect 91651 3424 91660 3464
rect 91700 3424 91709 3464
rect 91651 3423 91709 3424
rect 92035 3464 92093 3465
rect 92035 3424 92044 3464
rect 92084 3424 92093 3464
rect 92035 3423 92093 3424
rect 92419 3464 92477 3465
rect 92419 3424 92428 3464
rect 92468 3424 92477 3464
rect 92419 3423 92477 3424
rect 92803 3464 92861 3465
rect 92803 3424 92812 3464
rect 92852 3424 92861 3464
rect 92803 3423 92861 3424
rect 93187 3464 93245 3465
rect 93187 3424 93196 3464
rect 93236 3424 93245 3464
rect 93187 3423 93245 3424
rect 93571 3464 93629 3465
rect 93571 3424 93580 3464
rect 93620 3424 93629 3464
rect 93571 3423 93629 3424
rect 93955 3464 94013 3465
rect 93955 3424 93964 3464
rect 94004 3424 94013 3464
rect 93955 3423 94013 3424
rect 94339 3464 94397 3465
rect 94339 3424 94348 3464
rect 94388 3424 94397 3464
rect 94339 3423 94397 3424
rect 94723 3464 94781 3465
rect 94723 3424 94732 3464
rect 94772 3424 94781 3464
rect 94723 3423 94781 3424
rect 95107 3464 95165 3465
rect 95107 3424 95116 3464
rect 95156 3424 95165 3464
rect 95107 3423 95165 3424
rect 95491 3464 95549 3465
rect 95491 3424 95500 3464
rect 95540 3424 95549 3464
rect 95491 3423 95549 3424
rect 95875 3464 95933 3465
rect 95875 3424 95884 3464
rect 95924 3424 95933 3464
rect 95875 3423 95933 3424
rect 96259 3464 96317 3465
rect 96259 3424 96268 3464
rect 96308 3424 96317 3464
rect 96259 3423 96317 3424
rect 96643 3464 96701 3465
rect 96643 3424 96652 3464
rect 96692 3424 96701 3464
rect 96643 3423 96701 3424
rect 97027 3464 97085 3465
rect 97027 3424 97036 3464
rect 97076 3424 97085 3464
rect 97027 3423 97085 3424
rect 97411 3464 97469 3465
rect 97411 3424 97420 3464
rect 97460 3424 97469 3464
rect 97411 3423 97469 3424
rect 97795 3464 97853 3465
rect 97795 3424 97804 3464
rect 97844 3424 97853 3464
rect 97795 3423 97853 3424
rect 98179 3464 98237 3465
rect 98179 3424 98188 3464
rect 98228 3424 98237 3464
rect 98179 3423 98237 3424
rect 98563 3464 98621 3465
rect 98563 3424 98572 3464
rect 98612 3424 98621 3464
rect 98563 3423 98621 3424
rect 70541 3410 70599 3411
rect 17731 3380 17789 3381
rect 17731 3340 17740 3380
rect 17780 3340 17789 3380
rect 17731 3339 17789 3340
rect 17923 3380 17981 3381
rect 17923 3340 17932 3380
rect 17972 3340 17981 3380
rect 17923 3339 17981 3340
rect 34723 3380 34781 3381
rect 34723 3340 34732 3380
rect 34772 3340 34781 3380
rect 34723 3339 34781 3340
rect 34915 3380 34973 3381
rect 34915 3340 34924 3380
rect 34964 3340 34973 3380
rect 34915 3339 34973 3340
rect 46051 3380 46109 3381
rect 46051 3340 46060 3380
rect 46100 3340 46109 3380
rect 46051 3339 46109 3340
rect 46251 3380 46293 3389
rect 46251 3340 46252 3380
rect 46292 3340 46293 3380
rect 46251 3331 46293 3340
rect 46339 3380 46397 3381
rect 46339 3340 46348 3380
rect 46388 3340 46397 3380
rect 46339 3339 46397 3340
rect 47491 3380 47549 3381
rect 47491 3340 47500 3380
rect 47540 3340 47549 3380
rect 47491 3339 47549 3340
rect 49131 3380 49173 3389
rect 49131 3340 49132 3380
rect 49172 3340 49173 3380
rect 49131 3331 49173 3340
rect 49323 3380 49365 3389
rect 49323 3340 49324 3380
rect 49364 3340 49365 3380
rect 49323 3331 49365 3340
rect 49611 3380 49653 3389
rect 49611 3340 49612 3380
rect 49652 3340 49653 3380
rect 49611 3331 49653 3340
rect 50091 3380 50133 3389
rect 50091 3340 50092 3380
rect 50132 3340 50133 3380
rect 50091 3331 50133 3340
rect 52683 3380 52725 3389
rect 52683 3340 52684 3380
rect 52724 3340 52725 3380
rect 52683 3331 52725 3340
rect 54795 3380 54837 3389
rect 54795 3340 54796 3380
rect 54836 3340 54837 3380
rect 54795 3331 54837 3340
rect 57291 3380 57333 3389
rect 57291 3340 57292 3380
rect 57332 3340 57333 3380
rect 57291 3331 57333 3340
rect 59491 3380 59549 3381
rect 59491 3340 59500 3380
rect 59540 3340 59549 3380
rect 59491 3339 59549 3340
rect 59683 3380 59741 3381
rect 59683 3340 59692 3380
rect 59732 3340 59741 3380
rect 59683 3339 59741 3340
rect 60067 3380 60125 3381
rect 60067 3340 60076 3380
rect 60116 3340 60125 3380
rect 60067 3339 60125 3340
rect 60259 3380 60317 3381
rect 60259 3340 60268 3380
rect 60308 3340 60317 3380
rect 60259 3339 60317 3340
rect 62563 3380 62621 3381
rect 62563 3340 62572 3380
rect 62612 3340 62621 3380
rect 62563 3339 62621 3340
rect 62755 3380 62813 3381
rect 62755 3340 62764 3380
rect 62804 3340 62813 3380
rect 62755 3339 62813 3340
rect 81195 3380 81237 3389
rect 81195 3340 81196 3380
rect 81236 3340 81237 3380
rect 81195 3331 81237 3340
rect 84939 3380 84981 3389
rect 84939 3340 84940 3380
rect 84980 3340 84981 3380
rect 84939 3331 84981 3340
rect 85131 3380 85173 3389
rect 85131 3340 85132 3380
rect 85172 3340 85173 3380
rect 85131 3331 85173 3340
rect 46627 3296 46685 3297
rect 46627 3256 46636 3296
rect 46676 3256 46685 3296
rect 46627 3255 46685 3256
rect 49227 3296 49269 3305
rect 49227 3256 49228 3296
rect 49268 3256 49269 3296
rect 49227 3247 49269 3256
rect 1419 3212 1461 3221
rect 1419 3172 1420 3212
rect 1460 3172 1461 3212
rect 1419 3163 1461 3172
rect 1803 3212 1845 3221
rect 1803 3172 1804 3212
rect 1844 3172 1845 3212
rect 1803 3163 1845 3172
rect 2187 3212 2229 3221
rect 2187 3172 2188 3212
rect 2228 3172 2229 3212
rect 2187 3163 2229 3172
rect 2571 3212 2613 3221
rect 2571 3172 2572 3212
rect 2612 3172 2613 3212
rect 2571 3163 2613 3172
rect 2955 3212 2997 3221
rect 2955 3172 2956 3212
rect 2996 3172 2997 3212
rect 2955 3163 2997 3172
rect 3339 3212 3381 3221
rect 3339 3172 3340 3212
rect 3380 3172 3381 3212
rect 3339 3163 3381 3172
rect 3723 3212 3765 3221
rect 3723 3172 3724 3212
rect 3764 3172 3765 3212
rect 3723 3163 3765 3172
rect 4107 3212 4149 3221
rect 4107 3172 4108 3212
rect 4148 3172 4149 3212
rect 4107 3163 4149 3172
rect 4491 3212 4533 3221
rect 4491 3172 4492 3212
rect 4532 3172 4533 3212
rect 4491 3163 4533 3172
rect 4875 3212 4917 3221
rect 4875 3172 4876 3212
rect 4916 3172 4917 3212
rect 4875 3163 4917 3172
rect 5259 3212 5301 3221
rect 5259 3172 5260 3212
rect 5300 3172 5301 3212
rect 5259 3163 5301 3172
rect 5643 3212 5685 3221
rect 5643 3172 5644 3212
rect 5684 3172 5685 3212
rect 5643 3163 5685 3172
rect 6027 3212 6069 3221
rect 6027 3172 6028 3212
rect 6068 3172 6069 3212
rect 6027 3163 6069 3172
rect 6411 3212 6453 3221
rect 6411 3172 6412 3212
rect 6452 3172 6453 3212
rect 6411 3163 6453 3172
rect 6795 3212 6837 3221
rect 6795 3172 6796 3212
rect 6836 3172 6837 3212
rect 6795 3163 6837 3172
rect 7179 3212 7221 3221
rect 7179 3172 7180 3212
rect 7220 3172 7221 3212
rect 7179 3163 7221 3172
rect 7563 3212 7605 3221
rect 7563 3172 7564 3212
rect 7604 3172 7605 3212
rect 7563 3163 7605 3172
rect 7947 3212 7989 3221
rect 7947 3172 7948 3212
rect 7988 3172 7989 3212
rect 7947 3163 7989 3172
rect 8331 3212 8373 3221
rect 8331 3172 8332 3212
rect 8372 3172 8373 3212
rect 8331 3163 8373 3172
rect 8715 3212 8757 3221
rect 8715 3172 8716 3212
rect 8756 3172 8757 3212
rect 8715 3163 8757 3172
rect 9099 3212 9141 3221
rect 9099 3172 9100 3212
rect 9140 3172 9141 3212
rect 9099 3163 9141 3172
rect 9483 3212 9525 3221
rect 9483 3172 9484 3212
rect 9524 3172 9525 3212
rect 9483 3163 9525 3172
rect 9867 3212 9909 3221
rect 9867 3172 9868 3212
rect 9908 3172 9909 3212
rect 9867 3163 9909 3172
rect 10251 3212 10293 3221
rect 10251 3172 10252 3212
rect 10292 3172 10293 3212
rect 10251 3163 10293 3172
rect 10635 3212 10677 3221
rect 10635 3172 10636 3212
rect 10676 3172 10677 3212
rect 10635 3163 10677 3172
rect 11019 3212 11061 3221
rect 11019 3172 11020 3212
rect 11060 3172 11061 3212
rect 11019 3163 11061 3172
rect 11403 3212 11445 3221
rect 11403 3172 11404 3212
rect 11444 3172 11445 3212
rect 11403 3163 11445 3172
rect 11787 3212 11829 3221
rect 11787 3172 11788 3212
rect 11828 3172 11829 3212
rect 11787 3163 11829 3172
rect 12171 3212 12213 3221
rect 12171 3172 12172 3212
rect 12212 3172 12213 3212
rect 12171 3163 12213 3172
rect 12555 3212 12597 3221
rect 12555 3172 12556 3212
rect 12596 3172 12597 3212
rect 12555 3163 12597 3172
rect 12939 3212 12981 3221
rect 12939 3172 12940 3212
rect 12980 3172 12981 3212
rect 12939 3163 12981 3172
rect 13323 3212 13365 3221
rect 13323 3172 13324 3212
rect 13364 3172 13365 3212
rect 13323 3163 13365 3172
rect 13707 3212 13749 3221
rect 13707 3172 13708 3212
rect 13748 3172 13749 3212
rect 13707 3163 13749 3172
rect 14091 3212 14133 3221
rect 14091 3172 14092 3212
rect 14132 3172 14133 3212
rect 14091 3163 14133 3172
rect 14475 3212 14517 3221
rect 14475 3172 14476 3212
rect 14516 3172 14517 3212
rect 14475 3163 14517 3172
rect 14859 3212 14901 3221
rect 14859 3172 14860 3212
rect 14900 3172 14901 3212
rect 14859 3163 14901 3172
rect 15243 3212 15285 3221
rect 15243 3172 15244 3212
rect 15284 3172 15285 3212
rect 15243 3163 15285 3172
rect 15627 3212 15669 3221
rect 15627 3172 15628 3212
rect 15668 3172 15669 3212
rect 15627 3163 15669 3172
rect 16011 3212 16053 3221
rect 16011 3172 16012 3212
rect 16052 3172 16053 3212
rect 16011 3163 16053 3172
rect 16395 3212 16437 3221
rect 16395 3172 16396 3212
rect 16436 3172 16437 3212
rect 16395 3163 16437 3172
rect 16779 3212 16821 3221
rect 16779 3172 16780 3212
rect 16820 3172 16821 3212
rect 16779 3163 16821 3172
rect 17163 3212 17205 3221
rect 17163 3172 17164 3212
rect 17204 3172 17205 3212
rect 17163 3163 17205 3172
rect 17547 3212 17589 3221
rect 17547 3172 17548 3212
rect 17588 3172 17589 3212
rect 17547 3163 17589 3172
rect 18699 3212 18741 3221
rect 18699 3172 18700 3212
rect 18740 3172 18741 3212
rect 18699 3163 18741 3172
rect 19083 3212 19125 3221
rect 19083 3172 19084 3212
rect 19124 3172 19125 3212
rect 19083 3163 19125 3172
rect 19467 3212 19509 3221
rect 19467 3172 19468 3212
rect 19508 3172 19509 3212
rect 19467 3163 19509 3172
rect 19851 3212 19893 3221
rect 19851 3172 19852 3212
rect 19892 3172 19893 3212
rect 19851 3163 19893 3172
rect 20235 3212 20277 3221
rect 20235 3172 20236 3212
rect 20276 3172 20277 3212
rect 20235 3163 20277 3172
rect 20619 3212 20661 3221
rect 20619 3172 20620 3212
rect 20660 3172 20661 3212
rect 20619 3163 20661 3172
rect 21003 3212 21045 3221
rect 21003 3172 21004 3212
rect 21044 3172 21045 3212
rect 21003 3163 21045 3172
rect 21387 3212 21429 3221
rect 21387 3172 21388 3212
rect 21428 3172 21429 3212
rect 21387 3163 21429 3172
rect 21771 3212 21813 3221
rect 21771 3172 21772 3212
rect 21812 3172 21813 3212
rect 21771 3163 21813 3172
rect 22155 3212 22197 3221
rect 22155 3172 22156 3212
rect 22196 3172 22197 3212
rect 22155 3163 22197 3172
rect 22539 3212 22581 3221
rect 22539 3172 22540 3212
rect 22580 3172 22581 3212
rect 22539 3163 22581 3172
rect 22923 3212 22965 3221
rect 22923 3172 22924 3212
rect 22964 3172 22965 3212
rect 22923 3163 22965 3172
rect 23307 3212 23349 3221
rect 23307 3172 23308 3212
rect 23348 3172 23349 3212
rect 23307 3163 23349 3172
rect 23691 3212 23733 3221
rect 23691 3172 23692 3212
rect 23732 3172 23733 3212
rect 23691 3163 23733 3172
rect 24075 3212 24117 3221
rect 24075 3172 24076 3212
rect 24116 3172 24117 3212
rect 24075 3163 24117 3172
rect 24459 3212 24501 3221
rect 24459 3172 24460 3212
rect 24500 3172 24501 3212
rect 24459 3163 24501 3172
rect 24843 3212 24885 3221
rect 24843 3172 24844 3212
rect 24884 3172 24885 3212
rect 24843 3163 24885 3172
rect 25227 3212 25269 3221
rect 25227 3172 25228 3212
rect 25268 3172 25269 3212
rect 25227 3163 25269 3172
rect 25611 3212 25653 3221
rect 25611 3172 25612 3212
rect 25652 3172 25653 3212
rect 25611 3163 25653 3172
rect 25995 3212 26037 3221
rect 25995 3172 25996 3212
rect 26036 3172 26037 3212
rect 25995 3163 26037 3172
rect 26379 3212 26421 3221
rect 26379 3172 26380 3212
rect 26420 3172 26421 3212
rect 26379 3163 26421 3172
rect 26763 3212 26805 3221
rect 26763 3172 26764 3212
rect 26804 3172 26805 3212
rect 26763 3163 26805 3172
rect 27147 3212 27189 3221
rect 27147 3172 27148 3212
rect 27188 3172 27189 3212
rect 27147 3163 27189 3172
rect 27531 3212 27573 3221
rect 27531 3172 27532 3212
rect 27572 3172 27573 3212
rect 27531 3163 27573 3172
rect 27915 3212 27957 3221
rect 27915 3172 27916 3212
rect 27956 3172 27957 3212
rect 27915 3163 27957 3172
rect 28299 3212 28341 3221
rect 28299 3172 28300 3212
rect 28340 3172 28341 3212
rect 28299 3163 28341 3172
rect 28683 3212 28725 3221
rect 28683 3172 28684 3212
rect 28724 3172 28725 3212
rect 28683 3163 28725 3172
rect 29067 3212 29109 3221
rect 29067 3172 29068 3212
rect 29108 3172 29109 3212
rect 29067 3163 29109 3172
rect 29451 3212 29493 3221
rect 29451 3172 29452 3212
rect 29492 3172 29493 3212
rect 29451 3163 29493 3172
rect 29835 3212 29877 3221
rect 29835 3172 29836 3212
rect 29876 3172 29877 3212
rect 29835 3163 29877 3172
rect 30219 3212 30261 3221
rect 30219 3172 30220 3212
rect 30260 3172 30261 3212
rect 30219 3163 30261 3172
rect 30603 3212 30645 3221
rect 30603 3172 30604 3212
rect 30644 3172 30645 3212
rect 30603 3163 30645 3172
rect 30987 3212 31029 3221
rect 30987 3172 30988 3212
rect 31028 3172 31029 3212
rect 30987 3163 31029 3172
rect 31371 3212 31413 3221
rect 31371 3172 31372 3212
rect 31412 3172 31413 3212
rect 31371 3163 31413 3172
rect 31755 3212 31797 3221
rect 31755 3172 31756 3212
rect 31796 3172 31797 3212
rect 31755 3163 31797 3172
rect 32139 3212 32181 3221
rect 32139 3172 32140 3212
rect 32180 3172 32181 3212
rect 32139 3163 32181 3172
rect 32523 3212 32565 3221
rect 32523 3172 32524 3212
rect 32564 3172 32565 3212
rect 32523 3163 32565 3172
rect 32907 3212 32949 3221
rect 32907 3172 32908 3212
rect 32948 3172 32949 3212
rect 32907 3163 32949 3172
rect 33291 3212 33333 3221
rect 33291 3172 33292 3212
rect 33332 3172 33333 3212
rect 33291 3163 33333 3172
rect 33675 3212 33717 3221
rect 33675 3172 33676 3212
rect 33716 3172 33717 3212
rect 33675 3163 33717 3172
rect 34059 3212 34101 3221
rect 34059 3172 34060 3212
rect 34100 3172 34101 3212
rect 34059 3163 34101 3172
rect 34443 3212 34485 3221
rect 34443 3172 34444 3212
rect 34484 3172 34485 3212
rect 34443 3163 34485 3172
rect 34923 3212 34965 3221
rect 34923 3172 34924 3212
rect 34964 3172 34965 3212
rect 34923 3163 34965 3172
rect 35499 3212 35541 3221
rect 35499 3172 35500 3212
rect 35540 3172 35541 3212
rect 35499 3163 35541 3172
rect 35883 3212 35925 3221
rect 35883 3172 35884 3212
rect 35924 3172 35925 3212
rect 35883 3163 35925 3172
rect 36267 3212 36309 3221
rect 36267 3172 36268 3212
rect 36308 3172 36309 3212
rect 36267 3163 36309 3172
rect 36651 3212 36693 3221
rect 36651 3172 36652 3212
rect 36692 3172 36693 3212
rect 36651 3163 36693 3172
rect 37035 3212 37077 3221
rect 37035 3172 37036 3212
rect 37076 3172 37077 3212
rect 37035 3163 37077 3172
rect 37419 3212 37461 3221
rect 37419 3172 37420 3212
rect 37460 3172 37461 3212
rect 37419 3163 37461 3172
rect 37803 3212 37845 3221
rect 37803 3172 37804 3212
rect 37844 3172 37845 3212
rect 37803 3163 37845 3172
rect 38187 3212 38229 3221
rect 38187 3172 38188 3212
rect 38228 3172 38229 3212
rect 38187 3163 38229 3172
rect 38571 3212 38613 3221
rect 38571 3172 38572 3212
rect 38612 3172 38613 3212
rect 38571 3163 38613 3172
rect 38955 3212 38997 3221
rect 38955 3172 38956 3212
rect 38996 3172 38997 3212
rect 38955 3163 38997 3172
rect 39339 3212 39381 3221
rect 39339 3172 39340 3212
rect 39380 3172 39381 3212
rect 39339 3163 39381 3172
rect 39723 3212 39765 3221
rect 39723 3172 39724 3212
rect 39764 3172 39765 3212
rect 39723 3163 39765 3172
rect 40107 3212 40149 3221
rect 40107 3172 40108 3212
rect 40148 3172 40149 3212
rect 40107 3163 40149 3172
rect 40491 3212 40533 3221
rect 40491 3172 40492 3212
rect 40532 3172 40533 3212
rect 40491 3163 40533 3172
rect 40875 3212 40917 3221
rect 40875 3172 40876 3212
rect 40916 3172 40917 3212
rect 40875 3163 40917 3172
rect 41259 3212 41301 3221
rect 41259 3172 41260 3212
rect 41300 3172 41301 3212
rect 41259 3163 41301 3172
rect 41643 3212 41685 3221
rect 41643 3172 41644 3212
rect 41684 3172 41685 3212
rect 41643 3163 41685 3172
rect 42027 3212 42069 3221
rect 42027 3172 42028 3212
rect 42068 3172 42069 3212
rect 42027 3163 42069 3172
rect 42411 3212 42453 3221
rect 42411 3172 42412 3212
rect 42452 3172 42453 3212
rect 42411 3163 42453 3172
rect 42795 3212 42837 3221
rect 42795 3172 42796 3212
rect 42836 3172 42837 3212
rect 42795 3163 42837 3172
rect 43179 3212 43221 3221
rect 43179 3172 43180 3212
rect 43220 3172 43221 3212
rect 43179 3163 43221 3172
rect 43563 3212 43605 3221
rect 43563 3172 43564 3212
rect 43604 3172 43605 3212
rect 43563 3163 43605 3172
rect 43947 3212 43989 3221
rect 43947 3172 43948 3212
rect 43988 3172 43989 3212
rect 43947 3163 43989 3172
rect 44331 3212 44373 3221
rect 44331 3172 44332 3212
rect 44372 3172 44373 3212
rect 44331 3163 44373 3172
rect 44715 3212 44757 3221
rect 44715 3172 44716 3212
rect 44756 3172 44757 3212
rect 44715 3163 44757 3172
rect 45099 3212 45141 3221
rect 45099 3172 45100 3212
rect 45140 3172 45141 3212
rect 45099 3163 45141 3172
rect 45483 3212 45525 3221
rect 45483 3172 45484 3212
rect 45524 3172 45525 3212
rect 45483 3163 45525 3172
rect 45867 3212 45909 3221
rect 45867 3172 45868 3212
rect 45908 3172 45909 3212
rect 45867 3163 45909 3172
rect 46059 3212 46101 3221
rect 46059 3172 46060 3212
rect 46100 3172 46101 3212
rect 46059 3163 46101 3172
rect 48171 3212 48213 3221
rect 48171 3172 48172 3212
rect 48212 3172 48213 3212
rect 48171 3163 48213 3172
rect 48555 3212 48597 3221
rect 48555 3172 48556 3212
rect 48596 3172 48597 3212
rect 48555 3163 48597 3172
rect 48939 3212 48981 3221
rect 48939 3172 48940 3212
rect 48980 3172 48981 3212
rect 48939 3163 48981 3172
rect 50667 3212 50709 3221
rect 50667 3172 50668 3212
rect 50708 3172 50709 3212
rect 50667 3163 50709 3172
rect 51051 3212 51093 3221
rect 51051 3172 51052 3212
rect 51092 3172 51093 3212
rect 51051 3163 51093 3172
rect 51243 3212 51285 3221
rect 51243 3172 51244 3212
rect 51284 3172 51285 3212
rect 51243 3163 51285 3172
rect 51627 3212 51669 3221
rect 51627 3172 51628 3212
rect 51668 3172 51669 3212
rect 51627 3163 51669 3172
rect 52011 3212 52053 3221
rect 52011 3172 52012 3212
rect 52052 3172 52053 3212
rect 52011 3163 52053 3172
rect 52971 3212 53013 3221
rect 52971 3172 52972 3212
rect 53012 3172 53013 3212
rect 52971 3163 53013 3172
rect 53355 3212 53397 3221
rect 53355 3172 53356 3212
rect 53396 3172 53397 3212
rect 53355 3163 53397 3172
rect 53739 3212 53781 3221
rect 53739 3172 53740 3212
rect 53780 3172 53781 3212
rect 53739 3163 53781 3172
rect 54123 3212 54165 3221
rect 54123 3172 54124 3212
rect 54164 3172 54165 3212
rect 54123 3163 54165 3172
rect 54603 3212 54645 3221
rect 54603 3172 54604 3212
rect 54644 3172 54645 3212
rect 54603 3163 54645 3172
rect 55083 3212 55125 3221
rect 55083 3172 55084 3212
rect 55124 3172 55125 3212
rect 55083 3163 55125 3172
rect 55467 3212 55509 3221
rect 55467 3172 55468 3212
rect 55508 3172 55509 3212
rect 55467 3163 55509 3172
rect 55851 3212 55893 3221
rect 55851 3172 55852 3212
rect 55892 3172 55893 3212
rect 55851 3163 55893 3172
rect 56235 3212 56277 3221
rect 56235 3172 56236 3212
rect 56276 3172 56277 3212
rect 56235 3163 56277 3172
rect 56619 3212 56661 3221
rect 56619 3172 56620 3212
rect 56660 3172 56661 3212
rect 56619 3163 56661 3172
rect 57099 3212 57141 3221
rect 57099 3172 57100 3212
rect 57140 3172 57141 3212
rect 57099 3163 57141 3172
rect 57579 3212 57621 3221
rect 57579 3172 57580 3212
rect 57620 3172 57621 3212
rect 57579 3163 57621 3172
rect 57963 3212 58005 3221
rect 57963 3172 57964 3212
rect 58004 3172 58005 3212
rect 57963 3163 58005 3172
rect 58347 3212 58389 3221
rect 58347 3172 58348 3212
rect 58388 3172 58389 3212
rect 58347 3163 58389 3172
rect 58731 3212 58773 3221
rect 58731 3172 58732 3212
rect 58772 3172 58773 3212
rect 58731 3163 58773 3172
rect 59499 3212 59541 3221
rect 59499 3172 59500 3212
rect 59540 3172 59541 3212
rect 59499 3163 59541 3172
rect 60555 3212 60597 3221
rect 60555 3172 60556 3212
rect 60596 3172 60597 3212
rect 60555 3163 60597 3172
rect 60939 3212 60981 3221
rect 60939 3172 60940 3212
rect 60980 3172 60981 3212
rect 60939 3163 60981 3172
rect 61323 3212 61365 3221
rect 61323 3172 61324 3212
rect 61364 3172 61365 3212
rect 61323 3163 61365 3172
rect 61707 3212 61749 3221
rect 61707 3172 61708 3212
rect 61748 3172 61749 3212
rect 61707 3163 61749 3172
rect 62091 3212 62133 3221
rect 62091 3172 62092 3212
rect 62132 3172 62133 3212
rect 62091 3163 62133 3172
rect 63051 3212 63093 3221
rect 63051 3172 63052 3212
rect 63092 3172 63093 3212
rect 63051 3163 63093 3172
rect 63435 3212 63477 3221
rect 63435 3172 63436 3212
rect 63476 3172 63477 3212
rect 63435 3163 63477 3172
rect 63819 3212 63861 3221
rect 63819 3172 63820 3212
rect 63860 3172 63861 3212
rect 63819 3163 63861 3172
rect 64203 3212 64245 3221
rect 64203 3172 64204 3212
rect 64244 3172 64245 3212
rect 64203 3163 64245 3172
rect 64587 3212 64629 3221
rect 64587 3172 64588 3212
rect 64628 3172 64629 3212
rect 64587 3163 64629 3172
rect 65739 3212 65781 3221
rect 65739 3172 65740 3212
rect 65780 3172 65781 3212
rect 65739 3163 65781 3172
rect 66123 3212 66165 3221
rect 66123 3172 66124 3212
rect 66164 3172 66165 3212
rect 66123 3163 66165 3172
rect 66507 3212 66549 3221
rect 66507 3172 66508 3212
rect 66548 3172 66549 3212
rect 66507 3163 66549 3172
rect 66891 3212 66933 3221
rect 66891 3172 66892 3212
rect 66932 3172 66933 3212
rect 66891 3163 66933 3172
rect 67275 3212 67317 3221
rect 67275 3172 67276 3212
rect 67316 3172 67317 3212
rect 67275 3163 67317 3172
rect 67659 3212 67701 3221
rect 67659 3172 67660 3212
rect 67700 3172 67701 3212
rect 67659 3163 67701 3172
rect 68043 3212 68085 3221
rect 68043 3172 68044 3212
rect 68084 3172 68085 3212
rect 68043 3163 68085 3172
rect 68427 3212 68469 3221
rect 68427 3172 68428 3212
rect 68468 3172 68469 3212
rect 68427 3163 68469 3172
rect 68811 3212 68853 3221
rect 68811 3172 68812 3212
rect 68852 3172 68853 3212
rect 68811 3163 68853 3172
rect 69195 3212 69237 3221
rect 69195 3172 69196 3212
rect 69236 3172 69237 3212
rect 69195 3163 69237 3172
rect 69579 3212 69621 3221
rect 69579 3172 69580 3212
rect 69620 3172 69621 3212
rect 69579 3163 69621 3172
rect 69963 3212 70005 3221
rect 69963 3172 69964 3212
rect 70004 3172 70005 3212
rect 69963 3163 70005 3172
rect 70347 3212 70389 3221
rect 70347 3172 70348 3212
rect 70388 3172 70389 3212
rect 70347 3163 70389 3172
rect 70731 3212 70773 3221
rect 70731 3172 70732 3212
rect 70772 3172 70773 3212
rect 70731 3163 70773 3172
rect 71115 3212 71157 3221
rect 71115 3172 71116 3212
rect 71156 3172 71157 3212
rect 71115 3163 71157 3172
rect 71499 3212 71541 3221
rect 71499 3172 71500 3212
rect 71540 3172 71541 3212
rect 71499 3163 71541 3172
rect 71883 3212 71925 3221
rect 71883 3172 71884 3212
rect 71924 3172 71925 3212
rect 71883 3163 71925 3172
rect 72267 3212 72309 3221
rect 72267 3172 72268 3212
rect 72308 3172 72309 3212
rect 72267 3163 72309 3172
rect 72651 3212 72693 3221
rect 72651 3172 72652 3212
rect 72692 3172 72693 3212
rect 72651 3163 72693 3172
rect 73035 3212 73077 3221
rect 73035 3172 73036 3212
rect 73076 3172 73077 3212
rect 73035 3163 73077 3172
rect 73419 3212 73461 3221
rect 73419 3172 73420 3212
rect 73460 3172 73461 3212
rect 73419 3163 73461 3172
rect 73803 3212 73845 3221
rect 73803 3172 73804 3212
rect 73844 3172 73845 3212
rect 73803 3163 73845 3172
rect 74187 3212 74229 3221
rect 74187 3172 74188 3212
rect 74228 3172 74229 3212
rect 74187 3163 74229 3172
rect 74571 3212 74613 3221
rect 74571 3172 74572 3212
rect 74612 3172 74613 3212
rect 74571 3163 74613 3172
rect 74955 3212 74997 3221
rect 74955 3172 74956 3212
rect 74996 3172 74997 3212
rect 74955 3163 74997 3172
rect 75339 3212 75381 3221
rect 75339 3172 75340 3212
rect 75380 3172 75381 3212
rect 75339 3163 75381 3172
rect 75723 3212 75765 3221
rect 75723 3172 75724 3212
rect 75764 3172 75765 3212
rect 75723 3163 75765 3172
rect 76107 3212 76149 3221
rect 76107 3172 76108 3212
rect 76148 3172 76149 3212
rect 76107 3163 76149 3172
rect 76491 3212 76533 3221
rect 76491 3172 76492 3212
rect 76532 3172 76533 3212
rect 76491 3163 76533 3172
rect 76875 3212 76917 3221
rect 76875 3172 76876 3212
rect 76916 3172 76917 3212
rect 76875 3163 76917 3172
rect 77259 3212 77301 3221
rect 77259 3172 77260 3212
rect 77300 3172 77301 3212
rect 77259 3163 77301 3172
rect 77643 3212 77685 3221
rect 77643 3172 77644 3212
rect 77684 3172 77685 3212
rect 77643 3163 77685 3172
rect 78027 3212 78069 3221
rect 78027 3172 78028 3212
rect 78068 3172 78069 3212
rect 78027 3163 78069 3172
rect 78411 3212 78453 3221
rect 78411 3172 78412 3212
rect 78452 3172 78453 3212
rect 78411 3163 78453 3172
rect 78795 3212 78837 3221
rect 78795 3172 78796 3212
rect 78836 3172 78837 3212
rect 78795 3163 78837 3172
rect 79179 3212 79221 3221
rect 79179 3172 79180 3212
rect 79220 3172 79221 3212
rect 79179 3163 79221 3172
rect 79563 3212 79605 3221
rect 79563 3172 79564 3212
rect 79604 3172 79605 3212
rect 79563 3163 79605 3172
rect 79947 3212 79989 3221
rect 79947 3172 79948 3212
rect 79988 3172 79989 3212
rect 79947 3163 79989 3172
rect 80331 3212 80373 3221
rect 80331 3172 80332 3212
rect 80372 3172 80373 3212
rect 80331 3163 80373 3172
rect 82251 3212 82293 3221
rect 82251 3172 82252 3212
rect 82292 3172 82293 3212
rect 82251 3163 82293 3172
rect 83019 3212 83061 3221
rect 83019 3172 83020 3212
rect 83060 3172 83061 3212
rect 83019 3163 83061 3172
rect 83403 3212 83445 3221
rect 83403 3172 83404 3212
rect 83444 3172 83445 3212
rect 83403 3163 83445 3172
rect 83787 3212 83829 3221
rect 83787 3172 83788 3212
rect 83828 3172 83829 3212
rect 83787 3163 83829 3172
rect 84171 3212 84213 3221
rect 84171 3172 84172 3212
rect 84212 3172 84213 3212
rect 84171 3163 84213 3172
rect 84555 3212 84597 3221
rect 84555 3172 84556 3212
rect 84596 3172 84597 3212
rect 84555 3163 84597 3172
rect 85323 3212 85365 3221
rect 85323 3172 85324 3212
rect 85364 3172 85365 3212
rect 85323 3163 85365 3172
rect 85707 3212 85749 3221
rect 85707 3172 85708 3212
rect 85748 3172 85749 3212
rect 85707 3163 85749 3172
rect 86091 3212 86133 3221
rect 86091 3172 86092 3212
rect 86132 3172 86133 3212
rect 86091 3163 86133 3172
rect 86475 3212 86517 3221
rect 86475 3172 86476 3212
rect 86516 3172 86517 3212
rect 86475 3163 86517 3172
rect 86859 3212 86901 3221
rect 86859 3172 86860 3212
rect 86900 3172 86901 3212
rect 86859 3163 86901 3172
rect 87243 3212 87285 3221
rect 87243 3172 87244 3212
rect 87284 3172 87285 3212
rect 87243 3163 87285 3172
rect 87627 3212 87669 3221
rect 87627 3172 87628 3212
rect 87668 3172 87669 3212
rect 87627 3163 87669 3172
rect 88011 3212 88053 3221
rect 88011 3172 88012 3212
rect 88052 3172 88053 3212
rect 88011 3163 88053 3172
rect 88395 3212 88437 3221
rect 88395 3172 88396 3212
rect 88436 3172 88437 3212
rect 88395 3163 88437 3172
rect 88779 3212 88821 3221
rect 88779 3172 88780 3212
rect 88820 3172 88821 3212
rect 88779 3163 88821 3172
rect 89163 3212 89205 3221
rect 89163 3172 89164 3212
rect 89204 3172 89205 3212
rect 89163 3163 89205 3172
rect 89547 3212 89589 3221
rect 89547 3172 89548 3212
rect 89588 3172 89589 3212
rect 89547 3163 89589 3172
rect 89931 3212 89973 3221
rect 89931 3172 89932 3212
rect 89972 3172 89973 3212
rect 89931 3163 89973 3172
rect 90315 3212 90357 3221
rect 90315 3172 90316 3212
rect 90356 3172 90357 3212
rect 90315 3163 90357 3172
rect 90699 3212 90741 3221
rect 90699 3172 90700 3212
rect 90740 3172 90741 3212
rect 90699 3163 90741 3172
rect 91083 3212 91125 3221
rect 91083 3172 91084 3212
rect 91124 3172 91125 3212
rect 91083 3163 91125 3172
rect 91467 3212 91509 3221
rect 91467 3172 91468 3212
rect 91508 3172 91509 3212
rect 91467 3163 91509 3172
rect 91851 3212 91893 3221
rect 91851 3172 91852 3212
rect 91892 3172 91893 3212
rect 91851 3163 91893 3172
rect 92235 3212 92277 3221
rect 92235 3172 92236 3212
rect 92276 3172 92277 3212
rect 92235 3163 92277 3172
rect 92619 3212 92661 3221
rect 92619 3172 92620 3212
rect 92660 3172 92661 3212
rect 92619 3163 92661 3172
rect 93003 3212 93045 3221
rect 93003 3172 93004 3212
rect 93044 3172 93045 3212
rect 93003 3163 93045 3172
rect 93387 3212 93429 3221
rect 93387 3172 93388 3212
rect 93428 3172 93429 3212
rect 93387 3163 93429 3172
rect 93771 3212 93813 3221
rect 93771 3172 93772 3212
rect 93812 3172 93813 3212
rect 93771 3163 93813 3172
rect 94155 3212 94197 3221
rect 94155 3172 94156 3212
rect 94196 3172 94197 3212
rect 94155 3163 94197 3172
rect 94539 3212 94581 3221
rect 94539 3172 94540 3212
rect 94580 3172 94581 3212
rect 94539 3163 94581 3172
rect 94923 3212 94965 3221
rect 94923 3172 94924 3212
rect 94964 3172 94965 3212
rect 94923 3163 94965 3172
rect 95307 3212 95349 3221
rect 95307 3172 95308 3212
rect 95348 3172 95349 3212
rect 95307 3163 95349 3172
rect 95691 3212 95733 3221
rect 95691 3172 95692 3212
rect 95732 3172 95733 3212
rect 95691 3163 95733 3172
rect 96075 3212 96117 3221
rect 96075 3172 96076 3212
rect 96116 3172 96117 3212
rect 96075 3163 96117 3172
rect 96459 3212 96501 3221
rect 96459 3172 96460 3212
rect 96500 3172 96501 3212
rect 96459 3163 96501 3172
rect 96843 3212 96885 3221
rect 96843 3172 96844 3212
rect 96884 3172 96885 3212
rect 96843 3163 96885 3172
rect 97227 3212 97269 3221
rect 97227 3172 97228 3212
rect 97268 3172 97269 3212
rect 97227 3163 97269 3172
rect 97611 3212 97653 3221
rect 97611 3172 97612 3212
rect 97652 3172 97653 3212
rect 97611 3163 97653 3172
rect 97995 3212 98037 3221
rect 97995 3172 97996 3212
rect 98036 3172 98037 3212
rect 97995 3163 98037 3172
rect 98379 3212 98421 3221
rect 98379 3172 98380 3212
rect 98420 3172 98421 3212
rect 98379 3163 98421 3172
rect 1152 3044 98784 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 65408 3044
rect 65448 3004 65490 3044
rect 65530 3004 65572 3044
rect 65612 3004 65654 3044
rect 65694 3004 65736 3044
rect 65776 3004 80528 3044
rect 80568 3004 80610 3044
rect 80650 3004 80692 3044
rect 80732 3004 80774 3044
rect 80814 3004 80856 3044
rect 80896 3004 95648 3044
rect 95688 3004 95730 3044
rect 95770 3004 95812 3044
rect 95852 3004 95894 3044
rect 95934 3004 95976 3044
rect 96016 3004 98784 3044
rect 1152 2980 98784 3004
<< via1 >>
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 33928 11320 33968 11360
rect 34010 11320 34050 11360
rect 34092 11320 34132 11360
rect 34174 11320 34214 11360
rect 34256 11320 34296 11360
rect 49048 11320 49088 11360
rect 49130 11320 49170 11360
rect 49212 11320 49252 11360
rect 49294 11320 49334 11360
rect 49376 11320 49416 11360
rect 64168 11320 64208 11360
rect 64250 11320 64290 11360
rect 64332 11320 64372 11360
rect 64414 11320 64454 11360
rect 64496 11320 64536 11360
rect 79288 11320 79328 11360
rect 79370 11320 79410 11360
rect 79452 11320 79492 11360
rect 79534 11320 79574 11360
rect 79616 11320 79656 11360
rect 94408 11320 94448 11360
rect 94490 11320 94530 11360
rect 94572 11320 94612 11360
rect 94654 11320 94694 11360
rect 94736 11320 94776 11360
rect 11884 11152 11924 11192
rect 30892 11152 30932 11192
rect 19564 11068 19604 11108
rect 50092 10984 50132 11024
rect 11788 10900 11828 10940
rect 11980 10900 12020 10940
rect 12172 10900 12212 10940
rect 12364 10900 12404 10940
rect 15628 10900 15668 10940
rect 15820 10900 15860 10940
rect 17260 10900 17300 10940
rect 17452 10900 17492 10940
rect 19468 10900 19508 10940
rect 19660 10900 19700 10940
rect 24172 10900 24212 10940
rect 24364 10900 24404 10940
rect 24556 10900 24596 10940
rect 24748 10900 24788 10940
rect 24940 10900 24980 10940
rect 25132 10900 25172 10940
rect 28204 10900 28244 10940
rect 28396 10900 28436 10940
rect 30796 10900 30836 10940
rect 30988 10900 31028 10940
rect 31180 10900 31220 10940
rect 31372 10900 31412 10940
rect 36460 10900 36500 10940
rect 36652 10900 36692 10940
rect 36844 10900 36884 10940
rect 37036 10900 37076 10940
rect 39148 10900 39188 10940
rect 39340 10900 39380 10940
rect 61036 10900 61076 10940
rect 61228 10900 61268 10940
rect 71980 10900 72020 10940
rect 72172 10900 72212 10940
rect 82924 10900 82964 10940
rect 83116 10900 83156 10940
rect 12268 10816 12308 10856
rect 15724 10816 15764 10856
rect 24268 10816 24308 10856
rect 24652 10816 24692 10856
rect 25036 10816 25076 10856
rect 31276 10816 31316 10856
rect 36556 10816 36596 10856
rect 36940 10816 36980 10856
rect 50284 10732 50324 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 65408 10564 65448 10604
rect 65490 10564 65530 10604
rect 65572 10564 65612 10604
rect 65654 10564 65694 10604
rect 65736 10564 65776 10604
rect 80528 10564 80568 10604
rect 80610 10564 80650 10604
rect 80692 10564 80732 10604
rect 80774 10564 80814 10604
rect 80856 10564 80896 10604
rect 95648 10564 95688 10604
rect 95730 10564 95770 10604
rect 95812 10564 95852 10604
rect 95894 10564 95934 10604
rect 95976 10564 96016 10604
rect 57676 10396 57716 10436
rect 10924 10312 10964 10352
rect 19084 10312 19124 10352
rect 19852 10312 19892 10352
rect 23884 10312 23924 10352
rect 36076 10312 36116 10352
rect 36460 10312 36500 10352
rect 49420 10312 49460 10352
rect 84076 10312 84116 10352
rect 88300 10312 88340 10352
rect 10828 10228 10868 10268
rect 11020 10228 11060 10268
rect 11212 10228 11252 10268
rect 11404 10228 11444 10268
rect 11596 10228 11636 10268
rect 11788 10228 11828 10268
rect 11980 10228 12020 10268
rect 12172 10228 12212 10268
rect 12364 10249 12404 10289
rect 12556 10228 12596 10268
rect 12748 10228 12788 10268
rect 12940 10228 12980 10268
rect 14572 10228 14612 10268
rect 14764 10228 14804 10268
rect 14956 10228 14996 10268
rect 15148 10228 15188 10268
rect 15340 10228 15380 10268
rect 15532 10228 15572 10268
rect 15724 10228 15764 10268
rect 15916 10228 15956 10268
rect 16108 10228 16148 10268
rect 16300 10228 16340 10268
rect 18604 10228 18644 10268
rect 18796 10228 18836 10268
rect 18988 10228 19028 10268
rect 19180 10228 19220 10268
rect 19372 10228 19412 10268
rect 19564 10228 19604 10268
rect 19756 10228 19796 10268
rect 19948 10228 19988 10268
rect 20131 10213 20171 10253
rect 20332 10228 20372 10268
rect 21676 10228 21716 10268
rect 23788 10228 23828 10268
rect 23980 10228 24020 10268
rect 24172 10228 24212 10268
rect 24364 10249 24404 10289
rect 24556 10228 24596 10268
rect 24748 10228 24788 10268
rect 25420 10228 25460 10268
rect 30220 10228 30260 10268
rect 30412 10228 30452 10268
rect 30604 10228 30644 10268
rect 30796 10228 30836 10268
rect 30988 10228 31028 10268
rect 31180 10249 31220 10289
rect 31372 10228 31412 10268
rect 31564 10228 31604 10268
rect 32044 10228 32084 10268
rect 35596 10228 35636 10268
rect 35788 10228 35828 10268
rect 35980 10228 36020 10268
rect 36172 10228 36212 10268
rect 36364 10228 36404 10268
rect 36556 10228 36596 10268
rect 36748 10228 36788 10268
rect 36940 10228 36980 10268
rect 37420 10228 37460 10268
rect 37612 10228 37652 10268
rect 37804 10228 37844 10268
rect 37996 10228 38036 10268
rect 38188 10228 38228 10268
rect 38380 10228 38420 10268
rect 38572 10228 38612 10268
rect 38764 10228 38804 10268
rect 38956 10228 38996 10268
rect 39148 10228 39188 10268
rect 40588 10228 40628 10268
rect 41548 10228 41588 10268
rect 41836 10228 41876 10268
rect 42796 10228 42836 10268
rect 50284 10228 50324 10268
rect 52108 10228 52148 10268
rect 53068 10228 53108 10268
rect 57580 10228 57620 10268
rect 57772 10228 57812 10268
rect 58156 10228 58196 10268
rect 58618 10228 58658 10268
rect 58924 10228 58964 10268
rect 59116 10228 59156 10268
rect 59884 10228 59924 10268
rect 60076 10228 60116 10268
rect 60268 10228 60308 10268
rect 60460 10228 60500 10268
rect 68428 10228 68468 10268
rect 69580 10228 69620 10268
rect 69772 10228 69812 10268
rect 71308 10228 71348 10268
rect 71500 10228 71540 10268
rect 72940 10228 72980 10268
rect 73132 10228 73172 10268
rect 73324 10228 73364 10268
rect 73516 10228 73556 10268
rect 73804 10228 73844 10268
rect 73996 10228 74036 10268
rect 74284 10228 74324 10268
rect 74476 10228 74516 10268
rect 76492 10228 76532 10268
rect 76684 10228 76724 10268
rect 76876 10228 76916 10268
rect 77068 10228 77108 10268
rect 77260 10228 77300 10268
rect 77452 10228 77492 10268
rect 77644 10228 77684 10268
rect 77836 10228 77876 10268
rect 82540 10228 82580 10268
rect 82732 10228 82772 10268
rect 83212 10228 83252 10268
rect 83404 10228 83444 10268
rect 83596 10228 83636 10268
rect 83788 10228 83828 10268
rect 83980 10228 84020 10268
rect 84172 10228 84212 10268
rect 87820 10228 87860 10268
rect 88012 10228 88052 10268
rect 88204 10228 88244 10268
rect 88396 10228 88436 10268
rect 88588 10228 88628 10268
rect 88684 10228 88724 10268
rect 88780 10228 88820 10268
rect 88963 10213 89003 10253
rect 89164 10228 89204 10268
rect 89452 10228 89492 10268
rect 89644 10228 89684 10268
rect 12844 10144 12884 10184
rect 21484 10144 21524 10184
rect 25228 10144 25268 10184
rect 32236 10144 32276 10184
rect 15436 10060 15476 10100
rect 16204 10060 16244 10100
rect 21580 10060 21620 10100
rect 25324 10060 25364 10100
rect 30316 10060 30356 10100
rect 30700 10060 30740 10100
rect 37900 10060 37940 10100
rect 58156 10060 58196 10100
rect 58444 10060 58484 10100
rect 58636 10060 58676 10100
rect 60076 10060 60116 10100
rect 69100 10060 69140 10100
rect 74380 10060 74420 10100
rect 87916 10060 87956 10100
rect 89068 10060 89108 10100
rect 11308 9976 11348 10016
rect 11692 9976 11732 10016
rect 12076 9976 12116 10016
rect 12460 9976 12500 10016
rect 14668 9976 14708 10016
rect 15052 9976 15092 10016
rect 15820 9976 15860 10016
rect 18700 9976 18740 10016
rect 19468 9976 19508 10016
rect 20236 9976 20276 10016
rect 24268 9976 24308 10016
rect 24652 9976 24692 10016
rect 31084 9976 31124 10016
rect 31468 9976 31508 10016
rect 32044 9976 32084 10016
rect 35692 9976 35732 10016
rect 36844 9976 36884 10016
rect 37516 9976 37556 10016
rect 38284 9976 38324 10016
rect 38668 9976 38708 10016
rect 39052 9976 39092 10016
rect 57964 9976 58004 10016
rect 59116 9976 59156 10016
rect 60460 9976 60500 10016
rect 71404 9976 71444 10016
rect 73036 9976 73076 10016
rect 76588 9976 76628 10016
rect 76972 9976 77012 10016
rect 77356 9976 77396 10016
rect 77740 9976 77780 10016
rect 82636 9976 82676 10016
rect 83308 9976 83348 10016
rect 83692 9976 83732 10016
rect 89548 9976 89588 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 64168 9808 64208 9848
rect 64250 9808 64290 9848
rect 64332 9808 64372 9848
rect 64414 9808 64454 9848
rect 64496 9808 64536 9848
rect 79288 9808 79328 9848
rect 79370 9808 79410 9848
rect 79452 9808 79492 9848
rect 79534 9808 79574 9848
rect 79616 9808 79656 9848
rect 94408 9808 94448 9848
rect 94490 9808 94530 9848
rect 94572 9808 94612 9848
rect 94654 9808 94694 9848
rect 94736 9808 94776 9848
rect 34540 9640 34580 9680
rect 56236 9640 56276 9680
rect 56620 9640 56660 9680
rect 73804 9640 73844 9680
rect 77452 9640 77492 9680
rect 36364 9556 36404 9596
rect 48460 9556 48500 9596
rect 48652 9556 48692 9596
rect 51148 9556 51188 9596
rect 52300 9556 52340 9596
rect 55852 9556 55892 9596
rect 58732 9556 58772 9596
rect 59884 9556 59924 9596
rect 60364 9556 60404 9596
rect 60844 9556 60884 9596
rect 72076 9556 72116 9596
rect 40684 9472 40724 9512
rect 48268 9472 48308 9512
rect 49804 9472 49844 9512
rect 11596 9388 11636 9428
rect 11788 9388 11828 9428
rect 12076 9388 12116 9428
rect 12268 9388 12308 9428
rect 14572 9388 14612 9428
rect 14668 9388 14708 9428
rect 14764 9388 14804 9428
rect 14956 9388 14996 9428
rect 15148 9388 15188 9428
rect 15340 9388 15380 9428
rect 15532 9388 15572 9428
rect 15724 9388 15764 9428
rect 15916 9388 15956 9428
rect 16108 9388 16148 9428
rect 16300 9388 16340 9428
rect 18988 9388 19028 9428
rect 19180 9388 19220 9428
rect 19372 9388 19412 9428
rect 19564 9388 19604 9428
rect 19756 9388 19796 9428
rect 19948 9388 19988 9428
rect 24172 9388 24212 9428
rect 24364 9388 24404 9428
rect 24556 9388 24596 9428
rect 24748 9388 24788 9428
rect 25228 9388 25268 9428
rect 25420 9388 25460 9428
rect 30028 9388 30068 9428
rect 30220 9388 30260 9428
rect 30604 9388 30644 9428
rect 30796 9388 30836 9428
rect 30988 9375 31028 9415
rect 31084 9388 31124 9428
rect 31180 9388 31220 9428
rect 34444 9388 34484 9428
rect 34636 9388 34676 9428
rect 34828 9388 34868 9428
rect 35020 9388 35060 9428
rect 36268 9388 36308 9428
rect 36460 9388 36500 9428
rect 36652 9388 36692 9428
rect 36844 9388 36884 9428
rect 37132 9388 37172 9428
rect 37324 9388 37364 9428
rect 37996 9388 38036 9428
rect 38188 9388 38228 9428
rect 38380 9388 38420 9428
rect 38572 9388 38612 9428
rect 38764 9388 38804 9428
rect 38956 9388 38996 9428
rect 39340 9388 39380 9428
rect 40300 9388 40340 9428
rect 41548 9388 41588 9428
rect 42316 9388 42356 9428
rect 43276 9388 43316 9428
rect 48844 9388 48884 9428
rect 48940 9388 48980 9428
rect 49516 9388 49556 9428
rect 49612 9388 49652 9428
rect 51340 9388 51380 9428
rect 51436 9388 51476 9428
rect 52012 9388 52052 9428
rect 52108 9388 52148 9428
rect 52492 9388 52532 9428
rect 53452 9388 53492 9428
rect 54796 9388 54836 9428
rect 54988 9388 55028 9428
rect 55756 9388 55796 9428
rect 55948 9388 55988 9428
rect 56140 9388 56180 9428
rect 56332 9388 56372 9428
rect 56524 9388 56564 9428
rect 56716 9388 56756 9428
rect 58732 9388 58772 9428
rect 59020 9388 59060 9428
rect 59212 9388 59252 9428
rect 59404 9388 59444 9428
rect 59596 9388 59636 9428
rect 59884 9388 59924 9428
rect 60364 9388 60404 9428
rect 60844 9388 60884 9428
rect 62092 9388 62132 9428
rect 65164 9388 65204 9428
rect 66124 9388 66164 9428
rect 70540 9388 70580 9428
rect 70732 9388 70772 9428
rect 71596 9388 71636 9428
rect 71788 9388 71828 9428
rect 71980 9388 72020 9428
rect 72172 9388 72212 9428
rect 73132 9388 73172 9428
rect 73324 9388 73364 9428
rect 73708 9388 73748 9428
rect 73900 9388 73940 9428
rect 76972 9388 77012 9428
rect 77164 9388 77204 9428
rect 77356 9388 77396 9428
rect 77548 9388 77588 9428
rect 77740 9388 77780 9428
rect 77932 9388 77972 9428
rect 78316 9388 78356 9428
rect 78508 9388 78548 9428
rect 79276 9388 79316 9428
rect 80236 9388 80276 9428
rect 80620 9388 80660 9428
rect 80812 9388 80852 9428
rect 81004 9388 81044 9428
rect 81196 9388 81236 9428
rect 81868 9388 81908 9428
rect 82060 9388 82100 9428
rect 87148 9388 87188 9428
rect 87340 9388 87380 9428
rect 87724 9388 87764 9428
rect 87820 9388 87860 9428
rect 87916 9388 87956 9428
rect 88204 9388 88244 9428
rect 88396 9388 88436 9428
rect 88588 9388 88628 9428
rect 88780 9388 88820 9428
rect 88972 9388 89012 9428
rect 89164 9388 89204 9428
rect 89356 9388 89396 9428
rect 89548 9388 89588 9428
rect 89740 9388 89780 9428
rect 89932 9388 89972 9428
rect 11692 9304 11732 9344
rect 15052 9304 15092 9344
rect 15436 9304 15476 9344
rect 15820 9304 15860 9344
rect 16204 9304 16244 9344
rect 19084 9304 19124 9344
rect 19468 9304 19508 9344
rect 19852 9304 19892 9344
rect 24268 9304 24308 9344
rect 24652 9304 24692 9344
rect 30700 9304 30740 9344
rect 34924 9304 34964 9344
rect 36748 9304 36788 9344
rect 38092 9304 38132 9344
rect 38476 9304 38516 9344
rect 38860 9304 38900 9344
rect 54892 9304 54932 9344
rect 62956 9304 62996 9344
rect 71692 9304 71732 9344
rect 73228 9304 73268 9344
rect 77068 9304 77108 9344
rect 77836 9304 77876 9344
rect 78412 9304 78452 9344
rect 80716 9304 80756 9344
rect 81100 9304 81140 9344
rect 81964 9304 82004 9344
rect 87244 9304 87284 9344
rect 88300 9304 88340 9344
rect 88684 9304 88724 9344
rect 89068 9304 89108 9344
rect 89452 9304 89492 9344
rect 89836 9304 89876 9344
rect 48940 9220 48980 9260
rect 49516 9220 49556 9260
rect 51436 9220 51476 9260
rect 52012 9220 52052 9260
rect 58540 9220 58580 9260
rect 59116 9220 59156 9260
rect 59500 9220 59540 9260
rect 60076 9220 60116 9260
rect 60556 9220 60596 9260
rect 61036 9220 61076 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 65408 9052 65448 9092
rect 65490 9052 65530 9092
rect 65572 9052 65612 9092
rect 65654 9052 65694 9092
rect 65736 9052 65776 9092
rect 80528 9052 80568 9092
rect 80610 9052 80650 9092
rect 80692 9052 80732 9092
rect 80774 9052 80814 9092
rect 80856 9052 80896 9092
rect 95648 9052 95688 9092
rect 95730 9052 95770 9092
rect 95812 9052 95852 9092
rect 95894 9052 95934 9092
rect 95976 9052 96016 9092
rect 15340 8884 15380 8924
rect 31948 8884 31988 8924
rect 45196 8884 45236 8924
rect 49324 8884 49364 8924
rect 49900 8884 49940 8924
rect 52588 8884 52628 8924
rect 55468 8884 55508 8924
rect 58732 8884 58772 8924
rect 9772 8800 9812 8840
rect 11596 8800 11636 8840
rect 11980 8800 12020 8840
rect 12364 8800 12404 8840
rect 18700 8800 18740 8840
rect 25036 8800 25076 8840
rect 27916 8800 27956 8840
rect 28300 8800 28340 8840
rect 28684 8800 28724 8840
rect 34828 8800 34868 8840
rect 50188 8800 50228 8840
rect 70060 8800 70100 8840
rect 70540 8800 70580 8840
rect 70924 8800 70964 8840
rect 74668 8800 74708 8840
rect 75052 8800 75092 8840
rect 75436 8800 75476 8840
rect 78796 8800 78836 8840
rect 80908 8800 80948 8840
rect 81676 8800 81716 8840
rect 82060 8800 82100 8840
rect 83212 8800 83252 8840
rect 83596 8800 83636 8840
rect 86956 8800 86996 8840
rect 87724 8800 87764 8840
rect 89068 8800 89108 8840
rect 9676 8716 9716 8756
rect 9868 8716 9908 8756
rect 10060 8716 10100 8756
rect 10252 8716 10292 8756
rect 11116 8716 11156 8756
rect 11308 8716 11348 8756
rect 11500 8716 11540 8756
rect 11692 8716 11732 8756
rect 11884 8716 11924 8756
rect 12076 8716 12116 8756
rect 12268 8716 12308 8756
rect 12460 8716 12500 8756
rect 15724 8716 15764 8756
rect 18604 8716 18644 8756
rect 18796 8716 18836 8756
rect 20620 8716 20660 8756
rect 20812 8716 20852 8756
rect 24172 8716 24212 8756
rect 24364 8716 24404 8756
rect 24556 8716 24596 8756
rect 24748 8716 24788 8756
rect 24940 8716 24980 8756
rect 25132 8716 25172 8756
rect 25420 8716 25460 8756
rect 25612 8716 25652 8756
rect 27436 8716 27476 8756
rect 27628 8716 27668 8756
rect 27820 8716 27860 8756
rect 28012 8716 28052 8756
rect 28204 8716 28244 8756
rect 28396 8716 28436 8756
rect 28588 8716 28628 8756
rect 28780 8716 28820 8756
rect 29356 8716 29396 8756
rect 29548 8716 29588 8756
rect 32332 8716 32372 8756
rect 33964 8716 34004 8756
rect 34156 8716 34196 8756
rect 34348 8716 34388 8756
rect 34540 8716 34580 8756
rect 34732 8716 34772 8756
rect 34924 8716 34964 8756
rect 35116 8716 35156 8756
rect 35308 8716 35348 8756
rect 35500 8716 35540 8756
rect 35692 8716 35732 8756
rect 37036 8716 37076 8756
rect 37228 8716 37268 8756
rect 38284 8716 38324 8756
rect 38476 8716 38516 8756
rect 43372 8716 43412 8756
rect 43660 8716 43700 8756
rect 44620 8716 44660 8756
rect 44908 8716 44948 8756
rect 45100 8716 45140 8756
rect 45196 8716 45236 8756
rect 46156 8716 46196 8756
rect 47116 8716 47156 8756
rect 48364 8716 48404 8756
rect 49324 8716 49364 8756
rect 49420 8716 49460 8756
rect 49612 8716 49652 8756
rect 49996 8716 50036 8756
rect 50476 8716 50516 8756
rect 52588 8716 52628 8756
rect 52684 8716 52724 8756
rect 52876 8716 52916 8756
rect 54316 8716 54356 8756
rect 54508 8716 54548 8756
rect 54892 8724 54932 8764
rect 55276 8716 55316 8756
rect 55948 8716 55988 8756
rect 56140 8716 56180 8756
rect 56812 8724 56852 8764
rect 57196 8724 57236 8764
rect 59212 8716 59252 8756
rect 60076 8716 60116 8756
rect 66988 8716 67028 8756
rect 67180 8716 67220 8756
rect 69964 8716 70004 8756
rect 70156 8716 70196 8756
rect 70444 8716 70484 8756
rect 70636 8716 70676 8756
rect 70828 8716 70868 8756
rect 71020 8716 71060 8756
rect 73228 8716 73268 8756
rect 73420 8716 73460 8756
rect 74572 8716 74612 8756
rect 74764 8716 74804 8756
rect 74956 8716 74996 8756
rect 75148 8716 75188 8756
rect 75340 8716 75380 8756
rect 75532 8716 75572 8756
rect 75916 8716 75956 8756
rect 76108 8716 76148 8756
rect 76684 8716 76724 8756
rect 76876 8716 76916 8756
rect 77932 8716 77972 8756
rect 78124 8716 78164 8756
rect 78316 8729 78356 8769
rect 78508 8716 78548 8756
rect 78700 8716 78740 8756
rect 78892 8716 78932 8756
rect 80812 8716 80852 8756
rect 81004 8716 81044 8756
rect 81196 8716 81236 8756
rect 81292 8716 81332 8756
rect 81388 8716 81428 8756
rect 81580 8716 81620 8756
rect 81772 8716 81812 8756
rect 81964 8716 82004 8756
rect 82156 8716 82196 8756
rect 83116 8716 83156 8756
rect 83308 8716 83348 8756
rect 83500 8716 83540 8756
rect 83692 8716 83732 8756
rect 84076 8716 84116 8756
rect 84268 8716 84308 8756
rect 86860 8716 86900 8756
rect 87052 8716 87092 8756
rect 87244 8716 87284 8756
rect 87436 8716 87476 8756
rect 87628 8716 87668 8756
rect 87820 8716 87860 8756
rect 88012 8716 88052 8756
rect 88204 8729 88244 8769
rect 88972 8716 89012 8756
rect 89164 8716 89204 8756
rect 89356 8716 89396 8756
rect 89548 8716 89588 8756
rect 34060 8632 34100 8672
rect 42508 8632 42548 8672
rect 48748 8632 48788 8672
rect 54412 8632 54452 8672
rect 58924 8632 58964 8672
rect 48076 8548 48116 8588
rect 48940 8548 48980 8588
rect 54892 8548 54932 8588
rect 55276 8548 55316 8588
rect 56044 8548 56084 8588
rect 56620 8548 56660 8588
rect 56812 8548 56852 8588
rect 57196 8548 57236 8588
rect 84172 8548 84212 8588
rect 10156 8464 10196 8504
rect 11212 8464 11252 8504
rect 24268 8464 24308 8504
rect 24652 8464 24692 8504
rect 27532 8464 27572 8504
rect 34444 8464 34484 8504
rect 35212 8464 35252 8504
rect 35596 8464 35636 8504
rect 50956 8464 50996 8504
rect 54700 8464 54740 8504
rect 57388 8464 57428 8504
rect 73324 8464 73364 8504
rect 76780 8464 76820 8504
rect 78028 8464 78068 8504
rect 78412 8464 78452 8504
rect 87340 8464 87380 8504
rect 88108 8464 88148 8504
rect 89452 8464 89492 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 64168 8296 64208 8336
rect 64250 8296 64290 8336
rect 64332 8296 64372 8336
rect 64414 8296 64454 8336
rect 64496 8296 64536 8336
rect 79288 8296 79328 8336
rect 79370 8296 79410 8336
rect 79452 8296 79492 8336
rect 79534 8296 79574 8336
rect 79616 8296 79656 8336
rect 94408 8296 94448 8336
rect 94490 8296 94530 8336
rect 94572 8296 94612 8336
rect 94654 8296 94694 8336
rect 94736 8296 94776 8336
rect 30220 8128 30260 8168
rect 37036 8128 37076 8168
rect 50764 8128 50804 8168
rect 54604 8128 54644 8168
rect 58732 8128 58772 8168
rect 60172 8128 60212 8168
rect 72556 8128 72596 8168
rect 75052 8128 75092 8168
rect 81580 8128 81620 8168
rect 83692 8128 83732 8168
rect 86956 8128 86996 8168
rect 12460 8044 12500 8084
rect 22348 8044 22388 8084
rect 37708 8044 37748 8084
rect 46252 8044 46292 8084
rect 48172 8044 48212 8084
rect 51436 8044 51476 8084
rect 58924 8044 58964 8084
rect 85228 8044 85268 8084
rect 16300 7960 16340 8000
rect 32428 7960 32468 8000
rect 34924 7960 34964 8000
rect 35308 7960 35348 8000
rect 45580 7960 45620 8000
rect 50572 7960 50612 8000
rect 54412 7960 54452 8000
rect 58348 7960 58388 8000
rect 59980 7960 60020 8000
rect 84844 7960 84884 8000
rect 87532 7960 87572 8000
rect 8908 7876 8948 7916
rect 9100 7876 9140 7916
rect 9292 7876 9332 7916
rect 9484 7876 9524 7916
rect 9676 7876 9716 7916
rect 9868 7876 9908 7916
rect 10060 7876 10100 7916
rect 10252 7876 10292 7916
rect 10444 7876 10484 7916
rect 10636 7876 10676 7916
rect 11596 7876 11636 7916
rect 11788 7876 11828 7916
rect 11980 7876 12020 7916
rect 12172 7876 12212 7916
rect 12364 7876 12404 7916
rect 12556 7876 12596 7916
rect 12748 7876 12788 7916
rect 12940 7876 12980 7916
rect 13132 7876 13172 7916
rect 13324 7876 13364 7916
rect 13516 7876 13556 7916
rect 13708 7876 13748 7916
rect 14188 7876 14228 7916
rect 14380 7876 14420 7916
rect 17164 7876 17204 7916
rect 17836 7876 17876 7916
rect 18028 7876 18068 7916
rect 18220 7876 18260 7916
rect 18412 7876 18452 7916
rect 18604 7876 18644 7916
rect 18796 7876 18836 7916
rect 18988 7876 19028 7916
rect 19180 7876 19220 7916
rect 19372 7876 19412 7916
rect 19564 7876 19604 7916
rect 19756 7876 19796 7916
rect 19948 7863 19988 7903
rect 20428 7876 20468 7916
rect 20620 7876 20660 7916
rect 22540 7876 22580 7916
rect 22636 7876 22676 7916
rect 23212 7876 23252 7916
rect 23308 7876 23348 7916
rect 24556 7876 24596 7916
rect 24748 7876 24788 7916
rect 24940 7876 24980 7916
rect 25132 7876 25172 7916
rect 25324 7876 25364 7916
rect 25516 7876 25556 7916
rect 25708 7876 25748 7916
rect 25900 7876 25940 7916
rect 27628 7876 27668 7916
rect 27820 7876 27860 7916
rect 28012 7876 28052 7916
rect 28204 7876 28244 7916
rect 28396 7876 28436 7916
rect 28588 7876 28628 7916
rect 28780 7876 28820 7916
rect 28972 7876 29012 7916
rect 29932 7876 29972 7916
rect 30028 7876 30068 7916
rect 30796 7876 30836 7916
rect 30988 7876 31028 7916
rect 31180 7876 31220 7916
rect 31372 7876 31412 7916
rect 31564 7876 31604 7916
rect 31756 7876 31796 7916
rect 31948 7876 31988 7916
rect 32140 7876 32180 7916
rect 32332 7876 32372 7916
rect 32524 7876 32564 7916
rect 32716 7876 32756 7916
rect 32812 7876 32852 7916
rect 32908 7876 32948 7916
rect 33100 7876 33140 7916
rect 33196 7876 33236 7916
rect 33292 7876 33332 7916
rect 33580 7876 33620 7916
rect 33772 7876 33812 7916
rect 34444 7876 34484 7916
rect 34636 7876 34676 7916
rect 34828 7876 34868 7916
rect 35020 7876 35060 7916
rect 36172 7876 36212 7916
rect 36748 7876 36788 7916
rect 37420 7876 37460 7916
rect 9004 7792 9044 7832
rect 9388 7792 9428 7832
rect 9772 7792 9812 7832
rect 10156 7792 10196 7832
rect 10540 7792 10580 7832
rect 11692 7792 11732 7832
rect 12076 7792 12116 7832
rect 12844 7792 12884 7832
rect 13228 7792 13268 7832
rect 13612 7792 13652 7832
rect 17932 7792 17972 7832
rect 18316 7792 18356 7832
rect 18700 7792 18740 7832
rect 19084 7792 19124 7832
rect 19468 7792 19508 7832
rect 19852 7792 19892 7832
rect 23020 7792 23060 7832
rect 24652 7792 24692 7832
rect 25036 7792 25076 7832
rect 25420 7792 25460 7832
rect 25804 7792 25844 7832
rect 27724 7792 27764 7832
rect 28108 7792 28148 7832
rect 28492 7792 28532 7832
rect 28876 7792 28916 7832
rect 30892 7792 30932 7832
rect 31276 7792 31316 7832
rect 31660 7792 31700 7832
rect 32044 7792 32084 7832
rect 36844 7834 36884 7874
rect 37516 7876 37556 7916
rect 39436 7876 39476 7916
rect 39532 7876 39572 7916
rect 39724 7876 39764 7916
rect 39916 7876 39956 7916
rect 40876 7876 40916 7916
rect 41164 7876 41204 7916
rect 42028 7876 42068 7916
rect 42412 7876 42452 7916
rect 43372 7876 43412 7916
rect 44044 7876 44084 7916
rect 44236 7876 44276 7916
rect 44332 7876 44372 7916
rect 44908 7876 44948 7916
rect 45004 7876 45044 7916
rect 45196 7876 45236 7916
rect 45772 7876 45812 7916
rect 45868 7876 45908 7916
rect 46444 7876 46484 7916
rect 46540 7876 46580 7916
rect 46924 7876 46964 7916
rect 47116 7876 47156 7916
rect 47212 7876 47252 7916
rect 48364 7876 48404 7916
rect 48460 7876 48500 7916
rect 49228 7876 49268 7916
rect 50188 7876 50228 7916
rect 51244 7876 51284 7916
rect 51436 7876 51476 7916
rect 51628 7876 51668 7916
rect 51820 7876 51860 7916
rect 54796 7876 54836 7916
rect 54988 7876 55028 7916
rect 56044 7876 56084 7916
rect 56140 7876 56180 7916
rect 56236 7876 56276 7916
rect 56428 7876 56468 7916
rect 56620 7876 56660 7916
rect 56812 7876 56852 7916
rect 57004 7876 57044 7916
rect 57676 7876 57716 7916
rect 57868 7876 57908 7916
rect 58252 7876 58292 7916
rect 58444 7876 58484 7916
rect 58924 7876 58964 7916
rect 59500 7876 59540 7916
rect 59692 7876 59732 7916
rect 62668 7876 62708 7916
rect 63628 7876 63668 7916
rect 64012 7876 64052 7916
rect 64972 7876 65012 7916
rect 65260 7876 65300 7916
rect 66220 7876 66260 7916
rect 67180 7876 67220 7916
rect 67372 7876 67412 7916
rect 67660 7876 67700 7916
rect 67852 7876 67892 7916
rect 68716 7876 68756 7916
rect 68908 7876 68948 7916
rect 69772 7876 69812 7916
rect 69964 7876 70004 7916
rect 70156 7876 70196 7916
rect 70348 7876 70388 7916
rect 70540 7876 70580 7916
rect 70732 7876 70772 7916
rect 70924 7876 70964 7916
rect 71116 7876 71156 7916
rect 71692 7876 71732 7916
rect 71884 7876 71924 7916
rect 72076 7876 72116 7916
rect 72268 7876 72308 7916
rect 72748 7876 72788 7916
rect 73996 7876 74036 7916
rect 74188 7876 74228 7916
rect 74380 7876 74420 7916
rect 74572 7876 74612 7916
rect 74860 7876 74900 7916
rect 75244 7876 75284 7916
rect 75436 7876 75476 7916
rect 75724 7876 75764 7916
rect 75916 7876 75956 7916
rect 77548 7876 77588 7916
rect 77740 7876 77780 7916
rect 77932 7876 77972 7916
rect 78124 7876 78164 7916
rect 78412 7876 78452 7916
rect 78604 7876 78644 7916
rect 78796 7876 78836 7916
rect 78988 7876 79028 7916
rect 80716 7876 80756 7916
rect 80908 7876 80948 7916
rect 81100 7876 81140 7916
rect 81292 7876 81332 7916
rect 81484 7876 81524 7916
rect 81676 7876 81716 7916
rect 81868 7876 81908 7916
rect 82060 7876 82100 7916
rect 82444 7899 82484 7939
rect 82636 7876 82676 7916
rect 82828 7876 82868 7916
rect 83020 7876 83060 7916
rect 83212 7876 83252 7916
rect 83404 7876 83444 7916
rect 83596 7876 83636 7916
rect 83788 7876 83828 7916
rect 83980 7876 84020 7916
rect 84172 7876 84212 7916
rect 84364 7876 84404 7916
rect 84556 7876 84596 7916
rect 84748 7876 84788 7916
rect 84940 7876 84980 7916
rect 85132 7876 85172 7916
rect 85324 7876 85364 7916
rect 86764 7876 86804 7916
rect 87820 7876 87860 7916
rect 88012 7876 88052 7916
rect 88204 7876 88244 7916
rect 88396 7876 88436 7916
rect 88588 7876 88628 7916
rect 88684 7876 88724 7916
rect 88789 7863 88829 7903
rect 89068 7876 89108 7916
rect 89263 7899 89303 7939
rect 89452 7863 89492 7903
rect 89644 7876 89684 7916
rect 34540 7792 34580 7832
rect 49420 7792 49460 7832
rect 49996 7792 50036 7832
rect 69868 7792 69908 7832
rect 70252 7792 70292 7832
rect 70636 7792 70676 7832
rect 71020 7792 71060 7832
rect 74092 7792 74132 7832
rect 74476 7792 74516 7832
rect 75820 7792 75860 7832
rect 77644 7792 77684 7832
rect 78028 7792 78068 7832
rect 78892 7792 78932 7832
rect 80812 7792 80852 7832
rect 81196 7792 81236 7832
rect 81964 7792 82004 7832
rect 82540 7792 82580 7832
rect 82924 7792 82964 7832
rect 83308 7792 83348 7832
rect 84076 7792 84116 7832
rect 84460 7792 84500 7832
rect 87916 7792 87956 7832
rect 88300 7792 88340 7832
rect 89164 7792 89204 7832
rect 89548 7792 89588 7832
rect 22636 7708 22676 7748
rect 23308 7708 23348 7748
rect 36748 7708 36788 7748
rect 37420 7708 37460 7748
rect 39724 7708 39764 7748
rect 29740 7666 29780 7706
rect 44524 7666 44564 7706
rect 45868 7708 45908 7748
rect 46540 7708 46580 7748
rect 47212 7708 47252 7748
rect 48460 7708 48500 7748
rect 49612 7708 49652 7748
rect 44716 7666 44756 7706
rect 49804 7666 49844 7706
rect 54604 7708 54644 7748
rect 54892 7708 54932 7748
rect 56524 7708 56564 7748
rect 56908 7708 56948 7748
rect 57772 7708 57812 7748
rect 72844 7708 72884 7748
rect 74764 7708 74804 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 65408 7540 65448 7580
rect 65490 7540 65530 7580
rect 65572 7540 65612 7580
rect 65654 7540 65694 7580
rect 65736 7540 65776 7580
rect 80528 7540 80568 7580
rect 80610 7540 80650 7580
rect 80692 7540 80732 7580
rect 80774 7540 80814 7580
rect 80856 7540 80896 7580
rect 95648 7540 95688 7580
rect 95730 7540 95770 7580
rect 95812 7540 95852 7580
rect 95894 7540 95934 7580
rect 95976 7540 96016 7580
rect 23020 7372 23060 7412
rect 36652 7372 36692 7412
rect 42988 7372 43028 7412
rect 44620 7372 44660 7412
rect 46636 7372 46676 7412
rect 51340 7372 51380 7412
rect 59788 7372 59828 7412
rect 60556 7372 60596 7412
rect 77068 7414 77108 7454
rect 60844 7372 60884 7412
rect 61804 7372 61844 7412
rect 62092 7372 62132 7412
rect 78412 7372 78452 7412
rect 78892 7372 78932 7412
rect 79180 7372 79220 7412
rect 86860 7372 86900 7412
rect 89068 7372 89108 7412
rect 60460 7288 60500 7328
rect 78700 7288 78740 7328
rect 85708 7288 85748 7328
rect 9676 7204 9716 7244
rect 9868 7204 9908 7244
rect 10060 7204 10100 7244
rect 10252 7204 10292 7244
rect 10636 7204 10676 7244
rect 10828 7217 10868 7257
rect 11020 7204 11060 7244
rect 11212 7204 11252 7244
rect 11884 7204 11924 7244
rect 12076 7204 12116 7244
rect 12556 7204 12596 7244
rect 12748 7204 12788 7244
rect 13420 7204 13460 7244
rect 13612 7204 13652 7244
rect 18700 7204 18740 7244
rect 18892 7204 18932 7244
rect 22732 7204 22772 7244
rect 22924 7204 22964 7244
rect 23020 7204 23060 7244
rect 23980 7204 24020 7244
rect 24172 7204 24212 7244
rect 24364 7204 24404 7244
rect 24556 7204 24596 7244
rect 25036 7204 25076 7244
rect 25132 7204 25172 7244
rect 25228 7204 25268 7244
rect 26956 7204 26996 7244
rect 27148 7204 27188 7244
rect 30028 7204 30068 7244
rect 31180 7204 31220 7244
rect 31660 7204 31700 7244
rect 31860 7203 31900 7243
rect 32332 7204 32372 7244
rect 32620 7204 32660 7244
rect 32812 7204 32852 7244
rect 33868 7204 33908 7244
rect 34060 7204 34100 7244
rect 34252 7204 34292 7244
rect 34444 7204 34484 7244
rect 37324 7204 37364 7244
rect 37516 7204 37556 7244
rect 37708 7204 37748 7244
rect 37900 7204 37940 7244
rect 39148 7204 39188 7244
rect 40108 7204 40148 7244
rect 40396 7204 40436 7244
rect 41356 7204 41396 7244
rect 43468 7204 43508 7244
rect 44332 7204 44372 7244
rect 44524 7205 44564 7245
rect 44620 7204 44660 7244
rect 45772 7204 45812 7244
rect 45964 7204 46004 7244
rect 46540 7204 46580 7244
rect 46636 7204 46676 7244
rect 47116 7204 47156 7244
rect 47308 7204 47348 7244
rect 48556 7204 48596 7244
rect 48748 7204 48788 7244
rect 49036 7204 49076 7244
rect 49228 7204 49268 7244
rect 49324 7204 49364 7244
rect 49516 7204 49556 7244
rect 49708 7204 49748 7244
rect 50092 7204 50132 7244
rect 50380 7204 50420 7244
rect 50572 7204 50612 7244
rect 50764 7204 50804 7244
rect 50956 7204 50996 7244
rect 51244 7204 51284 7244
rect 51532 7204 51572 7244
rect 51724 7204 51764 7244
rect 51820 7204 51860 7244
rect 52012 7204 52052 7244
rect 52300 7204 52340 7244
rect 54316 7204 54356 7244
rect 54508 7204 54548 7244
rect 58348 7204 58388 7244
rect 59212 7204 59252 7244
rect 59404 7204 59444 7244
rect 59788 7204 59828 7244
rect 59980 7204 60020 7244
rect 60076 7204 60116 7244
rect 60268 7204 60308 7244
rect 60364 7204 60404 7244
rect 61900 7204 61940 7244
rect 63052 7204 63092 7244
rect 64012 7204 64052 7244
rect 64492 7204 64532 7244
rect 64684 7204 64724 7244
rect 64972 7204 65012 7244
rect 65164 7204 65204 7244
rect 66796 7204 66836 7244
rect 66988 7204 67028 7244
rect 68044 7204 68084 7244
rect 68236 7204 68276 7244
rect 68524 7204 68564 7244
rect 68716 7204 68756 7244
rect 69004 7204 69044 7244
rect 69196 7204 69236 7244
rect 70540 7225 70580 7265
rect 70732 7204 70772 7244
rect 74284 7204 74324 7244
rect 74476 7204 74516 7244
rect 74860 7204 74900 7244
rect 75052 7204 75092 7244
rect 75244 7204 75284 7244
rect 75436 7204 75476 7244
rect 77260 7204 77300 7244
rect 77356 7204 77396 7244
rect 77548 7204 77588 7244
rect 78028 7181 78068 7221
rect 78220 7204 78260 7244
rect 78508 7204 78548 7244
rect 78988 7204 79028 7244
rect 80812 7204 80852 7244
rect 81004 7204 81044 7244
rect 82636 7204 82676 7244
rect 82828 7204 82868 7244
rect 83020 7204 83060 7244
rect 83212 7204 83252 7244
rect 83404 7204 83444 7244
rect 83596 7204 83636 7244
rect 83788 7204 83828 7244
rect 83980 7204 84020 7244
rect 84172 7204 84212 7244
rect 84364 7204 84404 7244
rect 85612 7204 85652 7244
rect 85804 7204 85844 7244
rect 86380 7204 86420 7244
rect 87532 7204 87572 7244
rect 87724 7204 87764 7244
rect 88012 7204 88052 7244
rect 88204 7204 88244 7244
rect 89452 7204 89492 7244
rect 30412 7120 30452 7160
rect 33964 7120 34004 7160
rect 36460 7120 36500 7160
rect 46348 7120 46388 7160
rect 56236 7120 56276 7160
rect 56620 7120 56660 7160
rect 57196 7120 57236 7160
rect 61036 7120 61076 7160
rect 11980 7036 12020 7076
rect 29740 7036 29780 7076
rect 31852 7036 31892 7076
rect 32332 7036 32372 7076
rect 51820 7036 51860 7076
rect 58348 7036 58388 7076
rect 9772 6952 9812 6992
rect 10156 6952 10196 6992
rect 10732 6952 10772 6992
rect 11116 6952 11156 6992
rect 12652 6952 12692 6992
rect 18796 6952 18836 6992
rect 23980 6952 24020 6992
rect 24364 6952 24404 6992
rect 27148 6952 27188 6992
rect 32140 6952 32180 6992
rect 32716 6952 32756 6992
rect 34444 6952 34484 6992
rect 36652 6952 36692 6992
rect 37516 6952 37556 6992
rect 37900 6952 37940 6992
rect 49036 6952 49076 6992
rect 49516 6952 49556 6992
rect 52588 6952 52628 6992
rect 54412 6952 54452 6992
rect 56044 6952 56084 6992
rect 56428 6952 56468 6992
rect 57004 6952 57044 6992
rect 58540 6952 58580 6992
rect 60556 6952 60596 6992
rect 68236 6952 68276 6992
rect 68524 6952 68564 6992
rect 69004 6952 69044 6992
rect 70636 6952 70676 6992
rect 74476 6952 74516 6992
rect 74956 6952 74996 6992
rect 75340 6952 75380 6992
rect 78124 6952 78164 6992
rect 82828 6952 82868 6992
rect 83116 6952 83156 6992
rect 83500 6952 83540 6992
rect 83884 6952 83924 6992
rect 84268 6952 84308 6992
rect 88108 6952 88148 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 64168 6784 64208 6824
rect 64250 6784 64290 6824
rect 64332 6784 64372 6824
rect 64414 6784 64454 6824
rect 64496 6784 64536 6824
rect 79288 6784 79328 6824
rect 79370 6784 79410 6824
rect 79452 6784 79492 6824
rect 79534 6784 79574 6824
rect 79616 6784 79656 6824
rect 94408 6784 94448 6824
rect 94490 6784 94530 6824
rect 94572 6784 94612 6824
rect 94654 6784 94694 6824
rect 94736 6784 94776 6824
rect 15820 6616 15860 6656
rect 36652 6616 36692 6656
rect 48652 6616 48692 6656
rect 51436 6616 51476 6656
rect 51916 6616 51956 6656
rect 52108 6616 52148 6656
rect 52588 6616 52628 6656
rect 59308 6616 59348 6656
rect 62476 6616 62516 6656
rect 74188 6616 74228 6656
rect 77452 6616 77492 6656
rect 79468 6616 79508 6656
rect 87724 6616 87764 6656
rect 16396 6532 16436 6572
rect 18508 6532 18548 6572
rect 29932 6532 29972 6572
rect 32812 6532 32852 6572
rect 35500 6532 35540 6572
rect 35980 6532 36020 6572
rect 47884 6532 47924 6572
rect 49036 6532 49076 6572
rect 53260 6532 53300 6572
rect 54412 6532 54452 6572
rect 54988 6532 55028 6572
rect 57004 6532 57044 6572
rect 61228 6532 61268 6572
rect 62284 6532 62324 6572
rect 67276 6532 67316 6572
rect 71980 6532 72020 6572
rect 79276 6532 79316 6572
rect 79852 6532 79892 6572
rect 80236 6532 80276 6572
rect 82348 6532 82388 6572
rect 83308 6532 83348 6572
rect 1420 6448 1460 6488
rect 19468 6448 19508 6488
rect 20716 6448 20756 6488
rect 21100 6448 21140 6488
rect 35692 6448 35732 6488
rect 10444 6364 10484 6404
rect 10636 6364 10676 6404
rect 15628 6364 15668 6404
rect 15820 6364 15860 6404
rect 16012 6364 16052 6404
rect 16209 6361 16249 6401
rect 16396 6364 16436 6404
rect 16588 6364 16628 6404
rect 17740 6364 17780 6404
rect 17932 6364 17972 6404
rect 18124 6364 18164 6404
rect 18316 6364 18356 6404
rect 18508 6364 18548 6404
rect 18700 6364 18740 6404
rect 18892 6364 18932 6404
rect 19084 6364 19124 6404
rect 19660 6364 19700 6404
rect 19852 6364 19892 6404
rect 23212 6364 23252 6404
rect 23404 6364 23444 6404
rect 23596 6364 23636 6404
rect 24652 6406 24692 6446
rect 23788 6364 23828 6404
rect 24076 6364 24116 6404
rect 24268 6364 24308 6404
rect 24460 6364 24500 6404
rect 24748 6350 24788 6390
rect 24950 6365 24990 6405
rect 25132 6364 25172 6404
rect 25324 6364 25364 6404
rect 25516 6364 25556 6404
rect 26188 6364 26228 6404
rect 26380 6364 26420 6404
rect 26572 6364 26612 6404
rect 26764 6364 26804 6404
rect 26956 6364 26996 6404
rect 27148 6364 27188 6404
rect 27340 6364 27380 6404
rect 27532 6364 27572 6404
rect 27724 6364 27764 6404
rect 27916 6377 27956 6417
rect 28492 6364 28532 6404
rect 28684 6364 28724 6404
rect 29740 6364 29780 6404
rect 29932 6364 29972 6404
rect 30028 6364 30068 6404
rect 31468 6364 31508 6404
rect 31660 6364 31700 6404
rect 31852 6364 31892 6404
rect 32044 6364 32084 6404
rect 32236 6377 32276 6417
rect 32428 6364 32468 6404
rect 32620 6364 32660 6404
rect 32812 6364 32852 6404
rect 33196 6364 33236 6404
rect 33292 6364 33332 6404
rect 33676 6364 33716 6404
rect 33868 6364 33908 6404
rect 34060 6364 34100 6404
rect 34252 6364 34292 6404
rect 34444 6364 34484 6404
rect 34636 6353 34676 6393
rect 34828 6364 34868 6404
rect 35020 6364 35060 6404
rect 35884 6364 35924 6404
rect 37804 6406 37844 6446
rect 38764 6448 38804 6488
rect 46636 6448 46676 6488
rect 47212 6448 47252 6488
rect 47596 6448 47636 6488
rect 53068 6448 53108 6488
rect 57484 6448 57524 6488
rect 57964 6448 58004 6488
rect 58828 6448 58868 6488
rect 75724 6448 75764 6488
rect 78796 6448 78836 6488
rect 35980 6364 36020 6404
rect 36172 6364 36212 6404
rect 36364 6364 36404 6404
rect 37324 6364 37364 6404
rect 37612 6364 37652 6404
rect 37900 6364 37940 6404
rect 38092 6364 38132 6404
rect 38284 6364 38324 6404
rect 38668 6364 38708 6404
rect 38860 6364 38900 6404
rect 39340 6364 39380 6404
rect 40204 6364 40244 6404
rect 41644 6364 41684 6404
rect 41932 6364 41972 6404
rect 42796 6364 42836 6404
rect 43468 6364 43508 6404
rect 44332 6364 44372 6404
rect 44716 6364 44756 6404
rect 45676 6364 45716 6404
rect 46156 6364 46196 6404
rect 46348 6364 46388 6404
rect 47884 6364 47924 6404
rect 48076 6364 48116 6404
rect 48172 6364 48212 6404
rect 49324 6364 49364 6404
rect 50380 6364 50420 6404
rect 50668 6364 50708 6404
rect 50860 6364 50900 6404
rect 51148 6364 51188 6404
rect 51244 6364 51284 6404
rect 51436 6364 51476 6404
rect 51628 6364 51668 6404
rect 51916 6364 51956 6404
rect 52108 6350 52148 6390
rect 52300 6364 52340 6404
rect 52396 6364 52436 6404
rect 52588 6364 52628 6404
rect 52780 6364 52820 6404
rect 52876 6364 52916 6404
rect 53932 6364 53972 6404
rect 54124 6364 54164 6404
rect 54412 6364 54452 6404
rect 54988 6364 55028 6404
rect 55564 6364 55604 6404
rect 55756 6364 55796 6404
rect 56044 6364 56084 6404
rect 56236 6364 56276 6404
rect 56524 6364 56564 6404
rect 56716 6364 56756 6404
rect 57004 6364 57044 6404
rect 57388 6364 57428 6404
rect 57580 6364 57620 6404
rect 58252 6364 58292 6404
rect 58444 6364 58484 6404
rect 59884 6364 59924 6404
rect 60268 6364 60308 6404
rect 61036 6364 61076 6404
rect 61228 6364 61268 6404
rect 61804 6364 61844 6404
rect 61900 6364 61940 6404
rect 61996 6364 62036 6404
rect 62092 6364 62132 6404
rect 62668 6364 62708 6404
rect 62956 6364 62996 6404
rect 63148 6364 63188 6404
rect 64012 6364 64052 6404
rect 64972 6364 65012 6404
rect 65260 6364 65300 6404
rect 66220 6364 66260 6404
rect 66412 6364 66452 6404
rect 66604 6364 66644 6404
rect 67180 6364 67220 6404
rect 67372 6364 67412 6404
rect 67564 6364 67604 6404
rect 67756 6364 67796 6404
rect 68044 6364 68084 6404
rect 68236 6364 68276 6404
rect 68620 6364 68660 6404
rect 68812 6364 68852 6404
rect 69100 6364 69140 6404
rect 69292 6364 69332 6404
rect 69484 6364 69524 6404
rect 69676 6364 69716 6404
rect 71020 6364 71060 6404
rect 71788 6364 71828 6404
rect 71980 6364 72020 6404
rect 72652 6364 72692 6404
rect 72844 6364 72884 6404
rect 73228 6364 73268 6404
rect 73420 6364 73460 6404
rect 73996 6364 74036 6404
rect 74188 6364 74228 6404
rect 74373 6353 74413 6393
rect 74572 6364 74612 6404
rect 74764 6364 74804 6404
rect 74956 6364 74996 6404
rect 75148 6364 75188 6404
rect 75340 6364 75380 6404
rect 77452 6406 77492 6446
rect 79660 6448 79700 6488
rect 80044 6448 80084 6488
rect 80428 6448 80468 6488
rect 81964 6448 82004 6488
rect 83596 6448 83636 6488
rect 98476 6448 98516 6488
rect 76780 6364 76820 6404
rect 77644 6364 77684 6404
rect 77740 6364 77780 6404
rect 78700 6364 78740 6404
rect 78892 6364 78932 6404
rect 79084 6364 79124 6404
rect 79276 6364 79316 6404
rect 82156 6364 82196 6404
rect 82348 6364 82388 6404
rect 82732 6364 82772 6404
rect 82924 6364 82964 6404
rect 83116 6364 83156 6404
rect 83308 6364 83348 6404
rect 83500 6364 83540 6404
rect 83692 6364 83732 6404
rect 83884 6364 83924 6404
rect 84076 6364 84116 6404
rect 84652 6364 84692 6404
rect 86668 6364 86708 6404
rect 86860 6364 86900 6404
rect 87436 6364 87476 6404
rect 10540 6280 10580 6320
rect 16108 6280 16148 6320
rect 19756 6280 19796 6320
rect 27052 6280 27092 6320
rect 27436 6280 27476 6320
rect 27820 6280 27860 6320
rect 32332 6280 32372 6320
rect 34156 6280 34196 6320
rect 40780 6280 40820 6320
rect 50188 6280 50228 6320
rect 56140 6280 56180 6320
rect 56620 6280 56660 6320
rect 60556 6280 60596 6320
rect 63052 6280 63092 6320
rect 71308 6280 71348 6320
rect 72748 6280 72788 6320
rect 82828 6280 82868 6320
rect 83980 6280 84020 6320
rect 84844 6280 84884 6320
rect 86764 6280 86804 6320
rect 1228 6196 1268 6236
rect 17836 6196 17876 6236
rect 18220 6196 18260 6236
rect 18988 6196 19028 6236
rect 19276 6196 19316 6236
rect 20524 6196 20564 6236
rect 20908 6196 20948 6236
rect 23308 6196 23348 6236
rect 23692 6196 23732 6236
rect 24460 6196 24500 6236
rect 25036 6196 25076 6236
rect 25420 6196 25460 6236
rect 26284 6196 26324 6236
rect 26668 6196 26708 6236
rect 31564 6196 31604 6236
rect 31948 6196 31988 6236
rect 33004 6196 33044 6236
rect 33772 6196 33812 6236
rect 34540 6196 34580 6236
rect 34924 6196 34964 6236
rect 37612 6196 37652 6236
rect 38188 6196 38228 6236
rect 46828 6196 46868 6236
rect 47020 6196 47060 6236
rect 47404 6196 47444 6236
rect 47884 6196 47924 6236
rect 50476 6196 50516 6236
rect 51436 6196 51476 6236
rect 52588 6196 52628 6236
rect 54604 6196 54644 6236
rect 54796 6196 54836 6236
rect 57196 6196 57236 6236
rect 57772 6196 57812 6236
rect 58636 6196 58676 6236
rect 60748 6196 60788 6236
rect 62764 6196 62804 6236
rect 68140 6196 68180 6236
rect 69196 6196 69236 6236
rect 69580 6196 69620 6236
rect 71500 6196 71540 6236
rect 74476 6196 74516 6236
rect 74860 6196 74900 6236
rect 75244 6196 75284 6236
rect 75532 6196 75572 6236
rect 77068 6196 77108 6236
rect 77260 6196 77300 6236
rect 81772 6196 81812 6236
rect 84556 6196 84596 6236
rect 98668 6196 98708 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 65408 6028 65448 6068
rect 65490 6028 65530 6068
rect 65572 6028 65612 6068
rect 65654 6028 65694 6068
rect 65736 6028 65776 6068
rect 80528 6028 80568 6068
rect 80610 6028 80650 6068
rect 80692 6028 80732 6068
rect 80774 6028 80814 6068
rect 80856 6028 80896 6068
rect 95648 6028 95688 6068
rect 95730 6028 95770 6068
rect 95812 6028 95852 6068
rect 95894 6028 95934 6068
rect 95976 6028 96016 6068
rect 16972 5860 17012 5900
rect 23020 5860 23060 5900
rect 45388 5860 45428 5900
rect 53356 5860 53396 5900
rect 56812 5860 56852 5900
rect 61324 5860 61364 5900
rect 65068 5860 65108 5900
rect 72076 5860 72116 5900
rect 79372 5860 79412 5900
rect 41740 5776 41780 5816
rect 15340 5692 15380 5732
rect 15532 5692 15572 5732
rect 15724 5692 15764 5732
rect 15916 5692 15956 5732
rect 16108 5692 16148 5732
rect 16300 5692 16340 5732
rect 16492 5692 16532 5732
rect 16684 5692 16724 5732
rect 16876 5692 16916 5732
rect 17068 5692 17108 5732
rect 17260 5692 17300 5732
rect 17452 5692 17492 5732
rect 18124 5692 18164 5732
rect 18316 5692 18356 5732
rect 18604 5692 18644 5732
rect 18796 5692 18836 5732
rect 18988 5692 19028 5732
rect 19180 5692 19220 5732
rect 19372 5692 19412 5732
rect 19564 5692 19604 5732
rect 19756 5692 19796 5732
rect 19948 5692 19988 5732
rect 20140 5692 20180 5732
rect 20332 5692 20372 5732
rect 20524 5692 20564 5732
rect 20716 5692 20756 5732
rect 22732 5692 22772 5732
rect 23020 5692 23060 5732
rect 23212 5692 23252 5732
rect 23308 5692 23348 5732
rect 23788 5692 23828 5732
rect 23980 5692 24020 5732
rect 24172 5692 24212 5732
rect 24364 5692 24404 5732
rect 24748 5692 24788 5732
rect 24940 5692 24980 5732
rect 26572 5692 26612 5732
rect 26764 5692 26804 5732
rect 26956 5692 26996 5732
rect 27148 5692 27188 5732
rect 28492 5692 28532 5732
rect 28684 5692 28724 5732
rect 28972 5692 29012 5732
rect 29164 5692 29204 5732
rect 30124 5692 30164 5732
rect 30316 5692 30356 5732
rect 30604 5692 30644 5732
rect 30796 5692 30836 5732
rect 31084 5692 31124 5732
rect 31276 5692 31316 5732
rect 31468 5692 31508 5732
rect 31660 5692 31700 5732
rect 31852 5692 31892 5732
rect 32044 5692 32084 5732
rect 32236 5692 32276 5732
rect 32428 5692 32468 5732
rect 32620 5692 32660 5732
rect 32812 5692 32852 5732
rect 34156 5692 34196 5732
rect 34348 5692 34388 5732
rect 34540 5692 34580 5732
rect 34732 5692 34772 5732
rect 34924 5692 34964 5732
rect 35116 5692 35156 5732
rect 35404 5692 35444 5732
rect 35596 5692 35636 5732
rect 36076 5692 36116 5732
rect 36268 5692 36308 5732
rect 36460 5692 36500 5732
rect 36652 5692 36692 5732
rect 36844 5692 36884 5732
rect 37036 5703 37076 5743
rect 37228 5692 37268 5732
rect 37516 5692 37556 5732
rect 37708 5692 37748 5732
rect 37900 5692 37940 5732
rect 38092 5692 38132 5732
rect 38572 5692 38612 5732
rect 38764 5692 38804 5732
rect 39148 5692 39188 5732
rect 39340 5692 39380 5732
rect 42604 5692 42644 5732
rect 44044 5692 44084 5732
rect 44236 5692 44276 5732
rect 44332 5692 44372 5732
rect 44524 5692 44564 5732
rect 44716 5692 44756 5732
rect 44812 5692 44852 5732
rect 45100 5692 45140 5732
rect 45196 5692 45236 5732
rect 45388 5692 45428 5732
rect 45676 5692 45716 5732
rect 46636 5692 46676 5732
rect 48652 5692 48692 5732
rect 49612 5692 49652 5732
rect 52204 5692 52244 5732
rect 52396 5692 52436 5732
rect 52492 5692 52532 5732
rect 53740 5692 53780 5732
rect 53932 5692 53972 5732
rect 54316 5692 54356 5732
rect 54508 5692 54548 5732
rect 55660 5692 55700 5732
rect 55756 5692 55796 5732
rect 55852 5692 55892 5732
rect 56332 5692 56372 5732
rect 56524 5692 56564 5732
rect 56716 5692 56756 5732
rect 56908 5692 56948 5732
rect 57292 5692 57332 5732
rect 57676 5700 57716 5740
rect 58252 5692 58292 5732
rect 61228 5692 61268 5732
rect 61324 5692 61364 5732
rect 61996 5692 62036 5732
rect 64588 5692 64628 5732
rect 67276 5692 67316 5732
rect 67468 5692 67508 5732
rect 68332 5692 68372 5732
rect 68524 5692 68564 5732
rect 68716 5692 68756 5732
rect 68908 5692 68948 5732
rect 69580 5692 69620 5732
rect 69772 5692 69812 5732
rect 71308 5692 71348 5732
rect 71500 5692 71540 5732
rect 71980 5692 72020 5732
rect 72172 5692 72212 5732
rect 72364 5692 72404 5732
rect 72556 5692 72596 5732
rect 72748 5692 72788 5732
rect 72940 5692 72980 5732
rect 73420 5692 73460 5732
rect 73612 5692 73652 5732
rect 73804 5692 73844 5732
rect 73996 5692 74036 5732
rect 74284 5692 74324 5732
rect 74476 5692 74516 5732
rect 74956 5692 74996 5732
rect 75052 5692 75092 5732
rect 75724 5692 75764 5732
rect 75916 5692 75956 5732
rect 77260 5692 77300 5732
rect 77452 5692 77492 5732
rect 78028 5692 78068 5732
rect 78508 5692 78548 5732
rect 78700 5692 78740 5732
rect 78892 5692 78932 5732
rect 79084 5692 79124 5732
rect 79276 5692 79316 5732
rect 79468 5692 79508 5732
rect 79660 5692 79700 5732
rect 79852 5692 79892 5732
rect 80044 5692 80084 5732
rect 80236 5692 80276 5732
rect 80428 5692 80468 5732
rect 80620 5692 80660 5732
rect 80908 5692 80948 5732
rect 81100 5692 81140 5732
rect 81292 5692 81332 5732
rect 81484 5692 81524 5732
rect 81676 5692 81716 5732
rect 81868 5692 81908 5732
rect 82156 5692 82196 5732
rect 82348 5692 82388 5732
rect 82540 5692 82580 5732
rect 82732 5692 82772 5732
rect 82924 5692 82964 5732
rect 83116 5692 83156 5732
rect 83308 5692 83348 5732
rect 83500 5692 83540 5732
rect 83692 5692 83732 5732
rect 83884 5692 83924 5732
rect 84556 5692 84596 5732
rect 1708 5608 1748 5648
rect 2092 5608 2132 5648
rect 17740 5608 17780 5648
rect 19084 5608 19124 5648
rect 20236 5608 20276 5648
rect 21004 5608 21044 5648
rect 21388 5608 21428 5648
rect 28108 5608 28148 5648
rect 29548 5608 29588 5648
rect 29932 5608 29972 5648
rect 33772 5608 33812 5648
rect 39244 5608 39284 5648
rect 39724 5608 39764 5648
rect 40108 5608 40148 5648
rect 41260 5608 41300 5648
rect 42892 5608 42932 5648
rect 43276 5608 43316 5648
rect 43660 5608 43700 5648
rect 47116 5608 47156 5648
rect 47500 5608 47540 5648
rect 47884 5608 47924 5648
rect 48268 5608 48308 5648
rect 50092 5608 50132 5648
rect 53164 5608 53204 5648
rect 54892 5608 54932 5648
rect 55276 5608 55316 5648
rect 58732 5608 58772 5648
rect 59116 5608 59156 5648
rect 59500 5608 59540 5648
rect 59884 5608 59924 5648
rect 60268 5608 60308 5648
rect 60652 5608 60692 5648
rect 61804 5608 61844 5648
rect 62476 5608 62516 5648
rect 62860 5608 62900 5648
rect 63244 5608 63284 5648
rect 63628 5608 63668 5648
rect 64012 5608 64052 5648
rect 66988 5608 67028 5648
rect 67852 5608 67892 5648
rect 68812 5608 68852 5648
rect 69292 5608 69332 5648
rect 70156 5621 70196 5661
rect 70540 5608 70580 5648
rect 70924 5608 70964 5648
rect 73516 5608 73556 5648
rect 74860 5608 74900 5648
rect 75532 5608 75572 5648
rect 76300 5608 76340 5648
rect 76684 5608 76724 5648
rect 77068 5608 77108 5648
rect 77836 5608 77876 5648
rect 82636 5608 82676 5648
rect 84364 5608 84404 5648
rect 85036 5608 85076 5648
rect 85420 5608 85460 5648
rect 85804 5608 85844 5648
rect 86188 5608 86228 5648
rect 86590 5621 86630 5661
rect 97516 5608 97556 5648
rect 97900 5608 97940 5648
rect 98476 5608 98516 5648
rect 17260 5524 17300 5564
rect 19756 5524 19796 5564
rect 56524 5524 56564 5564
rect 57292 5550 57332 5590
rect 57676 5524 57716 5564
rect 57868 5524 57908 5564
rect 58252 5524 58292 5564
rect 61900 5524 61940 5564
rect 63820 5524 63860 5564
rect 74476 5524 74516 5564
rect 75916 5524 75956 5564
rect 79084 5524 79124 5564
rect 83884 5524 83924 5564
rect 1516 5440 1556 5480
rect 1900 5440 1940 5480
rect 15340 5440 15380 5480
rect 15724 5440 15764 5480
rect 16108 5440 16148 5480
rect 16492 5440 16532 5480
rect 17932 5440 17972 5480
rect 18124 5440 18164 5480
rect 18604 5440 18644 5480
rect 19372 5440 19412 5480
rect 20524 5440 20564 5480
rect 21196 5440 21236 5480
rect 21580 5440 21620 5480
rect 22444 5440 22484 5480
rect 23788 5440 23828 5480
rect 24172 5440 24212 5480
rect 26764 5440 26804 5480
rect 27148 5440 27188 5480
rect 28300 5440 28340 5480
rect 28492 5440 28532 5480
rect 29356 5440 29396 5480
rect 29740 5440 29780 5480
rect 31084 5440 31124 5480
rect 31660 5440 31700 5480
rect 32044 5440 32084 5480
rect 32428 5440 32468 5480
rect 32812 5440 32852 5480
rect 33964 5440 34004 5480
rect 34348 5440 34388 5480
rect 34732 5440 34772 5480
rect 35116 5440 35156 5480
rect 36268 5440 36308 5480
rect 36652 5440 36692 5480
rect 37036 5440 37076 5480
rect 37324 5440 37364 5480
rect 37708 5440 37748 5480
rect 38092 5440 38132 5480
rect 39532 5440 39572 5480
rect 39916 5440 39956 5480
rect 41068 5440 41108 5480
rect 43084 5440 43124 5480
rect 43468 5440 43508 5480
rect 43852 5440 43892 5480
rect 44236 5440 44276 5480
rect 44524 5440 44564 5480
rect 47308 5440 47348 5480
rect 47692 5440 47732 5480
rect 48076 5440 48116 5480
rect 48460 5440 48500 5480
rect 49900 5440 49940 5480
rect 52204 5440 52244 5480
rect 53932 5440 53972 5480
rect 54316 5440 54356 5480
rect 54700 5440 54740 5480
rect 55084 5440 55124 5480
rect 57100 5440 57140 5480
rect 58060 5440 58100 5480
rect 58540 5440 58580 5480
rect 58924 5440 58964 5480
rect 59308 5440 59348 5480
rect 59692 5440 59732 5480
rect 60076 5440 60116 5480
rect 60460 5440 60500 5480
rect 61036 5440 61076 5480
rect 62284 5440 62324 5480
rect 62668 5440 62708 5480
rect 63052 5440 63092 5480
rect 63436 5440 63476 5480
rect 66796 5440 66836 5480
rect 67660 5440 67700 5480
rect 68332 5440 68372 5480
rect 69100 5440 69140 5480
rect 69772 5440 69812 5480
rect 69964 5440 70004 5480
rect 70348 5440 70388 5480
rect 70732 5440 70772 5480
rect 72556 5440 72596 5480
rect 72940 5440 72980 5480
rect 73996 5440 74036 5480
rect 75340 5440 75380 5480
rect 76108 5440 76148 5480
rect 76492 5440 76532 5480
rect 76876 5440 76916 5480
rect 77452 5440 77492 5480
rect 78028 5440 78068 5480
rect 78700 5440 78740 5480
rect 79852 5440 79892 5480
rect 80044 5440 80084 5480
rect 80620 5440 80660 5480
rect 81100 5440 81140 5480
rect 81484 5440 81524 5480
rect 81868 5440 81908 5480
rect 82348 5440 82388 5480
rect 83116 5440 83156 5480
rect 83500 5440 83540 5480
rect 84556 5440 84596 5480
rect 84844 5440 84884 5480
rect 85228 5440 85268 5480
rect 85612 5440 85652 5480
rect 85996 5440 86036 5480
rect 86380 5440 86420 5480
rect 97708 5440 97748 5480
rect 98092 5440 98132 5480
rect 98284 5440 98324 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 64168 5272 64208 5312
rect 64250 5272 64290 5312
rect 64332 5272 64372 5312
rect 64414 5272 64454 5312
rect 64496 5272 64536 5312
rect 79288 5272 79328 5312
rect 79370 5272 79410 5312
rect 79452 5272 79492 5312
rect 79534 5272 79574 5312
rect 79616 5272 79656 5312
rect 94408 5272 94448 5312
rect 94490 5272 94530 5312
rect 94572 5272 94612 5312
rect 94654 5272 94694 5312
rect 94736 5272 94776 5312
rect 22828 5104 22868 5144
rect 27820 5104 27860 5144
rect 30508 5104 30548 5144
rect 57868 5104 57908 5144
rect 61804 5104 61844 5144
rect 67564 5104 67604 5144
rect 67948 5104 67988 5144
rect 70540 5104 70580 5144
rect 73324 5104 73364 5144
rect 19948 5020 19988 5060
rect 28396 5020 28436 5060
rect 31180 5020 31220 5060
rect 31660 5020 31700 5060
rect 41548 5020 41588 5060
rect 56716 5020 56756 5060
rect 65452 5020 65492 5060
rect 71692 5020 71732 5060
rect 79468 5020 79508 5060
rect 1708 4936 1748 4976
rect 2092 4936 2132 4976
rect 2476 4936 2516 4976
rect 2860 4936 2900 4976
rect 13708 4936 13748 4976
rect 13900 4936 13940 4976
rect 14284 4936 14324 4976
rect 14668 4936 14708 4976
rect 15052 4936 15092 4976
rect 15436 4936 15476 4976
rect 16396 4936 16436 4976
rect 16780 4936 16820 4976
rect 20332 4936 20372 4976
rect 21484 4936 21524 4976
rect 23788 4923 23828 4963
rect 24652 4936 24692 4976
rect 25900 4936 25940 4976
rect 26092 4936 26132 4976
rect 26476 4936 26516 4976
rect 26860 4936 26900 4976
rect 27244 4936 27284 4976
rect 29164 4936 29204 4976
rect 29548 4936 29588 4976
rect 29932 4936 29972 4976
rect 32236 4936 32276 4976
rect 32620 4936 32660 4976
rect 33004 4936 33044 4976
rect 33388 4936 33428 4976
rect 33772 4936 33812 4976
rect 34156 4936 34196 4976
rect 36652 4936 36692 4976
rect 37132 4936 37172 4976
rect 37516 4936 37556 4976
rect 37900 4936 37940 4976
rect 40204 4936 40244 4976
rect 40588 4936 40628 4976
rect 40972 4936 41012 4976
rect 41356 4936 41396 4976
rect 41740 4936 41780 4976
rect 47980 4936 48020 4976
rect 48364 4936 48404 4976
rect 48748 4936 48788 4976
rect 49132 4936 49172 4976
rect 52396 4936 52436 4976
rect 55756 4936 55796 4976
rect 56428 4936 56468 4976
rect 15820 4852 15860 4892
rect 16012 4852 16052 4892
rect 17164 4865 17204 4905
rect 17356 4852 17396 4892
rect 17548 4852 17588 4892
rect 17740 4841 17780 4881
rect 18028 4852 18068 4892
rect 18220 4852 18260 4892
rect 18604 4852 18644 4892
rect 18796 4852 18836 4892
rect 18988 4852 19028 4892
rect 19180 4852 19220 4892
rect 19372 4852 19412 4892
rect 19564 4852 19604 4892
rect 19948 4852 19988 4892
rect 20121 4852 20161 4892
rect 20716 4865 20756 4905
rect 20908 4852 20948 4892
rect 21100 4852 21140 4892
rect 21292 4852 21332 4892
rect 21868 4852 21908 4892
rect 22060 4852 22100 4892
rect 22252 4852 22292 4892
rect 22444 4852 22484 4892
rect 22636 4852 22676 4892
rect 22828 4852 22868 4892
rect 22924 4852 22964 4892
rect 23404 4852 23444 4892
rect 23596 4852 23636 4892
rect 24172 4852 24212 4892
rect 24364 4852 24404 4892
rect 24556 4852 24596 4892
rect 24748 4852 24788 4892
rect 24940 4852 24980 4892
rect 25132 4852 25172 4892
rect 25324 4852 25364 4892
rect 25516 4852 25556 4892
rect 27628 4852 27668 4892
rect 27820 4852 27860 4892
rect 28012 4852 28052 4892
rect 28204 4852 28244 4892
rect 28396 4852 28436 4892
rect 28588 4852 28628 4892
rect 28780 4852 28820 4892
rect 28972 4852 29012 4892
rect 30316 4852 30356 4892
rect 30508 4852 30548 4892
rect 30700 4852 30740 4892
rect 30892 4852 30932 4892
rect 31180 4852 31220 4892
rect 31372 4852 31412 4892
rect 31660 4841 31700 4881
rect 31852 4852 31892 4892
rect 34540 4852 34580 4892
rect 34732 4852 34772 4892
rect 34924 4852 34964 4892
rect 35116 4852 35156 4892
rect 35308 4841 35348 4881
rect 35500 4841 35540 4881
rect 35692 4852 35732 4892
rect 35884 4852 35924 4892
rect 36076 4852 36116 4892
rect 36268 4852 36308 4892
rect 36556 4852 36596 4892
rect 36748 4852 36788 4892
rect 38284 4852 38324 4892
rect 38476 4852 38516 4892
rect 38668 4852 38708 4892
rect 38860 4852 38900 4892
rect 39052 4852 39092 4892
rect 39244 4852 39284 4892
rect 39628 4852 39668 4892
rect 39820 4852 39860 4892
rect 42988 4852 43028 4892
rect 44332 4852 44372 4892
rect 45580 4852 45620 4892
rect 45868 4852 45908 4892
rect 46060 4852 46100 4892
rect 46156 4852 46196 4892
rect 46540 4852 46580 4892
rect 46828 4894 46868 4934
rect 56908 4936 56948 4976
rect 58828 4936 58868 4976
rect 59212 4936 59252 4976
rect 60364 4936 60404 4976
rect 60748 4936 60788 4976
rect 62764 4936 62804 4976
rect 63916 4936 63956 4976
rect 64300 4936 64340 4976
rect 66124 4936 66164 4976
rect 66508 4936 66548 4976
rect 66892 4936 66932 4976
rect 68908 4936 68948 4976
rect 69292 4936 69332 4976
rect 69676 4936 69716 4976
rect 70924 4936 70964 4976
rect 73708 4936 73748 4976
rect 75916 4936 75956 4976
rect 77548 4936 77588 4976
rect 78508 4936 78548 4976
rect 78892 4936 78932 4976
rect 79852 4936 79892 4976
rect 80236 4936 80276 4976
rect 80620 4936 80660 4976
rect 80908 4936 80948 4976
rect 82156 4936 82196 4976
rect 82540 4936 82580 4976
rect 85804 4936 85844 4976
rect 86188 4936 86228 4976
rect 86572 4936 86612 4976
rect 86956 4936 86996 4976
rect 87340 4936 87380 4976
rect 87724 4936 87764 4976
rect 88108 4936 88148 4976
rect 88492 4936 88532 4976
rect 97132 4936 97172 4976
rect 97708 4936 97748 4976
rect 98092 4936 98132 4976
rect 98476 4936 98516 4976
rect 46636 4852 46676 4892
rect 47020 4852 47060 4892
rect 47116 4852 47156 4892
rect 47308 4852 47348 4892
rect 47500 4852 47540 4892
rect 47596 4852 47636 4892
rect 47788 4852 47828 4892
rect 49516 4852 49556 4892
rect 49708 4852 49748 4892
rect 49900 4852 49940 4892
rect 50092 4852 50132 4892
rect 50284 4852 50324 4892
rect 50476 4852 50516 4892
rect 50668 4852 50708 4892
rect 50865 4865 50905 4905
rect 52780 4852 52820 4892
rect 54028 4852 54068 4892
rect 54988 4852 55028 4892
rect 55180 4852 55220 4892
rect 55372 4852 55412 4892
rect 55948 4852 55988 4892
rect 56140 4852 56180 4892
rect 56332 4852 56372 4892
rect 56524 4831 56564 4871
rect 57100 4852 57140 4892
rect 57292 4852 57332 4892
rect 57484 4852 57524 4892
rect 57676 4852 57716 4892
rect 57868 4852 57908 4892
rect 58060 4852 58100 4892
rect 58252 4852 58292 4892
rect 58444 4852 58484 4892
rect 59692 4852 59732 4892
rect 59884 4852 59924 4892
rect 61324 4852 61364 4892
rect 61708 4852 61748 4892
rect 61900 4831 61940 4871
rect 62092 4852 62132 4892
rect 62284 4852 62324 4892
rect 63244 4852 63284 4892
rect 63436 4852 63476 4892
rect 64780 4852 64820 4892
rect 67180 4852 67220 4892
rect 67372 4852 67412 4892
rect 67564 4852 67604 4892
rect 67756 4852 67796 4892
rect 67948 4852 67988 4892
rect 68140 4865 68180 4905
rect 68332 4852 68372 4892
rect 68524 4852 68564 4892
rect 69580 4852 69620 4892
rect 69772 4852 69812 4892
rect 69964 4852 70004 4892
rect 70156 4852 70196 4892
rect 70348 4852 70388 4892
rect 70540 4852 70580 4892
rect 71116 4852 71156 4892
rect 71308 4852 71348 4892
rect 71500 4852 71540 4892
rect 71692 4852 71732 4892
rect 71980 4852 72020 4892
rect 72172 4852 72212 4892
rect 72364 4852 72404 4892
rect 72556 4852 72596 4892
rect 72751 4841 72791 4881
rect 72940 4852 72980 4892
rect 73127 4865 73167 4905
rect 73324 4852 73364 4892
rect 74188 4852 74228 4892
rect 74380 4852 74420 4892
rect 74668 4852 74708 4892
rect 75820 4852 75860 4892
rect 76012 4852 76052 4892
rect 76207 4841 76247 4881
rect 76396 4852 76436 4892
rect 76588 4852 76628 4892
rect 76780 4852 76820 4892
rect 76972 4852 77012 4892
rect 77164 4852 77204 4892
rect 77836 4852 77876 4892
rect 78028 4852 78068 4892
rect 79276 4852 79316 4892
rect 79468 4852 79508 4892
rect 80812 4852 80852 4892
rect 81004 4852 81044 4892
rect 81196 4852 81236 4892
rect 81388 4865 81428 4905
rect 81580 4852 81620 4892
rect 81772 4852 81812 4892
rect 82732 4852 82772 4892
rect 82924 4852 82964 4892
rect 83308 4852 83348 4892
rect 83500 4852 83540 4892
rect 83692 4852 83732 4892
rect 83884 4852 83924 4892
rect 84556 4852 84596 4892
rect 19084 4768 19124 4808
rect 20812 4768 20852 4808
rect 35404 4768 35444 4808
rect 42220 4768 42260 4808
rect 43468 4768 43508 4808
rect 44716 4768 44756 4808
rect 49612 4768 49652 4808
rect 49996 4768 50036 4808
rect 53644 4768 53684 4808
rect 56044 4768 56084 4808
rect 72076 4768 72116 4808
rect 1516 4684 1556 4724
rect 1900 4684 1940 4724
rect 2284 4684 2324 4724
rect 2668 4684 2708 4724
rect 13516 4684 13556 4724
rect 14092 4684 14132 4724
rect 14476 4684 14516 4724
rect 14860 4684 14900 4724
rect 15244 4684 15284 4724
rect 15628 4684 15668 4724
rect 15916 4684 15956 4724
rect 16588 4684 16628 4724
rect 16972 4684 17012 4724
rect 17260 4684 17300 4724
rect 17644 4684 17684 4724
rect 18700 4684 18740 4724
rect 19468 4684 19508 4724
rect 20524 4684 20564 4724
rect 21196 4684 21236 4724
rect 21676 4684 21716 4724
rect 21964 4684 22004 4724
rect 22348 4684 22388 4724
rect 23500 4684 23540 4724
rect 23980 4684 24020 4724
rect 24268 4684 24308 4724
rect 25036 4684 25076 4724
rect 25420 4684 25460 4724
rect 25708 4684 25748 4724
rect 26284 4684 26324 4724
rect 26668 4684 26708 4724
rect 27052 4684 27092 4724
rect 27436 4684 27476 4724
rect 28108 4684 28148 4724
rect 28876 4684 28916 4724
rect 29356 4684 29396 4724
rect 29740 4684 29780 4724
rect 30124 4684 30164 4724
rect 30796 4684 30836 4724
rect 32428 4684 32468 4724
rect 32812 4684 32852 4724
rect 33196 4684 33236 4724
rect 33580 4684 33620 4724
rect 33964 4684 34004 4724
rect 34348 4684 34388 4724
rect 34636 4684 34676 4724
rect 35020 4684 35060 4724
rect 35788 4684 35828 4724
rect 37324 4684 37364 4724
rect 37708 4684 37748 4724
rect 38092 4684 38132 4724
rect 38380 4684 38420 4724
rect 38764 4684 38804 4724
rect 39724 4684 39764 4724
rect 40396 4684 40436 4724
rect 40780 4684 40820 4724
rect 41164 4684 41204 4724
rect 41932 4684 41972 4724
rect 45868 4684 45908 4724
rect 46828 4684 46868 4724
rect 47308 4684 47348 4724
rect 47788 4684 47828 4724
rect 48172 4684 48212 4724
rect 48556 4684 48596 4724
rect 48940 4684 48980 4724
rect 49324 4684 49364 4724
rect 50380 4684 50420 4724
rect 50764 4684 50804 4724
rect 52204 4684 52244 4724
rect 55276 4684 55316 4724
rect 55564 4684 55604 4724
rect 57196 4684 57236 4724
rect 57580 4684 57620 4724
rect 58348 4684 58388 4724
rect 58636 4684 58676 4724
rect 59020 4684 59060 4724
rect 59692 4684 59732 4724
rect 60172 4684 60212 4724
rect 60556 4684 60596 4724
rect 61228 4684 61268 4724
rect 61516 4684 61556 4724
rect 62572 4684 62612 4724
rect 63724 4684 63764 4724
rect 64108 4684 64148 4724
rect 65932 4684 65972 4724
rect 66316 4684 66356 4724
rect 66700 4684 66740 4724
rect 67276 4684 67316 4724
rect 68428 4684 68468 4724
rect 68716 4684 68756 4724
rect 69100 4684 69140 4724
rect 70060 4684 70100 4724
rect 70732 4684 70772 4724
rect 71212 4684 71252 4724
rect 72460 4684 72500 4724
rect 72844 4684 72884 4724
rect 73516 4684 73556 4724
rect 74284 4684 74324 4724
rect 75148 4684 75188 4724
rect 76300 4684 76340 4724
rect 76684 4684 76724 4724
rect 77068 4684 77108 4724
rect 77356 4684 77396 4724
rect 78316 4684 78356 4724
rect 78700 4684 78740 4724
rect 79660 4684 79700 4724
rect 80044 4684 80084 4724
rect 80428 4684 80468 4724
rect 81292 4684 81332 4724
rect 81676 4684 81716 4724
rect 81964 4684 82004 4724
rect 82348 4684 82388 4724
rect 82828 4684 82868 4724
rect 83404 4684 83444 4724
rect 83788 4684 83828 4724
rect 84940 4684 84980 4724
rect 85612 4684 85652 4724
rect 85996 4684 86036 4724
rect 86380 4684 86420 4724
rect 86764 4684 86804 4724
rect 87148 4684 87188 4724
rect 87532 4684 87572 4724
rect 87916 4684 87956 4724
rect 88300 4684 88340 4724
rect 97324 4684 97364 4724
rect 97516 4684 97556 4724
rect 97900 4684 97940 4724
rect 98284 4684 98324 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 65408 4516 65448 4556
rect 65490 4516 65530 4556
rect 65572 4516 65612 4556
rect 65654 4516 65694 4556
rect 65736 4516 65776 4556
rect 80528 4516 80568 4556
rect 80610 4516 80650 4556
rect 80692 4516 80732 4556
rect 80774 4516 80814 4556
rect 80856 4516 80896 4556
rect 95648 4516 95688 4556
rect 95730 4516 95770 4556
rect 95812 4516 95852 4556
rect 95894 4516 95934 4556
rect 95976 4516 96016 4556
rect 35020 4390 35060 4430
rect 34060 4348 34100 4388
rect 35788 4348 35828 4388
rect 45484 4348 45524 4388
rect 53164 4348 53204 4388
rect 55180 4348 55220 4388
rect 56716 4348 56756 4388
rect 61228 4348 61268 4388
rect 69004 4348 69044 4388
rect 70924 4348 70964 4388
rect 72844 4348 72884 4388
rect 85420 4348 85460 4388
rect 22732 4264 22772 4304
rect 47596 4264 47636 4304
rect 64204 4264 64244 4304
rect 77644 4264 77684 4304
rect 16972 4180 17012 4220
rect 17164 4180 17204 4220
rect 17356 4180 17396 4220
rect 17548 4191 17588 4231
rect 18892 4180 18932 4220
rect 19084 4180 19124 4220
rect 19564 4180 19604 4220
rect 19756 4180 19796 4220
rect 19948 4180 19988 4220
rect 20145 4180 20185 4220
rect 21100 4180 21140 4220
rect 21292 4180 21332 4220
rect 21484 4180 21524 4220
rect 21676 4180 21716 4220
rect 21868 4180 21908 4220
rect 22060 4180 22100 4220
rect 22252 4180 22292 4220
rect 22444 4180 22484 4220
rect 22636 4180 22676 4220
rect 22828 4180 22868 4220
rect 23788 4180 23828 4220
rect 23980 4180 24020 4220
rect 24172 4180 24212 4220
rect 24364 4180 24404 4220
rect 24556 4180 24596 4220
rect 24748 4180 24788 4220
rect 24940 4180 24980 4220
rect 25132 4180 25172 4220
rect 27244 4180 27284 4220
rect 27436 4180 27476 4220
rect 27628 4180 27668 4220
rect 27820 4180 27860 4220
rect 28012 4180 28052 4220
rect 28204 4180 28244 4220
rect 29260 4179 29300 4219
rect 29452 4180 29492 4220
rect 29932 4180 29972 4220
rect 30124 4180 30164 4220
rect 30316 4180 30356 4220
rect 30508 4180 30548 4220
rect 30700 4180 30740 4220
rect 30892 4180 30932 4220
rect 31084 4180 31124 4220
rect 31276 4180 31316 4220
rect 33868 4180 33908 4220
rect 34060 4180 34100 4220
rect 34444 4180 34484 4220
rect 34636 4180 34676 4220
rect 35020 4180 35060 4220
rect 35212 4180 35252 4220
rect 35588 4179 35628 4219
rect 35788 4180 35828 4220
rect 37612 4180 37652 4220
rect 37804 4180 37844 4220
rect 37996 4180 38036 4220
rect 38188 4180 38228 4220
rect 38380 4180 38420 4220
rect 38572 4180 38612 4220
rect 38764 4180 38804 4220
rect 38956 4180 38996 4220
rect 39148 4180 39188 4220
rect 39340 4180 39380 4220
rect 44620 4180 44660 4220
rect 45964 4180 46004 4220
rect 47116 4180 47156 4220
rect 48460 4180 48500 4220
rect 49036 4180 49076 4220
rect 49228 4180 49268 4220
rect 49516 4177 49556 4217
rect 49996 4180 50036 4220
rect 51532 4180 51572 4220
rect 52012 4180 52052 4220
rect 52108 4180 52148 4220
rect 52204 4180 52244 4220
rect 52396 4180 52436 4220
rect 52588 4180 52628 4220
rect 52972 4180 53012 4220
rect 53356 4180 53396 4220
rect 53548 4180 53588 4220
rect 54604 4180 54644 4220
rect 54796 4180 54836 4220
rect 55084 4180 55124 4220
rect 55276 4180 55316 4220
rect 56524 4180 56564 4220
rect 57004 4180 57044 4220
rect 57580 4180 57620 4220
rect 57964 4180 58004 4220
rect 58828 4180 58868 4220
rect 59212 4180 59252 4220
rect 60172 4180 60212 4220
rect 60460 4169 60500 4209
rect 60652 4180 60692 4220
rect 60940 4180 60980 4220
rect 61036 4180 61076 4220
rect 63436 4180 63476 4220
rect 64588 4180 64628 4220
rect 64780 4180 64820 4220
rect 66892 4180 66932 4220
rect 67084 4180 67124 4220
rect 67756 4180 67796 4220
rect 67948 4180 67988 4220
rect 68140 4180 68180 4220
rect 68332 4180 68372 4220
rect 68524 4180 68564 4220
rect 68716 4180 68756 4220
rect 68908 4180 68948 4220
rect 69100 4180 69140 4220
rect 70060 4180 70100 4220
rect 70252 4180 70292 4220
rect 70444 4180 70484 4220
rect 70636 4180 70676 4220
rect 70828 4180 70868 4220
rect 71020 4180 71060 4220
rect 71212 4180 71252 4220
rect 71404 4180 71444 4220
rect 71596 4180 71636 4220
rect 71788 4180 71828 4220
rect 71980 4180 72020 4220
rect 72172 4180 72212 4220
rect 72748 4180 72788 4220
rect 72940 4180 72980 4220
rect 73132 4180 73172 4220
rect 73324 4180 73364 4220
rect 73516 4180 73556 4220
rect 73708 4180 73748 4220
rect 74668 4180 74708 4220
rect 74860 4180 74900 4220
rect 75820 4180 75860 4220
rect 76012 4180 76052 4220
rect 76588 4180 76628 4220
rect 76780 4180 76820 4220
rect 77164 4180 77204 4220
rect 77356 4180 77396 4220
rect 78412 4180 78452 4220
rect 78796 4180 78836 4220
rect 78988 4180 79028 4220
rect 80716 4180 80756 4220
rect 80908 4180 80948 4220
rect 81292 4180 81332 4220
rect 83212 4180 83252 4220
rect 83404 4180 83444 4220
rect 84268 4180 84308 4220
rect 85324 4180 85364 4220
rect 85516 4180 85556 4220
rect 1516 4096 1556 4136
rect 1900 4096 1940 4136
rect 2284 4096 2324 4136
rect 2668 4096 2708 4136
rect 3052 4096 3092 4136
rect 3436 4096 3476 4136
rect 3820 4096 3860 4136
rect 4204 4096 4244 4136
rect 4588 4096 4628 4136
rect 4972 4096 5012 4136
rect 5356 4096 5396 4136
rect 5740 4096 5780 4136
rect 6124 4096 6164 4136
rect 6508 4096 6548 4136
rect 6892 4096 6932 4136
rect 7276 4096 7316 4136
rect 7660 4096 7700 4136
rect 8044 4096 8084 4136
rect 8428 4096 8468 4136
rect 8812 4096 8852 4136
rect 9196 4096 9236 4136
rect 9580 4096 9620 4136
rect 9964 4096 10004 4136
rect 10348 4096 10388 4136
rect 10732 4096 10772 4136
rect 11116 4096 11156 4136
rect 11500 4096 11540 4136
rect 11884 4096 11924 4136
rect 12268 4096 12308 4136
rect 12652 4096 12692 4136
rect 13036 4096 13076 4136
rect 13420 4096 13460 4136
rect 13804 4096 13844 4136
rect 14188 4096 14228 4136
rect 14572 4096 14612 4136
rect 14956 4096 14996 4136
rect 15340 4096 15380 4136
rect 15724 4096 15764 4136
rect 16108 4096 16148 4136
rect 16492 4096 16532 4136
rect 17740 4096 17780 4136
rect 18124 4096 18164 4136
rect 18508 4096 18548 4136
rect 20332 4096 20372 4136
rect 20716 4096 20756 4136
rect 22348 4096 22388 4136
rect 23020 4096 23060 4136
rect 23404 4096 23444 4136
rect 24268 4096 24308 4136
rect 25036 4096 25076 4136
rect 25324 4096 25364 4136
rect 25708 4096 25748 4136
rect 26092 4096 26132 4136
rect 26476 4096 26516 4136
rect 26860 4096 26900 4136
rect 28396 4096 28436 4136
rect 28780 4096 28820 4136
rect 31180 4096 31220 4136
rect 31468 4096 31508 4136
rect 31852 4096 31892 4136
rect 32236 4096 32276 4136
rect 32620 4096 32660 4136
rect 33004 4096 33044 4136
rect 33388 4096 33428 4136
rect 36076 4096 36116 4136
rect 36460 4109 36500 4149
rect 36844 4096 36884 4136
rect 37228 4109 37268 4149
rect 39532 4109 39572 4149
rect 39916 4096 39956 4136
rect 40300 4096 40340 4136
rect 40684 4096 40724 4136
rect 41068 4096 41108 4136
rect 41452 4096 41492 4136
rect 41836 4096 41876 4136
rect 42220 4096 42260 4136
rect 42604 4096 42644 4136
rect 42988 4096 43028 4136
rect 43372 4096 43412 4136
rect 50860 4096 50900 4136
rect 51244 4096 51284 4136
rect 51724 4096 51764 4136
rect 53932 4096 53972 4136
rect 54316 4096 54356 4136
rect 55660 4096 55700 4136
rect 56044 4096 56084 4136
rect 61612 4096 61652 4136
rect 61996 4096 62036 4136
rect 62380 4096 62420 4136
rect 62764 4096 62804 4136
rect 65260 4096 65300 4136
rect 65644 4096 65684 4136
rect 66028 4096 66068 4136
rect 66412 4096 66452 4136
rect 67564 4096 67604 4136
rect 69484 4096 69524 4136
rect 69868 4096 69908 4136
rect 71308 4096 71348 4136
rect 72556 4096 72596 4136
rect 74092 4096 74132 4136
rect 74476 4096 74516 4136
rect 75244 4096 75284 4136
rect 75628 4096 75668 4136
rect 76396 4096 76436 4136
rect 79372 4096 79412 4136
rect 79756 4096 79796 4136
rect 80140 4096 80180 4136
rect 80524 4096 80564 4136
rect 82636 4096 82676 4136
rect 83020 4096 83060 4136
rect 83788 4096 83828 4136
rect 85900 4096 85940 4136
rect 86284 4096 86324 4136
rect 86668 4096 86708 4136
rect 87052 4096 87092 4136
rect 87436 4096 87476 4136
rect 87820 4096 87860 4136
rect 88204 4096 88244 4136
rect 88588 4096 88628 4136
rect 88972 4109 89012 4149
rect 89356 4096 89396 4136
rect 89740 4096 89780 4136
rect 90124 4096 90164 4136
rect 90508 4096 90548 4136
rect 90892 4096 90932 4136
rect 91276 4096 91316 4136
rect 91660 4096 91700 4136
rect 92044 4096 92084 4136
rect 92428 4096 92468 4136
rect 92812 4096 92852 4136
rect 93196 4096 93236 4136
rect 93580 4096 93620 4136
rect 93964 4096 94004 4136
rect 94348 4096 94388 4136
rect 94732 4096 94772 4136
rect 95116 4096 95156 4136
rect 95500 4096 95540 4136
rect 95884 4096 95924 4136
rect 96268 4096 96308 4136
rect 96652 4096 96692 4136
rect 97036 4096 97076 4136
rect 97420 4109 97460 4149
rect 97804 4096 97844 4136
rect 98188 4096 98228 4136
rect 98572 4096 98612 4136
rect 21100 4012 21140 4052
rect 23980 4012 24020 4052
rect 28012 4012 28052 4052
rect 29260 4012 29300 4052
rect 30892 4012 30932 4052
rect 34444 4012 34484 4052
rect 38572 4012 38612 4052
rect 42796 4012 42836 4052
rect 49516 4012 49556 4052
rect 49996 4012 50036 4052
rect 50188 4012 50228 4052
rect 51628 4012 51668 4052
rect 52972 4012 53012 4052
rect 56524 4012 56564 4052
rect 57004 4012 57044 4052
rect 57580 4012 57620 4052
rect 60460 4012 60500 4052
rect 63628 4012 63668 4052
rect 64780 4012 64820 4052
rect 67084 4012 67124 4052
rect 68524 4012 68564 4052
rect 70444 4012 70484 4052
rect 74860 4012 74900 4052
rect 81580 4012 81620 4052
rect 84460 4012 84500 4052
rect 86092 4012 86132 4052
rect 94924 4012 94964 4052
rect 1708 3928 1748 3968
rect 2092 3928 2132 3968
rect 2476 3928 2516 3968
rect 2860 3928 2900 3968
rect 3244 3928 3284 3968
rect 3628 3928 3668 3968
rect 4012 3928 4052 3968
rect 4396 3928 4436 3968
rect 4780 3928 4820 3968
rect 5164 3928 5204 3968
rect 5548 3928 5588 3968
rect 5932 3928 5972 3968
rect 6316 3928 6356 3968
rect 6700 3928 6740 3968
rect 7084 3928 7124 3968
rect 7468 3928 7508 3968
rect 7852 3928 7892 3968
rect 8236 3928 8276 3968
rect 8620 3928 8660 3968
rect 9004 3928 9044 3968
rect 9388 3928 9428 3968
rect 9772 3928 9812 3968
rect 10156 3928 10196 3968
rect 10540 3928 10580 3968
rect 10924 3928 10964 3968
rect 11308 3928 11348 3968
rect 11692 3928 11732 3968
rect 12076 3928 12116 3968
rect 12460 3928 12500 3968
rect 12844 3928 12884 3968
rect 13228 3928 13268 3968
rect 13612 3928 13652 3968
rect 13996 3928 14036 3968
rect 14380 3928 14420 3968
rect 14764 3928 14804 3968
rect 15148 3928 15188 3968
rect 15532 3928 15572 3968
rect 15916 3928 15956 3968
rect 16300 3928 16340 3968
rect 16684 3928 16724 3968
rect 17356 3928 17396 3968
rect 17932 3928 17972 3968
rect 18316 3928 18356 3968
rect 18700 3928 18740 3968
rect 19756 3928 19796 3968
rect 19948 3928 19988 3968
rect 20524 3928 20564 3968
rect 20908 3928 20948 3968
rect 21484 3928 21524 3968
rect 21868 3928 21908 3968
rect 23212 3928 23252 3968
rect 23596 3928 23636 3968
rect 24556 3928 24596 3968
rect 25516 3928 25556 3968
rect 25900 3928 25940 3968
rect 26284 3928 26324 3968
rect 26668 3928 26708 3968
rect 27052 3928 27092 3968
rect 27436 3928 27476 3968
rect 27628 3928 27668 3968
rect 28588 3928 28628 3968
rect 28972 3928 29012 3968
rect 30124 3928 30164 3968
rect 30316 3928 30356 3968
rect 31660 3928 31700 3968
rect 32044 3928 32084 3968
rect 32428 3928 32468 3968
rect 32812 3928 32852 3968
rect 33196 3928 33236 3968
rect 33580 3928 33620 3968
rect 36268 3928 36308 3968
rect 36652 3928 36692 3968
rect 37036 3928 37076 3968
rect 37420 3928 37460 3968
rect 37804 3928 37844 3968
rect 38188 3928 38228 3968
rect 38956 3928 38996 3968
rect 39340 3928 39380 3968
rect 39724 3928 39764 3968
rect 40108 3928 40148 3968
rect 40492 3928 40532 3968
rect 40876 3928 40916 3968
rect 41260 3928 41300 3968
rect 41644 3928 41684 3968
rect 42028 3928 42068 3968
rect 42412 3928 42452 3968
rect 43180 3928 43220 3968
rect 43564 3928 43604 3968
rect 44236 3928 44276 3968
rect 46732 3928 46772 3968
rect 49228 3928 49268 3968
rect 49708 3928 49748 3968
rect 50668 3928 50708 3968
rect 51052 3928 51092 3968
rect 52396 3928 52436 3968
rect 53356 3928 53396 3968
rect 53740 3928 53780 3968
rect 54124 3928 54164 3968
rect 55468 3928 55508 3968
rect 55852 3928 55892 3968
rect 57196 3928 57236 3968
rect 57388 3928 57428 3968
rect 61420 3928 61460 3968
rect 61804 3928 61844 3968
rect 62188 3928 62228 3968
rect 62572 3928 62612 3968
rect 65068 3928 65108 3968
rect 65452 3928 65492 3968
rect 65836 3928 65876 3968
rect 66220 3928 66260 3968
rect 67372 3928 67412 3968
rect 67756 3928 67796 3968
rect 68140 3928 68180 3968
rect 69292 3928 69332 3968
rect 69676 3928 69716 3968
rect 70252 3928 70292 3968
rect 71788 3928 71828 3968
rect 72172 3928 72212 3968
rect 72364 3928 72404 3968
rect 73324 3928 73364 3968
rect 73708 3928 73748 3968
rect 73900 3928 73940 3968
rect 74284 3928 74324 3968
rect 75052 3928 75092 3968
rect 75436 3928 75476 3968
rect 76012 3928 76052 3968
rect 76204 3928 76244 3968
rect 76780 3928 76820 3968
rect 78796 3928 78836 3968
rect 79180 3928 79220 3968
rect 79564 3928 79604 3968
rect 79948 3928 79988 3968
rect 80332 3928 80372 3968
rect 80908 3928 80948 3968
rect 82444 3928 82484 3968
rect 82828 3928 82868 3968
rect 83404 3928 83444 3968
rect 83596 3928 83636 3968
rect 85708 3928 85748 3968
rect 86476 3928 86516 3968
rect 86860 3928 86900 3968
rect 87244 3928 87284 3968
rect 87628 3928 87668 3968
rect 88012 3928 88052 3968
rect 88396 3928 88436 3968
rect 88780 3928 88820 3968
rect 89164 3928 89204 3968
rect 89548 3928 89588 3968
rect 89932 3928 89972 3968
rect 90316 3928 90356 3968
rect 90700 3928 90740 3968
rect 91084 3928 91124 3968
rect 91468 3928 91508 3968
rect 91852 3928 91892 3968
rect 92236 3928 92276 3968
rect 92620 3928 92660 3968
rect 93004 3928 93044 3968
rect 93388 3928 93428 3968
rect 93772 3928 93812 3968
rect 94156 3928 94196 3968
rect 94540 3928 94580 3968
rect 95308 3928 95348 3968
rect 95692 3928 95732 3968
rect 96076 3928 96116 3968
rect 96460 3928 96500 3968
rect 96844 3928 96884 3968
rect 97228 3928 97268 3968
rect 97612 3928 97652 3968
rect 97996 3928 98036 3968
rect 98380 3928 98420 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 64168 3760 64208 3800
rect 64250 3760 64290 3800
rect 64332 3760 64372 3800
rect 64414 3760 64454 3800
rect 64496 3760 64536 3800
rect 79288 3760 79328 3800
rect 79370 3760 79410 3800
rect 79452 3760 79492 3800
rect 79534 3760 79574 3800
rect 79616 3760 79656 3800
rect 94408 3760 94448 3800
rect 94490 3760 94530 3800
rect 94572 3760 94612 3800
rect 94654 3760 94694 3800
rect 94736 3760 94776 3800
rect 49804 3592 49844 3632
rect 65356 3592 65396 3632
rect 81772 3592 81812 3632
rect 85132 3592 85172 3632
rect 49612 3508 49652 3548
rect 50092 3508 50132 3548
rect 50284 3508 50324 3548
rect 52492 3508 52532 3548
rect 52684 3508 52724 3548
rect 54796 3508 54836 3548
rect 57292 3508 57332 3548
rect 60268 3508 60308 3548
rect 64972 3508 65012 3548
rect 82636 3508 82676 3548
rect 1228 3424 1268 3464
rect 1612 3424 1652 3464
rect 1996 3424 2036 3464
rect 2380 3424 2420 3464
rect 2764 3424 2804 3464
rect 3148 3424 3188 3464
rect 3532 3424 3572 3464
rect 3916 3424 3956 3464
rect 4300 3424 4340 3464
rect 4684 3424 4724 3464
rect 5068 3424 5108 3464
rect 5452 3424 5492 3464
rect 5836 3424 5876 3464
rect 6220 3424 6260 3464
rect 6604 3424 6644 3464
rect 6988 3424 7028 3464
rect 7372 3424 7412 3464
rect 7756 3424 7796 3464
rect 8140 3424 8180 3464
rect 8524 3424 8564 3464
rect 8908 3424 8948 3464
rect 9292 3424 9332 3464
rect 9676 3424 9716 3464
rect 10060 3424 10100 3464
rect 10444 3424 10484 3464
rect 10828 3424 10868 3464
rect 11212 3424 11252 3464
rect 11596 3424 11636 3464
rect 11980 3424 12020 3464
rect 12364 3424 12404 3464
rect 12748 3424 12788 3464
rect 13132 3424 13172 3464
rect 13516 3424 13556 3464
rect 13900 3424 13940 3464
rect 14284 3424 14324 3464
rect 14668 3424 14708 3464
rect 15052 3424 15092 3464
rect 15436 3424 15476 3464
rect 15820 3424 15860 3464
rect 16204 3424 16244 3464
rect 16588 3424 16628 3464
rect 16972 3424 17012 3464
rect 17356 3424 17396 3464
rect 18508 3424 18548 3464
rect 18892 3424 18932 3464
rect 19276 3424 19316 3464
rect 19660 3424 19700 3464
rect 20044 3424 20084 3464
rect 20428 3424 20468 3464
rect 20812 3424 20852 3464
rect 21196 3424 21236 3464
rect 21580 3424 21620 3464
rect 21964 3424 22004 3464
rect 22348 3424 22388 3464
rect 22732 3424 22772 3464
rect 23116 3424 23156 3464
rect 23500 3424 23540 3464
rect 23884 3424 23924 3464
rect 24268 3424 24308 3464
rect 24652 3424 24692 3464
rect 25036 3424 25076 3464
rect 25420 3424 25460 3464
rect 25804 3424 25844 3464
rect 26188 3424 26228 3464
rect 26572 3424 26612 3464
rect 26956 3424 26996 3464
rect 27340 3424 27380 3464
rect 27724 3424 27764 3464
rect 28108 3424 28148 3464
rect 28492 3424 28532 3464
rect 28876 3424 28916 3464
rect 29260 3424 29300 3464
rect 29644 3424 29684 3464
rect 30028 3424 30068 3464
rect 30412 3424 30452 3464
rect 30796 3424 30836 3464
rect 31180 3424 31220 3464
rect 31564 3424 31604 3464
rect 31948 3424 31988 3464
rect 32332 3424 32372 3464
rect 32716 3424 32756 3464
rect 33100 3424 33140 3464
rect 33484 3424 33524 3464
rect 33868 3424 33908 3464
rect 34252 3424 34292 3464
rect 35308 3424 35348 3464
rect 35692 3424 35732 3464
rect 36076 3424 36116 3464
rect 36460 3424 36500 3464
rect 36844 3424 36884 3464
rect 37228 3424 37268 3464
rect 37612 3424 37652 3464
rect 37996 3424 38036 3464
rect 38380 3424 38420 3464
rect 38764 3424 38804 3464
rect 39148 3424 39188 3464
rect 39532 3424 39572 3464
rect 39916 3424 39956 3464
rect 40300 3424 40340 3464
rect 40684 3424 40724 3464
rect 41068 3424 41108 3464
rect 41452 3424 41492 3464
rect 41836 3424 41876 3464
rect 42220 3424 42260 3464
rect 42604 3424 42644 3464
rect 42988 3424 43028 3464
rect 43372 3424 43412 3464
rect 43756 3424 43796 3464
rect 44140 3424 44180 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 45292 3424 45332 3464
rect 45676 3424 45716 3464
rect 47980 3424 48020 3464
rect 48364 3424 48404 3464
rect 48748 3424 48788 3464
rect 50476 3424 50516 3464
rect 50860 3424 50900 3464
rect 51436 3424 51476 3464
rect 51820 3424 51860 3464
rect 52204 3424 52244 3464
rect 53164 3424 53204 3464
rect 53548 3424 53588 3464
rect 53932 3424 53972 3464
rect 54316 3424 54356 3464
rect 55276 3424 55316 3464
rect 55660 3424 55700 3464
rect 56044 3424 56084 3464
rect 56428 3424 56468 3464
rect 56812 3424 56852 3464
rect 57772 3424 57812 3464
rect 58156 3424 58196 3464
rect 58540 3424 58580 3464
rect 58924 3424 58964 3464
rect 60748 3424 60788 3464
rect 61132 3424 61172 3464
rect 61516 3424 61556 3464
rect 61900 3424 61940 3464
rect 62284 3424 62324 3464
rect 63244 3424 63284 3464
rect 63628 3424 63668 3464
rect 64012 3424 64052 3464
rect 64396 3424 64436 3464
rect 64780 3424 64820 3464
rect 65164 3424 65204 3464
rect 65548 3424 65588 3464
rect 65932 3424 65972 3464
rect 66316 3424 66356 3464
rect 66700 3424 66740 3464
rect 67084 3424 67124 3464
rect 67468 3424 67508 3464
rect 67852 3424 67892 3464
rect 68236 3424 68276 3464
rect 68620 3424 68660 3464
rect 69004 3424 69044 3464
rect 69388 3424 69428 3464
rect 69772 3424 69812 3464
rect 70156 3424 70196 3464
rect 70550 3411 70590 3451
rect 70924 3424 70964 3464
rect 71308 3424 71348 3464
rect 71692 3424 71732 3464
rect 72076 3424 72116 3464
rect 72460 3424 72500 3464
rect 72844 3424 72884 3464
rect 73228 3424 73268 3464
rect 73612 3424 73652 3464
rect 73996 3424 74036 3464
rect 74380 3424 74420 3464
rect 74764 3424 74804 3464
rect 75148 3424 75188 3464
rect 75532 3424 75572 3464
rect 75916 3435 75956 3475
rect 76300 3424 76340 3464
rect 76684 3424 76724 3464
rect 77068 3424 77108 3464
rect 77452 3424 77492 3464
rect 77836 3424 77876 3464
rect 78220 3424 78260 3464
rect 78604 3424 78644 3464
rect 78988 3424 79028 3464
rect 79372 3424 79412 3464
rect 79756 3424 79796 3464
rect 80140 3424 80180 3464
rect 80524 3424 80564 3464
rect 82444 3424 82484 3464
rect 82828 3424 82868 3464
rect 83212 3424 83252 3464
rect 83596 3424 83636 3464
rect 83980 3424 84020 3464
rect 84364 3424 84404 3464
rect 84748 3424 84788 3464
rect 85516 3424 85556 3464
rect 85900 3424 85940 3464
rect 86284 3424 86324 3464
rect 86668 3424 86708 3464
rect 87052 3424 87092 3464
rect 87436 3424 87476 3464
rect 87820 3424 87860 3464
rect 88204 3424 88244 3464
rect 88588 3424 88628 3464
rect 88972 3424 89012 3464
rect 89356 3424 89396 3464
rect 89740 3424 89780 3464
rect 90124 3424 90164 3464
rect 90508 3424 90548 3464
rect 90892 3424 90932 3464
rect 91276 3424 91316 3464
rect 91660 3424 91700 3464
rect 92044 3424 92084 3464
rect 92428 3424 92468 3464
rect 92812 3424 92852 3464
rect 93196 3424 93236 3464
rect 93580 3424 93620 3464
rect 93964 3424 94004 3464
rect 94348 3424 94388 3464
rect 94732 3424 94772 3464
rect 95116 3424 95156 3464
rect 95500 3424 95540 3464
rect 95884 3424 95924 3464
rect 96268 3424 96308 3464
rect 96652 3424 96692 3464
rect 97036 3424 97076 3464
rect 97420 3424 97460 3464
rect 97804 3424 97844 3464
rect 98188 3424 98228 3464
rect 98572 3424 98612 3464
rect 17740 3340 17780 3380
rect 17932 3340 17972 3380
rect 34732 3340 34772 3380
rect 34924 3340 34964 3380
rect 46060 3340 46100 3380
rect 46252 3340 46292 3380
rect 46348 3340 46388 3380
rect 47500 3340 47540 3380
rect 49132 3340 49172 3380
rect 49324 3340 49364 3380
rect 49612 3340 49652 3380
rect 50092 3340 50132 3380
rect 52684 3340 52724 3380
rect 54796 3340 54836 3380
rect 57292 3340 57332 3380
rect 59500 3340 59540 3380
rect 59692 3340 59732 3380
rect 60076 3340 60116 3380
rect 60268 3340 60308 3380
rect 62572 3340 62612 3380
rect 62764 3340 62804 3380
rect 81196 3340 81236 3380
rect 84940 3340 84980 3380
rect 85132 3340 85172 3380
rect 46636 3256 46676 3296
rect 49228 3256 49268 3296
rect 1420 3172 1460 3212
rect 1804 3172 1844 3212
rect 2188 3172 2228 3212
rect 2572 3172 2612 3212
rect 2956 3172 2996 3212
rect 3340 3172 3380 3212
rect 3724 3172 3764 3212
rect 4108 3172 4148 3212
rect 4492 3172 4532 3212
rect 4876 3172 4916 3212
rect 5260 3172 5300 3212
rect 5644 3172 5684 3212
rect 6028 3172 6068 3212
rect 6412 3172 6452 3212
rect 6796 3172 6836 3212
rect 7180 3172 7220 3212
rect 7564 3172 7604 3212
rect 7948 3172 7988 3212
rect 8332 3172 8372 3212
rect 8716 3172 8756 3212
rect 9100 3172 9140 3212
rect 9484 3172 9524 3212
rect 9868 3172 9908 3212
rect 10252 3172 10292 3212
rect 10636 3172 10676 3212
rect 11020 3172 11060 3212
rect 11404 3172 11444 3212
rect 11788 3172 11828 3212
rect 12172 3172 12212 3212
rect 12556 3172 12596 3212
rect 12940 3172 12980 3212
rect 13324 3172 13364 3212
rect 13708 3172 13748 3212
rect 14092 3172 14132 3212
rect 14476 3172 14516 3212
rect 14860 3172 14900 3212
rect 15244 3172 15284 3212
rect 15628 3172 15668 3212
rect 16012 3172 16052 3212
rect 16396 3172 16436 3212
rect 16780 3172 16820 3212
rect 17164 3172 17204 3212
rect 17548 3172 17588 3212
rect 18700 3172 18740 3212
rect 19084 3172 19124 3212
rect 19468 3172 19508 3212
rect 19852 3172 19892 3212
rect 20236 3172 20276 3212
rect 20620 3172 20660 3212
rect 21004 3172 21044 3212
rect 21388 3172 21428 3212
rect 21772 3172 21812 3212
rect 22156 3172 22196 3212
rect 22540 3172 22580 3212
rect 22924 3172 22964 3212
rect 23308 3172 23348 3212
rect 23692 3172 23732 3212
rect 24076 3172 24116 3212
rect 24460 3172 24500 3212
rect 24844 3172 24884 3212
rect 25228 3172 25268 3212
rect 25612 3172 25652 3212
rect 25996 3172 26036 3212
rect 26380 3172 26420 3212
rect 26764 3172 26804 3212
rect 27148 3172 27188 3212
rect 27532 3172 27572 3212
rect 27916 3172 27956 3212
rect 28300 3172 28340 3212
rect 28684 3172 28724 3212
rect 29068 3172 29108 3212
rect 29452 3172 29492 3212
rect 29836 3172 29876 3212
rect 30220 3172 30260 3212
rect 30604 3172 30644 3212
rect 30988 3172 31028 3212
rect 31372 3172 31412 3212
rect 31756 3172 31796 3212
rect 32140 3172 32180 3212
rect 32524 3172 32564 3212
rect 32908 3172 32948 3212
rect 33292 3172 33332 3212
rect 33676 3172 33716 3212
rect 34060 3172 34100 3212
rect 34444 3172 34484 3212
rect 34924 3172 34964 3212
rect 35500 3172 35540 3212
rect 35884 3172 35924 3212
rect 36268 3172 36308 3212
rect 36652 3172 36692 3212
rect 37036 3172 37076 3212
rect 37420 3172 37460 3212
rect 37804 3172 37844 3212
rect 38188 3172 38228 3212
rect 38572 3172 38612 3212
rect 38956 3172 38996 3212
rect 39340 3172 39380 3212
rect 39724 3172 39764 3212
rect 40108 3172 40148 3212
rect 40492 3172 40532 3212
rect 40876 3172 40916 3212
rect 41260 3172 41300 3212
rect 41644 3172 41684 3212
rect 42028 3172 42068 3212
rect 42412 3172 42452 3212
rect 42796 3172 42836 3212
rect 43180 3172 43220 3212
rect 43564 3172 43604 3212
rect 43948 3172 43988 3212
rect 44332 3172 44372 3212
rect 44716 3172 44756 3212
rect 45100 3172 45140 3212
rect 45484 3172 45524 3212
rect 45868 3172 45908 3212
rect 46060 3172 46100 3212
rect 48172 3172 48212 3212
rect 48556 3172 48596 3212
rect 48940 3172 48980 3212
rect 50668 3172 50708 3212
rect 51052 3172 51092 3212
rect 51244 3172 51284 3212
rect 51628 3172 51668 3212
rect 52012 3172 52052 3212
rect 52972 3172 53012 3212
rect 53356 3172 53396 3212
rect 53740 3172 53780 3212
rect 54124 3172 54164 3212
rect 54604 3172 54644 3212
rect 55084 3172 55124 3212
rect 55468 3172 55508 3212
rect 55852 3172 55892 3212
rect 56236 3172 56276 3212
rect 56620 3172 56660 3212
rect 57100 3172 57140 3212
rect 57580 3172 57620 3212
rect 57964 3172 58004 3212
rect 58348 3172 58388 3212
rect 58732 3172 58772 3212
rect 59500 3172 59540 3212
rect 60556 3172 60596 3212
rect 60940 3172 60980 3212
rect 61324 3172 61364 3212
rect 61708 3172 61748 3212
rect 62092 3172 62132 3212
rect 63052 3172 63092 3212
rect 63436 3172 63476 3212
rect 63820 3172 63860 3212
rect 64204 3172 64244 3212
rect 64588 3172 64628 3212
rect 65740 3172 65780 3212
rect 66124 3172 66164 3212
rect 66508 3172 66548 3212
rect 66892 3172 66932 3212
rect 67276 3172 67316 3212
rect 67660 3172 67700 3212
rect 68044 3172 68084 3212
rect 68428 3172 68468 3212
rect 68812 3172 68852 3212
rect 69196 3172 69236 3212
rect 69580 3172 69620 3212
rect 69964 3172 70004 3212
rect 70348 3172 70388 3212
rect 70732 3172 70772 3212
rect 71116 3172 71156 3212
rect 71500 3172 71540 3212
rect 71884 3172 71924 3212
rect 72268 3172 72308 3212
rect 72652 3172 72692 3212
rect 73036 3172 73076 3212
rect 73420 3172 73460 3212
rect 73804 3172 73844 3212
rect 74188 3172 74228 3212
rect 74572 3172 74612 3212
rect 74956 3172 74996 3212
rect 75340 3172 75380 3212
rect 75724 3172 75764 3212
rect 76108 3172 76148 3212
rect 76492 3172 76532 3212
rect 76876 3172 76916 3212
rect 77260 3172 77300 3212
rect 77644 3172 77684 3212
rect 78028 3172 78068 3212
rect 78412 3172 78452 3212
rect 78796 3172 78836 3212
rect 79180 3172 79220 3212
rect 79564 3172 79604 3212
rect 79948 3172 79988 3212
rect 80332 3172 80372 3212
rect 82252 3172 82292 3212
rect 83020 3172 83060 3212
rect 83404 3172 83444 3212
rect 83788 3172 83828 3212
rect 84172 3172 84212 3212
rect 84556 3172 84596 3212
rect 85324 3172 85364 3212
rect 85708 3172 85748 3212
rect 86092 3172 86132 3212
rect 86476 3172 86516 3212
rect 86860 3172 86900 3212
rect 87244 3172 87284 3212
rect 87628 3172 87668 3212
rect 88012 3172 88052 3212
rect 88396 3172 88436 3212
rect 88780 3172 88820 3212
rect 89164 3172 89204 3212
rect 89548 3172 89588 3212
rect 89932 3172 89972 3212
rect 90316 3172 90356 3212
rect 90700 3172 90740 3212
rect 91084 3172 91124 3212
rect 91468 3172 91508 3212
rect 91852 3172 91892 3212
rect 92236 3172 92276 3212
rect 92620 3172 92660 3212
rect 93004 3172 93044 3212
rect 93388 3172 93428 3212
rect 93772 3172 93812 3212
rect 94156 3172 94196 3212
rect 94540 3172 94580 3212
rect 94924 3172 94964 3212
rect 95308 3172 95348 3212
rect 95692 3172 95732 3212
rect 96076 3172 96116 3212
rect 96460 3172 96500 3212
rect 96844 3172 96884 3212
rect 97228 3172 97268 3212
rect 97612 3172 97652 3212
rect 97996 3172 98036 3212
rect 98380 3172 98420 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 65408 3004 65448 3044
rect 65490 3004 65530 3044
rect 65572 3004 65612 3044
rect 65654 3004 65694 3044
rect 65736 3004 65776 3044
rect 80528 3004 80568 3044
rect 80610 3004 80650 3044
rect 80692 3004 80732 3044
rect 80774 3004 80814 3044
rect 80856 3004 80896 3044
rect 95648 3004 95688 3044
rect 95730 3004 95770 3044
rect 95812 3004 95852 3044
rect 95894 3004 95934 3044
rect 95976 3004 96016 3044
<< metal2 >>
rect 6200 14920 6280 15000
rect 17144 14920 17224 15000
rect 28088 14920 28168 15000
rect 39032 14920 39112 15000
rect 49976 14920 50056 15000
rect 60920 14920 61000 15000
rect 71864 14920 71944 15000
rect 82808 14920 82888 15000
rect 93752 14920 93832 15000
rect 6220 11957 6260 14920
rect 6219 11948 6261 11957
rect 6219 11908 6220 11948
rect 6260 11908 6261 11948
rect 6219 11899 6261 11908
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 17164 11360 17204 14920
rect 18808 11360 19176 11369
rect 17164 11320 17300 11360
rect 3688 11311 4056 11320
rect 11884 11192 11924 11201
rect 11924 11152 12500 11192
rect 11884 11143 11924 11152
rect 11979 11024 12021 11033
rect 11979 10984 11980 11024
rect 12020 10984 12021 11024
rect 11979 10975 12021 10984
rect 11788 10940 11828 10949
rect 10731 10856 10773 10865
rect 10731 10816 10732 10856
rect 10772 10816 10773 10856
rect 10731 10807 10773 10816
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 7371 10184 7413 10193
rect 7371 10144 7372 10184
rect 7412 10144 7413 10184
rect 7371 10135 7413 10144
rect 3435 10016 3477 10025
rect 3435 9976 3436 10016
rect 3476 9976 3477 10016
rect 3435 9967 3477 9976
rect 3051 8840 3093 8849
rect 3051 8800 3052 8840
rect 3092 8800 3093 8840
rect 3051 8791 3093 8800
rect 1995 8168 2037 8177
rect 1995 8128 1996 8168
rect 2036 8128 2037 8168
rect 1995 8119 2037 8128
rect 1419 6488 1461 6497
rect 1419 6448 1420 6488
rect 1460 6448 1461 6488
rect 1419 6439 1461 6448
rect 1420 6354 1460 6439
rect 1228 6236 1268 6245
rect 844 6196 1228 6236
rect 844 80 884 6196
rect 1228 6187 1268 6196
rect 1707 5648 1749 5657
rect 1707 5608 1708 5648
rect 1748 5608 1749 5648
rect 1707 5599 1749 5608
rect 1708 5514 1748 5599
rect 1131 5480 1173 5489
rect 1516 5480 1556 5489
rect 1131 5440 1132 5480
rect 1172 5440 1173 5480
rect 1131 5431 1173 5440
rect 1324 5440 1516 5480
rect 1035 3380 1077 3389
rect 1035 3340 1036 3380
rect 1076 3340 1077 3380
rect 1035 3331 1077 3340
rect 1036 80 1076 3331
rect 1132 2792 1172 5431
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1228 3330 1268 3415
rect 1324 2792 1364 5440
rect 1516 5431 1556 5440
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 1900 5346 1940 5431
rect 1708 4976 1748 4985
rect 1611 4892 1653 4901
rect 1611 4852 1612 4892
rect 1652 4852 1653 4892
rect 1611 4843 1653 4852
rect 1516 4724 1556 4733
rect 1420 4684 1516 4724
rect 1420 3380 1460 4684
rect 1516 4675 1556 4684
rect 1516 4136 1556 4145
rect 1612 4136 1652 4843
rect 1708 4817 1748 4936
rect 1707 4808 1749 4817
rect 1707 4768 1708 4808
rect 1748 4768 1749 4808
rect 1707 4759 1749 4768
rect 1900 4724 1940 4733
rect 1556 4096 1652 4136
rect 1804 4684 1900 4724
rect 1516 4087 1556 4096
rect 1708 3968 1748 3977
rect 1612 3473 1652 3558
rect 1611 3464 1653 3473
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 1420 3340 1556 3380
rect 1419 3212 1461 3221
rect 1419 3172 1420 3212
rect 1460 3172 1461 3212
rect 1419 3163 1461 3172
rect 1420 3078 1460 3163
rect 1132 2752 1268 2792
rect 1324 2752 1460 2792
rect 1228 80 1268 2752
rect 1420 80 1460 2752
rect 1516 2372 1556 3340
rect 1611 3212 1653 3221
rect 1611 3172 1612 3212
rect 1652 3172 1653 3212
rect 1611 3163 1653 3172
rect 1612 2549 1652 3163
rect 1611 2540 1653 2549
rect 1611 2500 1612 2540
rect 1652 2500 1653 2540
rect 1611 2491 1653 2500
rect 1516 2332 1652 2372
rect 1612 80 1652 2332
rect 1708 2045 1748 3928
rect 1804 3380 1844 4684
rect 1900 4675 1940 4684
rect 1900 4136 1940 4145
rect 1996 4136 2036 8119
rect 2379 7748 2421 7757
rect 2379 7708 2380 7748
rect 2420 7708 2421 7748
rect 2379 7699 2421 7708
rect 2091 5648 2133 5657
rect 2091 5608 2092 5648
rect 2132 5608 2133 5648
rect 2091 5599 2133 5608
rect 2092 5514 2132 5599
rect 2091 4976 2133 4985
rect 2091 4936 2092 4976
rect 2132 4936 2133 4976
rect 2091 4927 2133 4936
rect 2092 4842 2132 4927
rect 2284 4724 2324 4733
rect 1940 4096 2036 4136
rect 2188 4684 2284 4724
rect 1900 4087 1940 4096
rect 2092 3968 2132 3977
rect 1995 3464 2037 3473
rect 1995 3424 1996 3464
rect 2036 3424 2037 3464
rect 1995 3415 2037 3424
rect 1804 3340 1940 3380
rect 1804 3212 1844 3221
rect 1804 2549 1844 3172
rect 1803 2540 1845 2549
rect 1803 2500 1804 2540
rect 1844 2500 1845 2540
rect 1803 2491 1845 2500
rect 1900 2372 1940 3340
rect 1996 3330 2036 3415
rect 1804 2332 1940 2372
rect 1707 2036 1749 2045
rect 1707 1996 1708 2036
rect 1748 1996 1749 2036
rect 1707 1987 1749 1996
rect 1804 80 1844 2332
rect 1995 2036 2037 2045
rect 1995 1996 1996 2036
rect 2036 1996 2037 2036
rect 1995 1987 2037 1996
rect 1996 80 2036 1987
rect 2092 1961 2132 3928
rect 2188 3380 2228 4684
rect 2284 4675 2324 4684
rect 2284 4136 2324 4145
rect 2380 4136 2420 7699
rect 2763 6404 2805 6413
rect 2763 6364 2764 6404
rect 2804 6364 2805 6404
rect 2763 6355 2805 6364
rect 2475 4976 2517 4985
rect 2475 4936 2476 4976
rect 2516 4936 2517 4976
rect 2475 4927 2517 4936
rect 2476 4842 2516 4927
rect 2668 4724 2708 4733
rect 2324 4096 2420 4136
rect 2572 4684 2668 4724
rect 2284 4087 2324 4096
rect 2476 3968 2516 3977
rect 2380 3473 2420 3558
rect 2379 3464 2421 3473
rect 2379 3424 2380 3464
rect 2420 3424 2421 3464
rect 2379 3415 2421 3424
rect 2188 3340 2324 3380
rect 2187 3212 2229 3221
rect 2187 3172 2188 3212
rect 2228 3172 2229 3212
rect 2187 3163 2229 3172
rect 2188 3078 2228 3163
rect 2284 2372 2324 3340
rect 2379 3212 2421 3221
rect 2379 3172 2380 3212
rect 2420 3172 2421 3212
rect 2379 3163 2421 3172
rect 2188 2332 2324 2372
rect 2091 1952 2133 1961
rect 2091 1912 2092 1952
rect 2132 1912 2133 1952
rect 2091 1903 2133 1912
rect 2188 80 2228 2332
rect 2380 2129 2420 3163
rect 2476 2540 2516 3928
rect 2572 3389 2612 4684
rect 2668 4675 2708 4684
rect 2667 4220 2709 4229
rect 2667 4180 2668 4220
rect 2708 4180 2709 4220
rect 2667 4171 2709 4180
rect 2668 4136 2708 4171
rect 2668 4085 2708 4096
rect 2764 3464 2804 6355
rect 2860 4976 2900 4985
rect 2900 4936 2996 4976
rect 2860 4927 2900 4936
rect 2764 3415 2804 3424
rect 2860 3968 2900 3977
rect 2571 3380 2613 3389
rect 2571 3340 2572 3380
rect 2612 3340 2613 3380
rect 2571 3331 2613 3340
rect 2571 3212 2613 3221
rect 2571 3172 2572 3212
rect 2612 3172 2613 3212
rect 2571 3163 2613 3172
rect 2572 3078 2612 3163
rect 2476 2500 2804 2540
rect 2571 2372 2613 2381
rect 2571 2332 2572 2372
rect 2612 2332 2613 2372
rect 2571 2323 2613 2332
rect 2379 2120 2421 2129
rect 2379 2080 2380 2120
rect 2420 2080 2421 2120
rect 2379 2071 2421 2080
rect 2379 1952 2421 1961
rect 2379 1912 2380 1952
rect 2420 1912 2421 1952
rect 2379 1903 2421 1912
rect 2380 80 2420 1903
rect 2572 80 2612 2323
rect 2764 80 2804 2500
rect 2860 1205 2900 3928
rect 2956 3380 2996 4936
rect 3052 4136 3092 8791
rect 3147 6656 3189 6665
rect 3147 6616 3148 6656
rect 3188 6616 3189 6656
rect 3147 6607 3189 6616
rect 3052 4087 3092 4096
rect 3148 3464 3188 6607
rect 3339 5480 3381 5489
rect 3339 5440 3340 5480
rect 3380 5440 3381 5480
rect 3339 5431 3381 5440
rect 3148 3415 3188 3424
rect 3244 3968 3284 3977
rect 2956 3340 3092 3380
rect 3052 3296 3092 3340
rect 3052 3256 3188 3296
rect 2956 3212 2996 3221
rect 2996 3172 3092 3212
rect 2956 3163 2996 3172
rect 2955 2540 2997 2549
rect 2955 2500 2956 2540
rect 2996 2500 2997 2540
rect 2955 2491 2997 2500
rect 2859 1196 2901 1205
rect 2859 1156 2860 1196
rect 2900 1156 2901 1196
rect 2859 1147 2901 1156
rect 2956 80 2996 2491
rect 3052 1289 3092 3172
rect 3148 1457 3188 3256
rect 3244 3137 3284 3928
rect 3340 3473 3380 5431
rect 3436 4136 3476 9967
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 6219 9512 6261 9521
rect 6219 9472 6220 9512
rect 6260 9472 6261 9512
rect 6219 9463 6261 9472
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 6123 8756 6165 8765
rect 6123 8716 6124 8756
rect 6164 8716 6165 8756
rect 6123 8707 6165 8716
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5355 7160 5397 7169
rect 5355 7120 5356 7160
rect 5396 7120 5397 7160
rect 5355 7111 5397 7120
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4779 6152 4821 6161
rect 4779 6112 4780 6152
rect 4820 6112 4821 6152
rect 4779 6103 4821 6112
rect 4107 5732 4149 5741
rect 4107 5692 4108 5732
rect 4148 5692 4149 5732
rect 4107 5683 4149 5692
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3819 5144 3861 5153
rect 3819 5104 3820 5144
rect 3860 5104 3861 5144
rect 3819 5095 3861 5104
rect 3436 4087 3476 4096
rect 3820 4136 3860 5095
rect 3820 4087 3860 4096
rect 4012 3977 4052 4062
rect 3628 3968 3668 3977
rect 3532 3928 3628 3968
rect 3532 3632 3572 3928
rect 3628 3919 3668 3928
rect 4011 3968 4053 3977
rect 4011 3928 4012 3968
rect 4052 3928 4053 3968
rect 4011 3919 4053 3928
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3532 3592 3860 3632
rect 3339 3464 3381 3473
rect 3339 3424 3340 3464
rect 3380 3424 3381 3464
rect 3339 3415 3381 3424
rect 3531 3464 3573 3473
rect 3531 3424 3532 3464
rect 3572 3424 3573 3464
rect 3531 3415 3573 3424
rect 3532 3330 3572 3415
rect 3340 3212 3380 3221
rect 3243 3128 3285 3137
rect 3243 3088 3244 3128
rect 3284 3088 3285 3128
rect 3243 3079 3285 3088
rect 3340 2540 3380 3172
rect 3627 3212 3669 3221
rect 3627 3172 3628 3212
rect 3668 3172 3669 3212
rect 3627 3163 3669 3172
rect 3724 3212 3764 3221
rect 3531 3128 3573 3137
rect 3531 3088 3532 3128
rect 3572 3088 3573 3128
rect 3531 3079 3573 3088
rect 3340 2500 3476 2540
rect 3339 2120 3381 2129
rect 3339 2080 3340 2120
rect 3380 2080 3381 2120
rect 3339 2071 3381 2080
rect 3147 1448 3189 1457
rect 3147 1408 3148 1448
rect 3188 1408 3189 1448
rect 3147 1399 3189 1408
rect 3051 1280 3093 1289
rect 3051 1240 3052 1280
rect 3092 1240 3093 1280
rect 3051 1231 3093 1240
rect 3147 1196 3189 1205
rect 3147 1156 3148 1196
rect 3188 1156 3189 1196
rect 3147 1147 3189 1156
rect 3148 80 3188 1147
rect 3340 80 3380 2071
rect 3436 1205 3476 2500
rect 3435 1196 3477 1205
rect 3435 1156 3436 1196
rect 3476 1156 3477 1196
rect 3435 1147 3477 1156
rect 3532 80 3572 3079
rect 3628 1364 3668 3163
rect 3724 1541 3764 3172
rect 3820 2036 3860 3592
rect 3916 3464 3956 3473
rect 4108 3464 4148 5683
rect 4203 5060 4245 5069
rect 4203 5020 4204 5060
rect 4244 5020 4245 5060
rect 4203 5011 4245 5020
rect 4204 4136 4244 5011
rect 4588 4145 4628 4230
rect 4204 4087 4244 4096
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4780 4136 4820 6103
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 5067 4388 5109 4397
rect 5067 4348 5068 4388
rect 5108 4348 5109 4388
rect 5067 4339 5109 4348
rect 4972 4136 5012 4145
rect 4780 4096 4972 4136
rect 4587 4087 4629 4096
rect 4972 4087 5012 4096
rect 4203 3968 4245 3977
rect 4203 3928 4204 3968
rect 4244 3928 4245 3968
rect 4203 3919 4245 3928
rect 4396 3968 4436 3977
rect 4780 3968 4820 3977
rect 4436 3928 4628 3968
rect 4396 3919 4436 3928
rect 3956 3424 4148 3464
rect 3916 3415 3956 3424
rect 4108 3212 4148 3221
rect 3820 1996 3956 2036
rect 3723 1532 3765 1541
rect 3723 1492 3724 1532
rect 3764 1492 3765 1532
rect 3723 1483 3765 1492
rect 3628 1324 3764 1364
rect 3724 80 3764 1324
rect 3916 80 3956 1996
rect 4108 1625 4148 3172
rect 4204 2036 4244 3919
rect 4299 3464 4341 3473
rect 4299 3424 4300 3464
rect 4340 3424 4341 3464
rect 4299 3415 4341 3424
rect 4300 3330 4340 3415
rect 4492 3212 4532 3221
rect 4204 1996 4340 2036
rect 4107 1616 4149 1625
rect 4107 1576 4108 1616
rect 4148 1576 4149 1616
rect 4107 1567 4149 1576
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 4108 80 4148 1231
rect 4300 80 4340 1996
rect 4492 1709 4532 3172
rect 4491 1700 4533 1709
rect 4491 1660 4492 1700
rect 4532 1660 4533 1700
rect 4491 1651 4533 1660
rect 4588 1616 4628 3928
rect 4683 3800 4725 3809
rect 4683 3760 4684 3800
rect 4724 3760 4725 3800
rect 4683 3751 4725 3760
rect 4684 3464 4724 3751
rect 4684 3415 4724 3424
rect 4683 3212 4725 3221
rect 4683 3172 4684 3212
rect 4724 3172 4725 3212
rect 4683 3163 4725 3172
rect 4684 1793 4724 3163
rect 4780 2036 4820 3928
rect 5068 3464 5108 4339
rect 5356 4136 5396 7111
rect 5739 6908 5781 6917
rect 5739 6868 5740 6908
rect 5780 6868 5781 6908
rect 5739 6859 5781 6868
rect 5451 6236 5493 6245
rect 5451 6196 5452 6236
rect 5492 6196 5493 6236
rect 5451 6187 5493 6196
rect 5452 4397 5492 6187
rect 5451 4388 5493 4397
rect 5451 4348 5452 4388
rect 5492 4348 5493 4388
rect 5451 4339 5493 4348
rect 5356 4087 5396 4096
rect 5740 4136 5780 6859
rect 5740 4087 5780 4096
rect 6124 4136 6164 8707
rect 6220 5069 6260 9463
rect 6507 6992 6549 7001
rect 6507 6952 6508 6992
rect 6548 6952 6549 6992
rect 6507 6943 6549 6952
rect 6219 5060 6261 5069
rect 6219 5020 6220 5060
rect 6260 5020 6261 5060
rect 6219 5011 6261 5020
rect 6124 4087 6164 4096
rect 6508 4136 6548 6943
rect 6891 6320 6933 6329
rect 6891 6280 6892 6320
rect 6932 6280 6933 6320
rect 6891 6271 6933 6280
rect 6508 4087 6548 4096
rect 6892 4136 6932 6271
rect 7372 6161 7412 10135
rect 7467 9932 7509 9941
rect 7467 9892 7468 9932
rect 7508 9892 7509 9932
rect 7467 9883 7509 9892
rect 7371 6152 7413 6161
rect 7371 6112 7372 6152
rect 7412 6112 7413 6152
rect 7371 6103 7413 6112
rect 7371 5396 7413 5405
rect 7371 5356 7372 5396
rect 7412 5356 7413 5396
rect 7371 5347 7413 5356
rect 7276 4145 7316 4230
rect 6892 4087 6932 4096
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 5164 3968 5204 3977
rect 5548 3968 5588 3977
rect 5204 3928 5396 3968
rect 5164 3919 5204 3928
rect 5068 3415 5108 3424
rect 4876 3221 4916 3306
rect 5260 3221 5300 3306
rect 4875 3212 4917 3221
rect 4875 3172 4876 3212
rect 4916 3172 4917 3212
rect 4875 3163 4917 3172
rect 5259 3212 5301 3221
rect 5259 3172 5260 3212
rect 5300 3172 5301 3212
rect 5259 3163 5301 3172
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 5356 2036 5396 3928
rect 5452 3464 5492 3473
rect 5452 2465 5492 3424
rect 5451 2456 5493 2465
rect 5451 2416 5452 2456
rect 5492 2416 5493 2456
rect 5451 2407 5493 2416
rect 4780 1996 5108 2036
rect 5356 1996 5492 2036
rect 4683 1784 4725 1793
rect 4683 1744 4684 1784
rect 4724 1744 4725 1784
rect 4683 1735 4725 1744
rect 4588 1576 4724 1616
rect 4491 1196 4533 1205
rect 4491 1156 4492 1196
rect 4532 1156 4533 1196
rect 4491 1147 4533 1156
rect 4492 80 4532 1147
rect 4684 80 4724 1576
rect 4875 1532 4917 1541
rect 4875 1492 4876 1532
rect 4916 1492 4917 1532
rect 4875 1483 4917 1492
rect 4876 80 4916 1483
rect 5068 80 5108 1996
rect 5259 1616 5301 1625
rect 5259 1576 5260 1616
rect 5300 1576 5301 1616
rect 5259 1567 5301 1576
rect 5260 80 5300 1567
rect 5452 80 5492 1996
rect 5548 1961 5588 3928
rect 5932 3968 5972 3977
rect 6316 3968 6356 3977
rect 6700 3968 6740 3977
rect 7084 3968 7124 3977
rect 5972 3928 6164 3968
rect 5932 3919 5972 3928
rect 5836 3464 5876 3473
rect 5644 3212 5684 3221
rect 5547 1952 5589 1961
rect 5547 1912 5548 1952
rect 5588 1912 5589 1952
rect 5547 1903 5589 1912
rect 5644 1877 5684 3172
rect 5739 3212 5781 3221
rect 5739 3172 5740 3212
rect 5780 3172 5781 3212
rect 5739 3163 5781 3172
rect 5740 2045 5780 3163
rect 5836 2381 5876 3424
rect 6028 3212 6068 3221
rect 5835 2372 5877 2381
rect 5835 2332 5836 2372
rect 5876 2332 5877 2372
rect 5835 2323 5877 2332
rect 5739 2036 5781 2045
rect 5739 1996 5740 2036
rect 5780 1996 5781 2036
rect 5739 1987 5781 1996
rect 6028 1961 6068 3172
rect 6124 2036 6164 3928
rect 6356 3928 6548 3968
rect 6316 3919 6356 3928
rect 6220 3464 6260 3473
rect 6220 2969 6260 3424
rect 6412 3212 6452 3221
rect 6219 2960 6261 2969
rect 6219 2920 6220 2960
rect 6260 2920 6261 2960
rect 6219 2911 6261 2920
rect 6412 2540 6452 3172
rect 6316 2500 6452 2540
rect 6124 1996 6260 2036
rect 5835 1952 5877 1961
rect 5835 1912 5836 1952
rect 5876 1912 5877 1952
rect 5835 1903 5877 1912
rect 6027 1952 6069 1961
rect 6027 1912 6028 1952
rect 6068 1912 6069 1952
rect 6027 1903 6069 1912
rect 5643 1868 5685 1877
rect 5643 1828 5644 1868
rect 5684 1828 5685 1868
rect 5643 1819 5685 1828
rect 5643 1700 5685 1709
rect 5643 1660 5644 1700
rect 5684 1660 5685 1700
rect 5643 1651 5685 1660
rect 5644 80 5684 1651
rect 5836 80 5876 1903
rect 6027 1784 6069 1793
rect 6027 1744 6028 1784
rect 6068 1744 6069 1784
rect 6027 1735 6069 1744
rect 6028 80 6068 1735
rect 6220 80 6260 1996
rect 6316 1709 6356 2500
rect 6411 2036 6453 2045
rect 6411 1996 6412 2036
rect 6452 1996 6453 2036
rect 6508 2036 6548 3928
rect 6740 3928 6932 3968
rect 6700 3919 6740 3928
rect 6604 3464 6644 3473
rect 6604 2540 6644 3424
rect 6796 3212 6836 3221
rect 6604 2500 6740 2540
rect 6508 1996 6644 2036
rect 6411 1987 6453 1996
rect 6315 1700 6357 1709
rect 6315 1660 6316 1700
rect 6356 1660 6357 1700
rect 6315 1651 6357 1660
rect 6412 80 6452 1987
rect 6604 80 6644 1996
rect 6700 1793 6740 2500
rect 6796 2045 6836 3172
rect 6795 2036 6837 2045
rect 6795 1996 6796 2036
rect 6836 1996 6837 2036
rect 6892 2036 6932 3928
rect 7124 3928 7316 3968
rect 7084 3919 7124 3928
rect 6987 3464 7029 3473
rect 6987 3424 6988 3464
rect 7028 3424 7029 3464
rect 6987 3415 7029 3424
rect 6988 3330 7028 3415
rect 7180 3212 7220 3221
rect 7180 2213 7220 3172
rect 7179 2204 7221 2213
rect 7179 2164 7180 2204
rect 7220 2164 7221 2204
rect 7179 2155 7221 2164
rect 6892 1996 7028 2036
rect 6795 1987 6837 1996
rect 6795 1868 6837 1877
rect 6795 1828 6796 1868
rect 6836 1828 6837 1868
rect 6795 1819 6837 1828
rect 6699 1784 6741 1793
rect 6699 1744 6700 1784
rect 6740 1744 6741 1784
rect 6699 1735 6741 1744
rect 6796 80 6836 1819
rect 6988 80 7028 1996
rect 7179 1952 7221 1961
rect 7179 1912 7180 1952
rect 7220 1912 7221 1952
rect 7276 1952 7316 3928
rect 7372 3809 7412 5347
rect 7468 5153 7508 9883
rect 9195 9428 9237 9437
rect 9195 9388 9196 9428
rect 9236 9388 9237 9428
rect 9195 9379 9237 9388
rect 7563 9008 7605 9017
rect 7563 8968 7564 9008
rect 7604 8968 7605 9008
rect 7563 8959 7605 8968
rect 7564 7757 7604 8959
rect 8811 8840 8853 8849
rect 8811 8800 8812 8840
rect 8852 8800 8853 8840
rect 8811 8791 8853 8800
rect 8427 8252 8469 8261
rect 8427 8212 8428 8252
rect 8468 8212 8469 8252
rect 8427 8203 8469 8212
rect 7563 7748 7605 7757
rect 7563 7708 7564 7748
rect 7604 7708 7605 7748
rect 7563 7699 7605 7708
rect 8043 7748 8085 7757
rect 8043 7708 8044 7748
rect 8084 7708 8085 7748
rect 8043 7699 8085 7708
rect 7467 5144 7509 5153
rect 7467 5104 7468 5144
rect 7508 5104 7509 5144
rect 7467 5095 7509 5104
rect 7659 4304 7701 4313
rect 7659 4264 7660 4304
rect 7700 4264 7701 4304
rect 7659 4255 7701 4264
rect 7660 4136 7700 4255
rect 7660 4087 7700 4096
rect 8044 4136 8084 7699
rect 8044 4087 8084 4096
rect 8428 4136 8468 8203
rect 8812 8177 8852 8791
rect 8811 8168 8853 8177
rect 8811 8128 8812 8168
rect 8852 8128 8853 8168
rect 8811 8119 8853 8128
rect 8907 7916 8949 7925
rect 8907 7876 8908 7916
rect 8948 7876 8949 7916
rect 8907 7867 8949 7876
rect 9100 7916 9140 7927
rect 8908 7782 8948 7867
rect 9100 7841 9140 7876
rect 9004 7832 9044 7841
rect 9004 6161 9044 7792
rect 9099 7832 9141 7841
rect 9099 7792 9100 7832
rect 9140 7792 9141 7832
rect 9099 7783 9141 7792
rect 9003 6152 9045 6161
rect 9003 6112 9004 6152
rect 9044 6112 9045 6152
rect 9003 6103 9045 6112
rect 8907 5312 8949 5321
rect 8907 5272 8908 5312
rect 8948 5272 8949 5312
rect 8907 5263 8949 5272
rect 8811 4976 8853 4985
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 8428 4087 8468 4096
rect 8812 4136 8852 4927
rect 8812 4087 8852 4096
rect 7468 3968 7508 3977
rect 7371 3800 7413 3809
rect 7371 3760 7372 3800
rect 7412 3760 7413 3800
rect 7371 3751 7413 3760
rect 7372 3464 7412 3473
rect 7372 3137 7412 3424
rect 7371 3128 7413 3137
rect 7371 3088 7372 3128
rect 7412 3088 7413 3128
rect 7371 3079 7413 3088
rect 7371 2960 7413 2969
rect 7371 2920 7372 2960
rect 7412 2920 7413 2960
rect 7371 2911 7413 2920
rect 7372 2129 7412 2911
rect 7371 2120 7413 2129
rect 7371 2080 7372 2120
rect 7412 2080 7413 2120
rect 7371 2071 7413 2080
rect 7468 2036 7508 3928
rect 7852 3968 7892 3977
rect 8236 3968 8276 3977
rect 7892 3928 8084 3968
rect 7852 3919 7892 3928
rect 7756 3464 7796 3473
rect 7756 3305 7796 3424
rect 7755 3296 7797 3305
rect 7755 3256 7756 3296
rect 7796 3256 7797 3296
rect 7755 3247 7797 3256
rect 7563 3212 7605 3221
rect 7563 3172 7564 3212
rect 7604 3172 7605 3212
rect 7563 3163 7605 3172
rect 7948 3212 7988 3221
rect 7564 3078 7604 3163
rect 7948 2381 7988 3172
rect 7947 2372 7989 2381
rect 7947 2332 7948 2372
rect 7988 2332 7989 2372
rect 7947 2323 7989 2332
rect 7947 2036 7989 2045
rect 7468 1996 7796 2036
rect 7276 1912 7412 1952
rect 7179 1903 7221 1912
rect 7180 80 7220 1903
rect 7372 80 7412 1912
rect 7563 1700 7605 1709
rect 7563 1660 7564 1700
rect 7604 1660 7605 1700
rect 7563 1651 7605 1660
rect 7564 80 7604 1651
rect 7756 80 7796 1996
rect 7947 1996 7948 2036
rect 7988 1996 7989 2036
rect 8044 2036 8084 3928
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8140 3330 8180 3415
rect 8236 2372 8276 3928
rect 8620 3968 8660 3977
rect 8524 3464 8564 3473
rect 8428 3424 8524 3464
rect 8332 3212 8372 3221
rect 8332 2633 8372 3172
rect 8428 3053 8468 3424
rect 8524 3415 8564 3424
rect 8523 3212 8565 3221
rect 8523 3172 8524 3212
rect 8564 3172 8565 3212
rect 8523 3163 8565 3172
rect 8427 3044 8469 3053
rect 8427 3004 8428 3044
rect 8468 3004 8469 3044
rect 8427 2995 8469 3004
rect 8331 2624 8373 2633
rect 8331 2584 8332 2624
rect 8372 2584 8373 2624
rect 8331 2575 8373 2584
rect 8236 2332 8468 2372
rect 8331 2204 8373 2213
rect 8331 2164 8332 2204
rect 8372 2164 8373 2204
rect 8331 2155 8373 2164
rect 8044 1996 8180 2036
rect 7947 1987 7989 1996
rect 7948 80 7988 1987
rect 8140 80 8180 1996
rect 8332 80 8372 2155
rect 8428 1532 8468 2332
rect 8524 1616 8564 3163
rect 8620 2036 8660 3928
rect 8908 3464 8948 5263
rect 9196 5237 9236 9379
rect 9579 9344 9621 9353
rect 9579 9304 9580 9344
rect 9620 9304 9621 9344
rect 9579 9295 9621 9304
rect 9483 8336 9525 8345
rect 9483 8296 9484 8336
rect 9524 8296 9525 8336
rect 9483 8287 9525 8296
rect 9291 8168 9333 8177
rect 9291 8128 9292 8168
rect 9332 8128 9333 8168
rect 9291 8119 9333 8128
rect 9292 7925 9332 8119
rect 9291 7916 9333 7925
rect 9291 7876 9292 7916
rect 9332 7876 9333 7916
rect 9291 7867 9333 7876
rect 9484 7916 9524 8287
rect 9484 7867 9524 7876
rect 9292 7782 9332 7867
rect 9388 7832 9428 7841
rect 9195 5228 9237 5237
rect 9195 5188 9196 5228
rect 9236 5188 9237 5228
rect 9195 5179 9237 5188
rect 9291 5144 9333 5153
rect 9291 5104 9292 5144
rect 9332 5104 9333 5144
rect 9291 5095 9333 5104
rect 9195 4724 9237 4733
rect 9195 4684 9196 4724
rect 9236 4684 9237 4724
rect 9195 4675 9237 4684
rect 9196 4136 9236 4675
rect 9196 4087 9236 4096
rect 9004 3968 9044 3977
rect 9044 3928 9236 3968
rect 9004 3919 9044 3928
rect 8908 3415 8948 3424
rect 8716 3212 8756 3221
rect 8716 2213 8756 3172
rect 9100 3212 9140 3221
rect 9196 3212 9236 3928
rect 9292 3464 9332 5095
rect 9388 4649 9428 7792
rect 9580 7748 9620 9295
rect 9771 9260 9813 9269
rect 9771 9220 9772 9260
rect 9812 9220 9813 9260
rect 9771 9211 9813 9220
rect 9772 8840 9812 9211
rect 9772 8791 9812 8800
rect 9675 8756 9717 8765
rect 9675 8716 9676 8756
rect 9716 8716 9717 8756
rect 9675 8707 9717 8716
rect 9868 8756 9908 8765
rect 10059 8756 10101 8765
rect 9908 8716 10004 8756
rect 9868 8707 9908 8716
rect 9676 8622 9716 8707
rect 9867 8000 9909 8009
rect 9867 7960 9868 8000
rect 9908 7960 9909 8000
rect 9867 7951 9909 7960
rect 9675 7916 9717 7925
rect 9675 7876 9676 7916
rect 9716 7876 9717 7916
rect 9675 7867 9717 7876
rect 9868 7916 9908 7951
rect 9676 7782 9716 7867
rect 9868 7865 9908 7876
rect 9772 7832 9812 7841
rect 9484 7708 9620 7748
rect 9484 7085 9524 7708
rect 9772 7412 9812 7792
rect 9580 7372 9812 7412
rect 9964 7412 10004 8716
rect 10059 8716 10060 8756
rect 10100 8716 10101 8756
rect 10059 8707 10101 8716
rect 10252 8756 10292 8765
rect 10635 8756 10677 8765
rect 10292 8716 10484 8756
rect 10252 8707 10292 8716
rect 10060 8177 10100 8707
rect 10156 8504 10196 8513
rect 10196 8464 10388 8504
rect 10156 8455 10196 8464
rect 10155 8336 10197 8345
rect 10155 8296 10156 8336
rect 10196 8296 10197 8336
rect 10155 8287 10197 8296
rect 10059 8168 10101 8177
rect 10059 8128 10060 8168
rect 10100 8128 10101 8168
rect 10059 8119 10101 8128
rect 10156 8000 10196 8287
rect 10060 7960 10196 8000
rect 10251 8000 10293 8009
rect 10251 7960 10252 8000
rect 10292 7960 10293 8000
rect 10060 7916 10100 7960
rect 10251 7951 10293 7960
rect 10060 7867 10100 7876
rect 10252 7916 10292 7951
rect 10156 7832 10196 7841
rect 10059 7412 10101 7421
rect 9964 7372 10060 7412
rect 10100 7372 10101 7412
rect 9483 7076 9525 7085
rect 9483 7036 9484 7076
rect 9524 7036 9525 7076
rect 9483 7027 9525 7036
rect 9580 5657 9620 7372
rect 10059 7363 10101 7372
rect 9675 7244 9717 7253
rect 9675 7204 9676 7244
rect 9716 7204 9717 7244
rect 9675 7195 9717 7204
rect 9867 7244 9909 7253
rect 9867 7204 9868 7244
rect 9908 7204 9909 7244
rect 9867 7195 9909 7204
rect 10060 7244 10100 7363
rect 10156 7337 10196 7792
rect 10155 7328 10197 7337
rect 10155 7288 10156 7328
rect 10196 7288 10197 7328
rect 10155 7279 10197 7288
rect 10060 7195 10100 7204
rect 10252 7244 10292 7876
rect 10348 7673 10388 8464
rect 10444 7916 10484 8716
rect 10635 8716 10636 8756
rect 10676 8716 10677 8756
rect 10635 8707 10677 8716
rect 10636 8009 10676 8707
rect 10635 8000 10677 8009
rect 10635 7960 10636 8000
rect 10676 7960 10677 8000
rect 10635 7951 10677 7960
rect 10347 7664 10389 7673
rect 10347 7624 10348 7664
rect 10388 7624 10389 7664
rect 10347 7615 10389 7624
rect 10444 7589 10484 7876
rect 10636 7916 10676 7951
rect 10636 7866 10676 7876
rect 10540 7832 10580 7841
rect 10443 7580 10485 7589
rect 10443 7540 10444 7580
rect 10484 7540 10485 7580
rect 10443 7531 10485 7540
rect 10540 7412 10580 7792
rect 10635 7580 10677 7589
rect 10635 7540 10636 7580
rect 10676 7540 10677 7580
rect 10635 7531 10677 7540
rect 10444 7372 10580 7412
rect 10347 7328 10389 7337
rect 10347 7288 10348 7328
rect 10388 7288 10389 7328
rect 10347 7279 10389 7288
rect 10252 7195 10292 7204
rect 9676 7110 9716 7195
rect 9868 7110 9908 7195
rect 9963 7076 10005 7085
rect 9963 7036 9964 7076
rect 10004 7036 10005 7076
rect 9963 7027 10005 7036
rect 9771 6992 9813 7001
rect 9771 6952 9772 6992
rect 9812 6952 9813 6992
rect 9771 6943 9813 6952
rect 9772 6858 9812 6943
rect 9675 5900 9717 5909
rect 9675 5860 9676 5900
rect 9716 5860 9717 5900
rect 9675 5851 9717 5860
rect 9579 5648 9621 5657
rect 9579 5608 9580 5648
rect 9620 5608 9621 5648
rect 9579 5599 9621 5608
rect 9579 5228 9621 5237
rect 9579 5188 9580 5228
rect 9620 5188 9621 5228
rect 9579 5179 9621 5188
rect 9387 4640 9429 4649
rect 9387 4600 9388 4640
rect 9428 4600 9429 4640
rect 9387 4591 9429 4600
rect 9580 4136 9620 5179
rect 9580 4087 9620 4096
rect 9292 3415 9332 3424
rect 9388 3968 9428 3977
rect 9196 3172 9332 3212
rect 9100 2540 9140 3172
rect 9100 2500 9236 2540
rect 9099 2372 9141 2381
rect 9099 2332 9100 2372
rect 9140 2332 9141 2372
rect 9099 2323 9141 2332
rect 8715 2204 8757 2213
rect 8715 2164 8716 2204
rect 8756 2164 8757 2204
rect 8715 2155 8757 2164
rect 8620 1996 8948 2036
rect 8524 1576 8756 1616
rect 8428 1492 8564 1532
rect 8524 80 8564 1492
rect 8716 80 8756 1576
rect 8908 80 8948 1996
rect 9100 80 9140 2323
rect 9196 1373 9236 2500
rect 9195 1364 9237 1373
rect 9195 1324 9196 1364
rect 9236 1324 9237 1364
rect 9195 1315 9237 1324
rect 9292 80 9332 3172
rect 9388 1037 9428 3928
rect 9676 3464 9716 5851
rect 9964 4136 10004 7027
rect 10156 6992 10196 7001
rect 10059 6740 10101 6749
rect 10059 6700 10060 6740
rect 10100 6700 10101 6740
rect 10059 6691 10101 6700
rect 10060 4136 10100 6691
rect 10156 6497 10196 6952
rect 10251 6572 10293 6581
rect 10251 6532 10252 6572
rect 10292 6532 10293 6572
rect 10251 6523 10293 6532
rect 10155 6488 10197 6497
rect 10155 6448 10156 6488
rect 10196 6448 10197 6488
rect 10155 6439 10197 6448
rect 10252 4901 10292 6523
rect 10251 4892 10293 4901
rect 10251 4852 10252 4892
rect 10292 4852 10293 4892
rect 10251 4843 10293 4852
rect 10348 4817 10388 7279
rect 10444 6581 10484 7372
rect 10539 7244 10581 7253
rect 10539 7204 10540 7244
rect 10580 7204 10581 7244
rect 10539 7195 10581 7204
rect 10636 7244 10676 7531
rect 10636 7195 10676 7204
rect 10540 6992 10580 7195
rect 10732 7160 10772 10807
rect 11788 10781 11828 10900
rect 11980 10940 12020 10975
rect 10827 10772 10869 10781
rect 10827 10732 10828 10772
rect 10868 10732 10869 10772
rect 10827 10723 10869 10732
rect 11499 10772 11541 10781
rect 11499 10732 11500 10772
rect 11540 10732 11541 10772
rect 11499 10723 11541 10732
rect 11787 10772 11829 10781
rect 11787 10732 11788 10772
rect 11828 10732 11829 10772
rect 11787 10723 11829 10732
rect 10828 10268 10868 10723
rect 10923 10604 10965 10613
rect 10923 10564 10924 10604
rect 10964 10564 10965 10604
rect 10923 10555 10965 10564
rect 10924 10352 10964 10555
rect 11211 10520 11253 10529
rect 11211 10480 11212 10520
rect 11252 10480 11253 10520
rect 11211 10471 11253 10480
rect 10924 10303 10964 10312
rect 10828 10219 10868 10228
rect 11020 10268 11060 10277
rect 11212 10268 11252 10471
rect 11060 10228 11212 10268
rect 11020 10219 11060 10228
rect 11212 10219 11252 10228
rect 11403 10268 11445 10277
rect 11403 10228 11404 10268
rect 11444 10228 11445 10268
rect 11403 10219 11445 10228
rect 11404 10134 11444 10219
rect 11308 10016 11348 10025
rect 11308 8933 11348 9976
rect 11403 9596 11445 9605
rect 11403 9556 11404 9596
rect 11444 9556 11445 9596
rect 11403 9547 11445 9556
rect 11307 8924 11349 8933
rect 11307 8884 11308 8924
rect 11348 8884 11349 8924
rect 11307 8875 11349 8884
rect 11115 8756 11157 8765
rect 11115 8716 11116 8756
rect 11156 8716 11157 8756
rect 11115 8707 11157 8716
rect 11308 8756 11348 8765
rect 11116 8622 11156 8707
rect 11308 8597 11348 8716
rect 11307 8588 11349 8597
rect 11307 8548 11308 8588
rect 11348 8548 11349 8588
rect 11307 8539 11349 8548
rect 11212 8504 11252 8513
rect 11019 8420 11061 8429
rect 11019 8380 11020 8420
rect 11060 8380 11061 8420
rect 11019 8371 11061 8380
rect 10923 8336 10965 8345
rect 10923 8296 10924 8336
rect 10964 8296 10965 8336
rect 10923 8287 10965 8296
rect 10828 7337 10868 7352
rect 10827 7328 10869 7337
rect 10827 7288 10828 7328
rect 10868 7288 10869 7328
rect 10827 7279 10869 7288
rect 10828 7257 10868 7279
rect 10828 7208 10868 7217
rect 10732 7120 10868 7160
rect 10732 6992 10772 7001
rect 10540 6952 10676 6992
rect 10443 6572 10485 6581
rect 10443 6532 10444 6572
rect 10484 6532 10485 6572
rect 10443 6523 10485 6532
rect 10443 6404 10485 6413
rect 10443 6364 10444 6404
rect 10484 6364 10485 6404
rect 10443 6355 10485 6364
rect 10636 6404 10676 6952
rect 10636 6355 10676 6364
rect 10444 6270 10484 6355
rect 10540 6320 10580 6329
rect 10347 4808 10389 4817
rect 10347 4768 10348 4808
rect 10388 4768 10389 4808
rect 10347 4759 10389 4768
rect 10540 4145 10580 6280
rect 10732 4313 10772 6952
rect 10731 4304 10773 4313
rect 10731 4264 10732 4304
rect 10772 4264 10773 4304
rect 10731 4255 10773 4264
rect 10348 4136 10388 4145
rect 10060 4096 10348 4136
rect 9964 4087 10004 4096
rect 10348 4087 10388 4096
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10732 4136 10772 4145
rect 10828 4136 10868 7120
rect 10924 6413 10964 8287
rect 11020 7925 11060 8371
rect 11019 7916 11061 7925
rect 11019 7876 11020 7916
rect 11060 7876 11061 7916
rect 11019 7867 11061 7876
rect 11020 7244 11060 7867
rect 11212 7412 11252 8464
rect 11212 7372 11348 7412
rect 11020 7195 11060 7204
rect 11211 7244 11253 7253
rect 11211 7204 11212 7244
rect 11252 7204 11253 7244
rect 11211 7195 11253 7204
rect 11212 7001 11252 7195
rect 11116 6992 11156 7001
rect 10923 6404 10965 6413
rect 10923 6364 10924 6404
rect 10964 6364 10965 6404
rect 10923 6355 10965 6364
rect 11116 6329 11156 6952
rect 11211 6992 11253 7001
rect 11211 6952 11212 6992
rect 11252 6952 11253 6992
rect 11211 6943 11253 6952
rect 11115 6320 11157 6329
rect 11115 6280 11116 6320
rect 11156 6280 11157 6320
rect 11115 6271 11157 6280
rect 11308 5648 11348 7372
rect 11404 6488 11444 9547
rect 11500 9428 11540 10723
rect 11595 10688 11637 10697
rect 11595 10648 11596 10688
rect 11636 10648 11637 10688
rect 11595 10639 11637 10648
rect 11596 10277 11636 10639
rect 11595 10268 11637 10277
rect 11595 10228 11596 10268
rect 11636 10228 11637 10268
rect 11595 10219 11637 10228
rect 11788 10268 11828 10277
rect 11980 10268 12020 10900
rect 12171 10940 12213 10949
rect 12171 10900 12172 10940
rect 12212 10900 12213 10940
rect 12171 10891 12213 10900
rect 12364 10940 12404 10949
rect 12172 10806 12212 10891
rect 12268 10856 12308 10865
rect 12268 10604 12308 10816
rect 12364 10697 12404 10900
rect 12363 10688 12405 10697
rect 12363 10648 12364 10688
rect 12404 10648 12405 10688
rect 12363 10639 12405 10648
rect 12076 10564 12308 10604
rect 12076 10277 12116 10564
rect 12363 10520 12405 10529
rect 12363 10480 12364 10520
rect 12404 10480 12405 10520
rect 12363 10471 12405 10480
rect 12171 10436 12213 10445
rect 12171 10396 12172 10436
rect 12212 10396 12213 10436
rect 12171 10387 12213 10396
rect 11828 10228 11980 10268
rect 11788 10219 11828 10228
rect 11980 10219 12020 10228
rect 12075 10268 12117 10277
rect 12075 10228 12076 10268
rect 12116 10228 12117 10268
rect 12075 10219 12117 10228
rect 12172 10268 12212 10387
rect 12364 10289 12404 10471
rect 12212 10228 12308 10268
rect 12364 10240 12404 10249
rect 12172 10219 12212 10228
rect 11596 10134 11636 10219
rect 11787 10100 11829 10109
rect 11787 10060 11788 10100
rect 11828 10060 11829 10100
rect 11787 10051 11829 10060
rect 11692 10016 11732 10025
rect 11692 9605 11732 9976
rect 11691 9596 11733 9605
rect 11691 9556 11692 9596
rect 11732 9556 11733 9596
rect 11691 9547 11733 9556
rect 11596 9428 11636 9437
rect 11500 9388 11596 9428
rect 11596 9379 11636 9388
rect 11788 9428 11828 10051
rect 12076 10016 12116 10025
rect 12116 9976 12212 10016
rect 12076 9967 12116 9976
rect 12076 9428 12116 9437
rect 11788 9379 11828 9388
rect 11884 9388 12076 9428
rect 11692 9344 11732 9353
rect 11692 9185 11732 9304
rect 11691 9176 11733 9185
rect 11691 9136 11692 9176
rect 11732 9136 11733 9176
rect 11691 9127 11733 9136
rect 11787 8924 11829 8933
rect 11787 8884 11788 8924
rect 11828 8884 11829 8924
rect 11787 8875 11829 8884
rect 11500 8765 11540 8850
rect 11595 8840 11637 8849
rect 11595 8800 11596 8840
rect 11636 8800 11637 8840
rect 11595 8791 11637 8800
rect 11499 8756 11541 8765
rect 11499 8716 11500 8756
rect 11540 8716 11541 8756
rect 11499 8707 11541 8716
rect 11596 8706 11636 8791
rect 11692 8756 11732 8765
rect 11692 8168 11732 8716
rect 11788 8504 11828 8875
rect 11884 8765 11924 9388
rect 12076 9379 12116 9388
rect 11979 9008 12021 9017
rect 11979 8968 11980 9008
rect 12020 8968 12021 9008
rect 11979 8959 12021 8968
rect 11980 8840 12020 8959
rect 11980 8791 12020 8800
rect 11883 8756 11925 8765
rect 11883 8716 11884 8756
rect 11924 8716 11925 8756
rect 11883 8707 11925 8716
rect 12076 8756 12116 8765
rect 11884 8622 11924 8707
rect 11788 8464 11924 8504
rect 11596 8128 11732 8168
rect 11596 7916 11636 8128
rect 11596 7757 11636 7876
rect 11788 7916 11828 7925
rect 11691 7832 11733 7841
rect 11691 7792 11692 7832
rect 11732 7792 11733 7832
rect 11691 7783 11733 7792
rect 11595 7748 11637 7757
rect 11595 7708 11596 7748
rect 11636 7708 11637 7748
rect 11595 7699 11637 7708
rect 11692 7698 11732 7783
rect 11691 7496 11733 7505
rect 11691 7456 11692 7496
rect 11732 7456 11733 7496
rect 11691 7447 11733 7456
rect 11404 6448 11540 6488
rect 11020 5608 11348 5648
rect 11020 4229 11060 5608
rect 11211 5060 11253 5069
rect 11211 5020 11212 5060
rect 11252 5020 11253 5060
rect 11211 5011 11253 5020
rect 11019 4220 11061 4229
rect 11019 4180 11020 4220
rect 11060 4180 11061 4220
rect 11019 4171 11061 4180
rect 11116 4145 11156 4230
rect 10772 4096 10868 4136
rect 11115 4136 11157 4145
rect 11115 4096 11116 4136
rect 11156 4096 11157 4136
rect 10732 4087 10772 4096
rect 11115 4087 11157 4096
rect 9676 3415 9716 3424
rect 9772 3968 9812 3977
rect 9484 3212 9524 3221
rect 9524 3172 9620 3212
rect 9484 3163 9524 3172
rect 9483 2540 9525 2549
rect 9483 2500 9484 2540
rect 9524 2500 9525 2540
rect 9483 2491 9525 2500
rect 9387 1028 9429 1037
rect 9387 988 9388 1028
rect 9428 988 9429 1028
rect 9387 979 9429 988
rect 9484 80 9524 2491
rect 9580 1625 9620 3172
rect 9675 2204 9717 2213
rect 9675 2164 9676 2204
rect 9716 2164 9717 2204
rect 9675 2155 9717 2164
rect 9579 1616 9621 1625
rect 9579 1576 9580 1616
rect 9620 1576 9621 1616
rect 9579 1567 9621 1576
rect 9676 1196 9716 2155
rect 9772 1280 9812 3928
rect 10156 3968 10196 3977
rect 10540 3968 10580 3977
rect 10924 3968 10964 3977
rect 10196 3928 10388 3968
rect 10156 3919 10196 3928
rect 10059 3464 10101 3473
rect 10059 3424 10060 3464
rect 10100 3424 10101 3464
rect 10059 3415 10101 3424
rect 10060 3330 10100 3415
rect 9868 3212 9908 3221
rect 9868 1709 9908 3172
rect 10252 3212 10292 3221
rect 9867 1700 9909 1709
rect 9867 1660 9868 1700
rect 9908 1660 9909 1700
rect 9867 1651 9909 1660
rect 10252 1541 10292 3172
rect 10348 2036 10388 3928
rect 10580 3928 10772 3968
rect 10540 3919 10580 3928
rect 10444 3464 10484 3473
rect 10444 3137 10484 3424
rect 10636 3212 10676 3221
rect 10443 3128 10485 3137
rect 10443 3088 10444 3128
rect 10484 3088 10485 3128
rect 10443 3079 10485 3088
rect 10348 1996 10484 2036
rect 10251 1532 10293 1541
rect 10251 1492 10252 1532
rect 10292 1492 10293 1532
rect 10251 1483 10293 1492
rect 10251 1364 10293 1373
rect 10251 1324 10252 1364
rect 10292 1324 10293 1364
rect 10251 1315 10293 1324
rect 9772 1240 10100 1280
rect 9676 1156 9908 1196
rect 9675 1028 9717 1037
rect 9675 988 9676 1028
rect 9716 988 9717 1028
rect 9675 979 9717 988
rect 9676 80 9716 979
rect 9868 80 9908 1156
rect 10060 80 10100 1240
rect 10252 80 10292 1315
rect 10444 80 10484 1996
rect 10636 1793 10676 3172
rect 10732 2036 10772 3928
rect 10964 3928 11156 3968
rect 10924 3919 10964 3928
rect 10828 3464 10868 3473
rect 10828 3305 10868 3424
rect 10827 3296 10869 3305
rect 10827 3256 10828 3296
rect 10868 3256 10869 3296
rect 10827 3247 10869 3256
rect 11020 3212 11060 3221
rect 10732 1996 10868 2036
rect 10635 1784 10677 1793
rect 10635 1744 10636 1784
rect 10676 1744 10677 1784
rect 10635 1735 10677 1744
rect 10635 1616 10677 1625
rect 10635 1576 10636 1616
rect 10676 1576 10677 1616
rect 10635 1567 10677 1576
rect 10636 80 10676 1567
rect 10828 80 10868 1996
rect 11020 1877 11060 3172
rect 11116 2036 11156 3928
rect 11212 3464 11252 5011
rect 11500 4136 11540 6448
rect 11595 5228 11637 5237
rect 11595 5188 11596 5228
rect 11636 5188 11637 5228
rect 11595 5179 11637 5188
rect 11500 4087 11540 4096
rect 11308 3968 11348 3977
rect 11348 3928 11540 3968
rect 11308 3919 11348 3928
rect 11212 3415 11252 3424
rect 11404 3212 11444 3221
rect 11116 1996 11252 2036
rect 11019 1868 11061 1877
rect 11019 1828 11020 1868
rect 11060 1828 11061 1868
rect 11019 1819 11061 1828
rect 11019 1700 11061 1709
rect 11019 1660 11020 1700
rect 11060 1660 11061 1700
rect 11019 1651 11061 1660
rect 11020 80 11060 1651
rect 11212 80 11252 1996
rect 11404 1709 11444 3172
rect 11500 2540 11540 3928
rect 11596 3464 11636 5179
rect 11692 4136 11732 7447
rect 11788 7001 11828 7876
rect 11884 7505 11924 8464
rect 11979 8168 12021 8177
rect 11979 8128 11980 8168
rect 12020 8128 12021 8168
rect 11979 8119 12021 8128
rect 11980 7916 12020 8119
rect 12076 8009 12116 8716
rect 12172 8084 12212 9976
rect 12268 9428 12308 10228
rect 12460 10184 12500 11152
rect 12747 10940 12789 10949
rect 15628 10940 15668 10949
rect 12747 10900 12748 10940
rect 12788 10900 12789 10940
rect 12747 10891 12789 10900
rect 15532 10900 15628 10940
rect 12555 10436 12597 10445
rect 12555 10396 12556 10436
rect 12596 10396 12597 10436
rect 12555 10387 12597 10396
rect 12556 10268 12596 10387
rect 12556 10219 12596 10228
rect 12748 10268 12788 10891
rect 14571 10772 14613 10781
rect 14571 10732 14572 10772
rect 14612 10732 14613 10772
rect 14571 10723 14613 10732
rect 15147 10772 15189 10781
rect 15147 10732 15148 10772
rect 15188 10732 15189 10772
rect 15147 10723 15189 10732
rect 14475 10604 14517 10613
rect 14475 10564 14476 10604
rect 14516 10564 14517 10604
rect 14475 10555 14517 10564
rect 12939 10436 12981 10445
rect 12939 10396 12940 10436
rect 12980 10396 12981 10436
rect 12939 10387 12981 10396
rect 12268 9379 12308 9388
rect 12364 10144 12500 10184
rect 12364 9260 12404 10144
rect 12748 10109 12788 10228
rect 12940 10268 12980 10387
rect 12940 10219 12980 10228
rect 14476 10193 14516 10555
rect 14572 10277 14612 10723
rect 14955 10688 14997 10697
rect 14955 10648 14956 10688
rect 14996 10648 14997 10688
rect 14955 10639 14997 10648
rect 14763 10604 14805 10613
rect 14763 10564 14764 10604
rect 14804 10564 14805 10604
rect 14763 10555 14805 10564
rect 14571 10268 14613 10277
rect 14571 10228 14572 10268
rect 14612 10228 14613 10268
rect 14571 10219 14613 10228
rect 14764 10268 14804 10555
rect 12843 10184 12885 10193
rect 12843 10144 12844 10184
rect 12884 10144 12885 10184
rect 12843 10135 12885 10144
rect 14475 10184 14517 10193
rect 14475 10144 14476 10184
rect 14516 10144 14517 10184
rect 14475 10135 14517 10144
rect 12747 10100 12789 10109
rect 12747 10060 12748 10100
rect 12788 10060 12789 10100
rect 12747 10051 12789 10060
rect 12844 10050 12884 10135
rect 14572 10134 14612 10219
rect 12460 10016 12500 10025
rect 14668 10016 14708 10025
rect 12500 9976 12596 10016
rect 12460 9967 12500 9976
rect 12364 9220 12500 9260
rect 12363 9092 12405 9101
rect 12363 9052 12364 9092
rect 12404 9052 12405 9092
rect 12363 9043 12405 9052
rect 12364 8840 12404 9043
rect 12460 8933 12500 9220
rect 12459 8924 12501 8933
rect 12459 8884 12460 8924
rect 12500 8884 12501 8924
rect 12459 8875 12501 8884
rect 12556 8849 12596 9976
rect 13996 9976 14668 10016
rect 13035 9260 13077 9269
rect 13035 9220 13036 9260
rect 13076 9220 13077 9260
rect 13035 9211 13077 9220
rect 12364 8791 12404 8800
rect 12555 8840 12597 8849
rect 12555 8800 12556 8840
rect 12596 8800 12597 8840
rect 12555 8791 12597 8800
rect 12267 8756 12309 8765
rect 12267 8716 12268 8756
rect 12308 8716 12309 8756
rect 12267 8707 12309 8716
rect 12459 8756 12501 8765
rect 12459 8716 12460 8756
rect 12500 8716 12501 8756
rect 12459 8707 12501 8716
rect 12651 8756 12693 8765
rect 12651 8716 12652 8756
rect 12692 8716 12693 8756
rect 12651 8707 12693 8716
rect 12268 8622 12308 8707
rect 12460 8622 12500 8707
rect 12459 8084 12501 8093
rect 12172 8044 12308 8084
rect 12075 8000 12117 8009
rect 12075 7960 12076 8000
rect 12116 7960 12117 8000
rect 12075 7951 12117 7960
rect 11980 7867 12020 7876
rect 12172 7916 12212 7925
rect 12075 7832 12117 7841
rect 12075 7792 12076 7832
rect 12116 7792 12117 7832
rect 12075 7783 12117 7792
rect 12076 7698 12116 7783
rect 12172 7757 12212 7876
rect 12171 7748 12213 7757
rect 12171 7708 12172 7748
rect 12212 7708 12213 7748
rect 12171 7699 12213 7708
rect 11883 7496 11925 7505
rect 11883 7456 11884 7496
rect 11924 7456 11925 7496
rect 11883 7447 11925 7456
rect 11883 7328 11925 7337
rect 11883 7288 11884 7328
rect 11924 7288 11925 7328
rect 11883 7279 11925 7288
rect 11884 7244 11924 7279
rect 11884 7193 11924 7204
rect 12076 7244 12116 7253
rect 11980 7076 12020 7085
rect 11787 6992 11829 7001
rect 11787 6952 11788 6992
rect 11828 6952 11829 6992
rect 11787 6943 11829 6952
rect 11980 4985 12020 7036
rect 12076 7001 12116 7204
rect 12268 7169 12308 8044
rect 12459 8044 12460 8084
rect 12500 8044 12501 8084
rect 12459 8035 12501 8044
rect 12460 7950 12500 8035
rect 12363 7916 12405 7925
rect 12363 7876 12364 7916
rect 12404 7876 12405 7916
rect 12363 7867 12405 7876
rect 12556 7916 12596 7925
rect 12364 7782 12404 7867
rect 12556 7832 12596 7876
rect 12553 7792 12596 7832
rect 12553 7664 12593 7792
rect 12553 7624 12596 7664
rect 12556 7505 12596 7624
rect 12555 7496 12597 7505
rect 12555 7456 12556 7496
rect 12596 7456 12597 7496
rect 12555 7447 12597 7456
rect 12652 7328 12692 8707
rect 12939 8252 12981 8261
rect 12939 8212 12940 8252
rect 12980 8212 12981 8252
rect 12939 8203 12981 8212
rect 12747 8168 12789 8177
rect 12747 8128 12748 8168
rect 12788 8128 12789 8168
rect 12747 8119 12789 8128
rect 12748 7916 12788 8119
rect 12940 7925 12980 8203
rect 12748 7867 12788 7876
rect 12939 7916 12981 7925
rect 12939 7876 12940 7916
rect 12980 7876 12981 7916
rect 12939 7867 12981 7876
rect 12844 7832 12884 7841
rect 12747 7496 12789 7505
rect 12747 7456 12748 7496
rect 12788 7456 12789 7496
rect 12747 7447 12789 7456
rect 12556 7288 12692 7328
rect 12556 7244 12596 7288
rect 12556 7195 12596 7204
rect 12748 7244 12788 7447
rect 12267 7160 12309 7169
rect 12267 7120 12268 7160
rect 12308 7120 12309 7160
rect 12267 7111 12309 7120
rect 12748 7001 12788 7204
rect 12844 7169 12884 7792
rect 12940 7782 12980 7867
rect 13036 7664 13076 9211
rect 13323 8756 13365 8765
rect 13323 8716 13324 8756
rect 13364 8716 13365 8756
rect 13323 8707 13365 8716
rect 13131 8168 13173 8177
rect 13131 8128 13132 8168
rect 13172 8128 13173 8168
rect 13131 8119 13173 8128
rect 13132 7916 13172 8119
rect 13324 8093 13364 8707
rect 13707 8672 13749 8681
rect 13707 8632 13708 8672
rect 13748 8632 13749 8672
rect 13707 8623 13749 8632
rect 13515 8168 13557 8177
rect 13515 8128 13516 8168
rect 13556 8128 13557 8168
rect 13515 8119 13557 8128
rect 13323 8084 13365 8093
rect 13323 8044 13324 8084
rect 13364 8044 13365 8084
rect 13323 8035 13365 8044
rect 13132 7867 13172 7876
rect 13324 7916 13364 8035
rect 13324 7867 13364 7876
rect 13516 7916 13556 8119
rect 13516 7867 13556 7876
rect 13708 7916 13748 8623
rect 12940 7624 13076 7664
rect 13228 7832 13268 7841
rect 12843 7160 12885 7169
rect 12843 7120 12844 7160
rect 12884 7120 12885 7160
rect 12843 7111 12885 7120
rect 12075 6992 12117 7001
rect 12075 6952 12076 6992
rect 12116 6952 12117 6992
rect 12075 6943 12117 6952
rect 12652 6992 12692 7001
rect 12267 6572 12309 6581
rect 12267 6532 12268 6572
rect 12308 6532 12309 6572
rect 12267 6523 12309 6532
rect 11979 4976 12021 4985
rect 11979 4936 11980 4976
rect 12020 4936 12021 4976
rect 11979 4927 12021 4936
rect 11884 4136 11924 4145
rect 11692 4096 11884 4136
rect 11884 4087 11924 4096
rect 12268 4136 12308 6523
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12556 6245 12596 6439
rect 12555 6236 12597 6245
rect 12555 6196 12556 6236
rect 12596 6196 12597 6236
rect 12555 6187 12597 6196
rect 12652 4733 12692 6952
rect 12747 6992 12789 7001
rect 12747 6952 12748 6992
rect 12788 6952 12789 6992
rect 12747 6943 12789 6952
rect 12651 4724 12693 4733
rect 12651 4684 12652 4724
rect 12692 4684 12693 4724
rect 12651 4675 12693 4684
rect 12363 4640 12405 4649
rect 12363 4600 12364 4640
rect 12404 4600 12405 4640
rect 12363 4591 12405 4600
rect 12268 4087 12308 4096
rect 11692 3968 11732 3977
rect 12076 3968 12116 3977
rect 11732 3928 11924 3968
rect 11692 3919 11732 3928
rect 11596 3415 11636 3424
rect 11788 3212 11828 3221
rect 11500 2500 11636 2540
rect 11403 1700 11445 1709
rect 11403 1660 11404 1700
rect 11444 1660 11445 1700
rect 11403 1651 11445 1660
rect 11403 1532 11445 1541
rect 11403 1492 11404 1532
rect 11444 1492 11445 1532
rect 11403 1483 11445 1492
rect 11404 80 11444 1483
rect 11596 80 11636 2500
rect 11788 1961 11828 3172
rect 11884 2540 11924 3928
rect 12116 3928 12308 3968
rect 12076 3919 12116 3928
rect 11979 3632 12021 3641
rect 11979 3592 11980 3632
rect 12020 3592 12021 3632
rect 11979 3583 12021 3592
rect 11980 3464 12020 3583
rect 11980 3415 12020 3424
rect 12172 3212 12212 3221
rect 11884 2500 12020 2540
rect 11787 1952 11829 1961
rect 11787 1912 11788 1952
rect 11828 1912 11829 1952
rect 11787 1903 11829 1912
rect 11787 1784 11829 1793
rect 11787 1744 11788 1784
rect 11828 1744 11829 1784
rect 11787 1735 11829 1744
rect 11788 80 11828 1735
rect 11980 80 12020 2500
rect 12172 2297 12212 3172
rect 12268 2540 12308 3928
rect 12364 3464 12404 4591
rect 12652 4136 12692 4145
rect 12940 4136 12980 7624
rect 13131 7160 13173 7169
rect 13131 7120 13132 7160
rect 13172 7120 13173 7160
rect 13131 7111 13173 7120
rect 13035 4472 13077 4481
rect 13035 4432 13036 4472
rect 13076 4432 13077 4472
rect 13035 4423 13077 4432
rect 12692 4096 12980 4136
rect 13036 4136 13076 4423
rect 12652 4087 12692 4096
rect 13036 4087 13076 4096
rect 12460 3968 12500 3977
rect 12844 3968 12884 3977
rect 12500 3928 12692 3968
rect 12460 3919 12500 3928
rect 12364 3415 12404 3424
rect 12556 3212 12596 3221
rect 12556 2540 12596 3172
rect 12268 2500 12404 2540
rect 12171 2288 12213 2297
rect 12171 2248 12172 2288
rect 12212 2248 12213 2288
rect 12171 2239 12213 2248
rect 12171 1868 12213 1877
rect 12171 1828 12172 1868
rect 12212 1828 12213 1868
rect 12171 1819 12213 1828
rect 12172 80 12212 1819
rect 12364 80 12404 2500
rect 12460 2500 12596 2540
rect 12460 533 12500 2500
rect 12555 1700 12597 1709
rect 12555 1660 12556 1700
rect 12596 1660 12597 1700
rect 12555 1651 12597 1660
rect 12459 524 12501 533
rect 12459 484 12460 524
rect 12500 484 12501 524
rect 12459 475 12501 484
rect 12556 80 12596 1651
rect 12652 1280 12692 3928
rect 12748 3464 12788 3473
rect 12748 1709 12788 3424
rect 12747 1700 12789 1709
rect 12747 1660 12748 1700
rect 12788 1660 12789 1700
rect 12747 1651 12789 1660
rect 12652 1240 12788 1280
rect 12748 80 12788 1240
rect 12844 617 12884 3928
rect 13132 3464 13172 7111
rect 13228 6413 13268 7792
rect 13612 7832 13652 7841
rect 13323 7664 13365 7673
rect 13323 7624 13324 7664
rect 13364 7624 13365 7664
rect 13323 7615 13365 7624
rect 13227 6404 13269 6413
rect 13227 6364 13228 6404
rect 13268 6364 13269 6404
rect 13227 6355 13269 6364
rect 13324 4136 13364 7615
rect 13612 7421 13652 7792
rect 13708 7673 13748 7876
rect 13707 7664 13749 7673
rect 13707 7624 13708 7664
rect 13748 7624 13749 7664
rect 13707 7615 13749 7624
rect 13611 7412 13653 7421
rect 13611 7372 13612 7412
rect 13652 7372 13653 7412
rect 13611 7363 13653 7372
rect 13708 7337 13748 7615
rect 13707 7328 13749 7337
rect 13707 7288 13708 7328
rect 13748 7288 13749 7328
rect 13707 7279 13749 7288
rect 13420 7244 13460 7253
rect 13420 7001 13460 7204
rect 13611 7244 13653 7253
rect 13611 7204 13612 7244
rect 13652 7204 13653 7244
rect 13611 7195 13653 7204
rect 13612 7110 13652 7195
rect 13419 6992 13461 7001
rect 13419 6952 13420 6992
rect 13460 6952 13461 6992
rect 13419 6943 13461 6952
rect 13707 6152 13749 6161
rect 13707 6112 13708 6152
rect 13748 6112 13749 6152
rect 13707 6103 13749 6112
rect 13708 4976 13748 6103
rect 13900 4985 13940 5070
rect 13708 4927 13748 4936
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 13996 4808 14036 9976
rect 14668 9967 14708 9976
rect 14572 9428 14612 9437
rect 14475 9176 14517 9185
rect 14475 9136 14476 9176
rect 14516 9136 14517 9176
rect 14475 9127 14517 9136
rect 14379 8588 14421 8597
rect 14379 8548 14380 8588
rect 14420 8548 14421 8588
rect 14379 8539 14421 8548
rect 14187 8168 14229 8177
rect 14187 8128 14188 8168
rect 14228 8128 14229 8168
rect 14187 8119 14229 8128
rect 14188 7916 14228 8119
rect 14188 7867 14228 7876
rect 14380 7916 14420 8539
rect 14380 7867 14420 7876
rect 14283 7832 14325 7841
rect 14283 7792 14284 7832
rect 14324 7792 14325 7832
rect 14283 7783 14325 7792
rect 14187 7412 14229 7421
rect 14187 7372 14188 7412
rect 14228 7372 14229 7412
rect 14187 7363 14229 7372
rect 13900 4768 14036 4808
rect 13516 4724 13556 4733
rect 13420 4136 13460 4145
rect 13324 4096 13420 4136
rect 13420 4087 13460 4096
rect 13132 3415 13172 3424
rect 13228 3968 13268 3977
rect 12940 3212 12980 3221
rect 12940 2540 12980 3172
rect 12940 2500 13076 2540
rect 12939 1952 12981 1961
rect 12939 1912 12940 1952
rect 12980 1912 12981 1952
rect 12939 1903 12981 1912
rect 12843 608 12885 617
rect 12843 568 12844 608
rect 12884 568 12885 608
rect 12843 559 12885 568
rect 12940 80 12980 1903
rect 13036 1541 13076 2500
rect 13131 1700 13173 1709
rect 13131 1660 13132 1700
rect 13172 1660 13173 1700
rect 13131 1651 13173 1660
rect 13035 1532 13077 1541
rect 13035 1492 13036 1532
rect 13076 1492 13077 1532
rect 13035 1483 13077 1492
rect 13132 785 13172 1651
rect 13228 1289 13268 3928
rect 13516 3632 13556 4684
rect 13803 4388 13845 4397
rect 13803 4348 13804 4388
rect 13844 4348 13845 4388
rect 13803 4339 13845 4348
rect 13804 4136 13844 4339
rect 13804 4087 13844 4096
rect 13420 3592 13556 3632
rect 13612 3968 13652 3977
rect 13324 3212 13364 3221
rect 13324 2456 13364 3172
rect 13420 2540 13460 3592
rect 13516 3464 13556 3473
rect 13516 3053 13556 3424
rect 13515 3044 13557 3053
rect 13515 3004 13516 3044
rect 13556 3004 13557 3044
rect 13515 2995 13557 3004
rect 13612 2549 13652 3928
rect 13900 3464 13940 4768
rect 14092 4724 14132 4733
rect 13900 3415 13940 3424
rect 13996 3968 14036 3977
rect 13708 3212 13748 3221
rect 13611 2540 13653 2549
rect 13420 2500 13556 2540
rect 13324 2416 13460 2456
rect 13323 2288 13365 2297
rect 13323 2248 13324 2288
rect 13364 2248 13365 2288
rect 13323 2239 13365 2248
rect 13227 1280 13269 1289
rect 13227 1240 13228 1280
rect 13268 1240 13269 1280
rect 13227 1231 13269 1240
rect 13131 776 13173 785
rect 13131 736 13132 776
rect 13172 736 13173 776
rect 13131 727 13173 736
rect 13131 608 13173 617
rect 13131 568 13132 608
rect 13172 568 13173 608
rect 13131 559 13173 568
rect 13132 80 13172 559
rect 13324 80 13364 2239
rect 13420 1625 13460 2416
rect 13419 1616 13461 1625
rect 13419 1576 13420 1616
rect 13460 1576 13461 1616
rect 13419 1567 13461 1576
rect 13516 80 13556 2500
rect 13611 2500 13612 2540
rect 13652 2500 13653 2540
rect 13708 2540 13748 3172
rect 13899 3128 13941 3137
rect 13899 3088 13900 3128
rect 13940 3088 13941 3128
rect 13899 3079 13941 3088
rect 13900 2885 13940 3079
rect 13899 2876 13941 2885
rect 13899 2836 13900 2876
rect 13940 2836 13941 2876
rect 13899 2827 13941 2836
rect 13708 2500 13844 2540
rect 13611 2491 13653 2500
rect 13707 1280 13749 1289
rect 13707 1240 13708 1280
rect 13748 1240 13749 1280
rect 13707 1231 13749 1240
rect 13708 80 13748 1231
rect 13804 1037 13844 2500
rect 13996 1373 14036 3928
rect 14092 3632 14132 4684
rect 14188 4136 14228 7363
rect 14284 4976 14324 7783
rect 14476 6161 14516 9127
rect 14572 8849 14612 9388
rect 14667 9428 14709 9437
rect 14667 9388 14668 9428
rect 14708 9388 14709 9428
rect 14667 9379 14709 9388
rect 14764 9428 14804 10228
rect 14956 10268 14996 10639
rect 14859 10100 14901 10109
rect 14859 10060 14860 10100
rect 14900 10060 14901 10100
rect 14859 10051 14901 10060
rect 14764 9379 14804 9388
rect 14668 9294 14708 9379
rect 14571 8840 14613 8849
rect 14571 8800 14572 8840
rect 14612 8800 14613 8840
rect 14571 8791 14613 8800
rect 14860 7076 14900 10051
rect 14956 9428 14996 10228
rect 15148 10268 15188 10723
rect 15532 10697 15572 10900
rect 15628 10891 15668 10900
rect 15820 10940 15860 10949
rect 15723 10856 15765 10865
rect 15723 10816 15724 10856
rect 15764 10816 15765 10856
rect 15723 10807 15765 10816
rect 15627 10772 15669 10781
rect 15627 10732 15628 10772
rect 15668 10732 15669 10772
rect 15627 10723 15669 10732
rect 15531 10688 15573 10697
rect 15531 10648 15532 10688
rect 15572 10648 15573 10688
rect 15531 10639 15573 10648
rect 15531 10352 15573 10361
rect 15531 10312 15532 10352
rect 15572 10312 15573 10352
rect 15531 10303 15573 10312
rect 15339 10268 15381 10277
rect 15148 10219 15188 10228
rect 15244 10228 15340 10268
rect 15380 10228 15381 10268
rect 15052 10016 15092 10025
rect 15092 9976 15188 10016
rect 15052 9967 15092 9976
rect 15148 9857 15188 9976
rect 15147 9848 15189 9857
rect 15147 9808 15148 9848
rect 15188 9808 15189 9848
rect 15147 9799 15189 9808
rect 15147 9680 15189 9689
rect 15147 9640 15148 9680
rect 15188 9640 15189 9680
rect 15147 9631 15189 9640
rect 14956 8849 14996 9388
rect 15148 9428 15188 9631
rect 15148 9379 15188 9388
rect 15052 9344 15092 9353
rect 15052 9260 15092 9304
rect 15052 9220 15188 9260
rect 14955 8840 14997 8849
rect 14955 8800 14956 8840
rect 14996 8800 14997 8840
rect 14955 8791 14997 8800
rect 14860 7036 14996 7076
rect 14475 6152 14517 6161
rect 14475 6112 14476 6152
rect 14516 6112 14517 6152
rect 14475 6103 14517 6112
rect 14763 6152 14805 6161
rect 14763 6112 14764 6152
rect 14804 6112 14805 6152
rect 14763 6103 14805 6112
rect 14284 4927 14324 4936
rect 14667 4976 14709 4985
rect 14667 4936 14668 4976
rect 14708 4936 14709 4976
rect 14667 4927 14709 4936
rect 14668 4842 14708 4927
rect 14188 4087 14228 4096
rect 14476 4724 14516 4733
rect 14187 3968 14229 3977
rect 14187 3928 14188 3968
rect 14228 3928 14229 3968
rect 14187 3919 14229 3928
rect 14380 3968 14420 3977
rect 14188 3716 14228 3919
rect 14188 3676 14324 3716
rect 14092 3592 14228 3632
rect 14091 3212 14133 3221
rect 14091 3172 14092 3212
rect 14132 3172 14133 3212
rect 14091 3163 14133 3172
rect 14092 3078 14132 3163
rect 14188 2540 14228 3592
rect 14284 3464 14324 3676
rect 14284 3415 14324 3424
rect 14380 3389 14420 3928
rect 14476 3632 14516 4684
rect 14667 4556 14709 4565
rect 14667 4516 14668 4556
rect 14708 4516 14709 4556
rect 14667 4507 14709 4516
rect 14571 4220 14613 4229
rect 14571 4180 14572 4220
rect 14612 4180 14613 4220
rect 14571 4171 14613 4180
rect 14572 4136 14612 4171
rect 14572 4085 14612 4096
rect 14476 3592 14612 3632
rect 14379 3380 14421 3389
rect 14379 3340 14380 3380
rect 14420 3340 14421 3380
rect 14379 3331 14421 3340
rect 14379 3212 14421 3221
rect 14379 3172 14380 3212
rect 14420 3172 14421 3212
rect 14379 3163 14421 3172
rect 14476 3212 14516 3221
rect 14092 2500 14228 2540
rect 13995 1364 14037 1373
rect 13995 1324 13996 1364
rect 14036 1324 14037 1364
rect 13995 1315 14037 1324
rect 13803 1028 13845 1037
rect 13803 988 13804 1028
rect 13844 988 13845 1028
rect 13803 979 13845 988
rect 13899 524 13941 533
rect 13899 484 13900 524
rect 13940 484 13941 524
rect 13899 475 13941 484
rect 13900 80 13940 475
rect 14092 80 14132 2500
rect 14283 2456 14325 2465
rect 14283 2416 14284 2456
rect 14324 2416 14325 2456
rect 14283 2407 14325 2416
rect 14284 80 14324 2407
rect 14380 1121 14420 3163
rect 14476 1709 14516 3172
rect 14572 2540 14612 3592
rect 14668 3464 14708 4507
rect 14764 4145 14804 6103
rect 14860 4724 14900 4733
rect 14763 4136 14805 4145
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 14763 3968 14805 3977
rect 14763 3928 14764 3968
rect 14804 3928 14805 3968
rect 14763 3919 14805 3928
rect 14764 3834 14804 3919
rect 14860 3632 14900 4684
rect 14956 4136 14996 7036
rect 15148 6581 15188 9220
rect 15244 8924 15284 10228
rect 15339 10219 15381 10228
rect 15532 10268 15572 10303
rect 15340 10134 15380 10219
rect 15435 10100 15477 10109
rect 15435 10060 15436 10100
rect 15476 10060 15477 10100
rect 15435 10051 15477 10060
rect 15436 9966 15476 10051
rect 15340 9428 15380 9437
rect 15340 9092 15380 9388
rect 15532 9428 15572 10228
rect 15628 9428 15668 10723
rect 15724 10722 15764 10807
rect 15723 10268 15765 10277
rect 15723 10228 15724 10268
rect 15764 10228 15765 10268
rect 15820 10268 15860 10900
rect 17260 10940 17300 11320
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 28108 11360 28148 14920
rect 28395 11444 28437 11453
rect 28395 11404 28396 11444
rect 28436 11404 28437 11444
rect 28395 11395 28437 11404
rect 28108 11320 28244 11360
rect 18808 11311 19176 11320
rect 19563 11108 19605 11117
rect 19563 11068 19564 11108
rect 19604 11068 19605 11108
rect 19563 11059 19605 11068
rect 21195 11108 21237 11117
rect 21195 11068 21196 11108
rect 21236 11068 21237 11108
rect 21195 11059 21237 11068
rect 24363 11108 24405 11117
rect 25419 11108 25461 11117
rect 24363 11068 24364 11108
rect 24404 11068 24405 11108
rect 24363 11059 24405 11068
rect 24556 11068 24980 11108
rect 19275 11024 19317 11033
rect 19275 10984 19276 11024
rect 19316 10984 19317 11024
rect 19275 10975 19317 10984
rect 17260 10891 17300 10900
rect 17451 10940 17493 10949
rect 17451 10900 17452 10940
rect 17492 10900 17493 10940
rect 17451 10891 17493 10900
rect 17452 10806 17492 10891
rect 18603 10772 18645 10781
rect 18603 10732 18604 10772
rect 18644 10732 18645 10772
rect 18603 10723 18645 10732
rect 16299 10436 16341 10445
rect 16299 10396 16300 10436
rect 16340 10396 16341 10436
rect 16299 10387 16341 10396
rect 15915 10268 15957 10277
rect 15820 10228 15916 10268
rect 15956 10228 15957 10268
rect 15723 10219 15765 10228
rect 15915 10219 15957 10228
rect 16107 10268 16149 10277
rect 16107 10228 16108 10268
rect 16148 10228 16149 10268
rect 16107 10219 16149 10228
rect 16300 10268 16340 10387
rect 16300 10219 16340 10228
rect 18604 10268 18644 10723
rect 19083 10688 19125 10697
rect 19083 10648 19084 10688
rect 19124 10648 19125 10688
rect 19083 10639 19125 10648
rect 18795 10436 18837 10445
rect 18795 10396 18796 10436
rect 18836 10396 18837 10436
rect 18795 10387 18837 10396
rect 18604 10219 18644 10228
rect 18796 10268 18836 10387
rect 19084 10352 19124 10639
rect 19179 10520 19221 10529
rect 19179 10480 19180 10520
rect 19220 10480 19221 10520
rect 19179 10471 19221 10480
rect 19084 10303 19124 10312
rect 18796 10219 18836 10228
rect 18988 10268 19028 10277
rect 15724 9848 15764 10219
rect 15916 10134 15956 10219
rect 16108 10134 16148 10219
rect 17643 10184 17685 10193
rect 17643 10144 17644 10184
rect 17684 10144 17685 10184
rect 17643 10135 17685 10144
rect 16203 10100 16245 10109
rect 16203 10060 16204 10100
rect 16244 10060 16245 10100
rect 16203 10051 16245 10060
rect 15820 10016 15860 10025
rect 15860 9976 16052 10016
rect 15820 9967 15860 9976
rect 15724 9808 15956 9848
rect 15916 9437 15956 9808
rect 15724 9428 15764 9437
rect 15628 9388 15724 9428
rect 15532 9379 15572 9388
rect 15724 9379 15764 9388
rect 15915 9428 15957 9437
rect 15915 9388 15916 9428
rect 15956 9388 15957 9428
rect 15915 9379 15957 9388
rect 15435 9344 15477 9353
rect 15435 9304 15436 9344
rect 15476 9304 15477 9344
rect 15435 9295 15477 9304
rect 15820 9344 15860 9353
rect 15436 9210 15476 9295
rect 15340 9052 15476 9092
rect 15340 8924 15380 8933
rect 15244 8884 15340 8924
rect 15340 8875 15380 8884
rect 15436 8849 15476 9052
rect 15531 8924 15573 8933
rect 15531 8884 15532 8924
rect 15572 8884 15573 8924
rect 15531 8875 15573 8884
rect 15435 8840 15477 8849
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 15243 8756 15285 8765
rect 15243 8716 15244 8756
rect 15284 8716 15285 8756
rect 15243 8707 15285 8716
rect 15244 6749 15284 8707
rect 15532 7076 15572 8875
rect 15724 8756 15764 8765
rect 15724 8597 15764 8716
rect 15723 8588 15765 8597
rect 15723 8548 15724 8588
rect 15764 8548 15765 8588
rect 15723 8539 15765 8548
rect 15436 7036 15572 7076
rect 15243 6740 15285 6749
rect 15243 6700 15244 6740
rect 15284 6700 15285 6740
rect 15243 6691 15285 6700
rect 15147 6572 15189 6581
rect 15147 6532 15148 6572
rect 15188 6532 15189 6572
rect 15147 6523 15189 6532
rect 15051 6404 15093 6413
rect 15051 6364 15052 6404
rect 15092 6364 15093 6404
rect 15051 6355 15093 6364
rect 15052 4976 15092 6355
rect 15147 6236 15189 6245
rect 15147 6196 15148 6236
rect 15188 6196 15189 6236
rect 15147 6187 15189 6196
rect 15052 4927 15092 4936
rect 15051 4808 15093 4817
rect 15051 4768 15052 4808
rect 15092 4768 15093 4808
rect 15051 4759 15093 4768
rect 14956 4087 14996 4096
rect 15052 3893 15092 4759
rect 15148 4136 15188 6187
rect 15339 5816 15381 5825
rect 15339 5776 15340 5816
rect 15380 5776 15381 5816
rect 15339 5767 15381 5776
rect 15340 5732 15380 5767
rect 15340 5681 15380 5692
rect 15340 5480 15380 5489
rect 15340 5069 15380 5440
rect 15436 5144 15476 7036
rect 15531 6908 15573 6917
rect 15531 6868 15532 6908
rect 15572 6868 15573 6908
rect 15531 6859 15573 6868
rect 15532 5732 15572 6859
rect 15820 6824 15860 9304
rect 15916 9294 15956 9379
rect 15724 6784 15860 6824
rect 15627 6572 15669 6581
rect 15627 6532 15628 6572
rect 15668 6532 15669 6572
rect 15627 6523 15669 6532
rect 15628 6404 15668 6523
rect 15628 5900 15668 6364
rect 15724 6245 15764 6784
rect 15819 6656 15861 6665
rect 15819 6616 15820 6656
rect 15860 6616 15861 6656
rect 15819 6607 15861 6616
rect 15820 6522 15860 6607
rect 16012 6572 16052 9976
rect 16204 9966 16244 10051
rect 16299 9680 16341 9689
rect 16299 9640 16300 9680
rect 16340 9640 16341 9680
rect 16299 9631 16341 9640
rect 16107 9428 16149 9437
rect 16107 9388 16108 9428
rect 16148 9388 16149 9428
rect 16107 9379 16149 9388
rect 16300 9428 16340 9631
rect 16300 9379 16340 9388
rect 16108 9294 16148 9379
rect 16204 9344 16244 9353
rect 16204 6749 16244 9304
rect 16299 8840 16341 8849
rect 16299 8800 16300 8840
rect 16340 8800 16341 8840
rect 16299 8791 16341 8800
rect 16779 8840 16821 8849
rect 16779 8800 16780 8840
rect 16820 8800 16821 8840
rect 16779 8791 16821 8800
rect 16300 8000 16340 8791
rect 16300 7951 16340 7960
rect 16587 6908 16629 6917
rect 16587 6868 16588 6908
rect 16628 6868 16629 6908
rect 16587 6859 16629 6868
rect 16203 6740 16245 6749
rect 16203 6700 16204 6740
rect 16244 6700 16245 6740
rect 16203 6691 16245 6700
rect 16396 6581 16436 6666
rect 15916 6532 16052 6572
rect 16395 6572 16437 6581
rect 16395 6532 16396 6572
rect 16436 6532 16437 6572
rect 15819 6404 15861 6413
rect 15819 6364 15820 6404
rect 15860 6364 15861 6404
rect 15819 6355 15861 6364
rect 15820 6270 15860 6355
rect 15723 6236 15765 6245
rect 15723 6196 15724 6236
rect 15764 6196 15765 6236
rect 15723 6187 15765 6196
rect 15916 5993 15956 6532
rect 16395 6523 16437 6532
rect 16011 6404 16053 6413
rect 16011 6364 16012 6404
rect 16052 6364 16053 6404
rect 16011 6355 16053 6364
rect 16209 6404 16249 6410
rect 16299 6404 16341 6413
rect 16396 6404 16436 6413
rect 16209 6401 16300 6404
rect 16249 6364 16300 6401
rect 16340 6364 16345 6404
rect 16012 6270 16052 6355
rect 16209 6352 16249 6361
rect 16299 6355 16345 6364
rect 16107 6320 16149 6329
rect 16107 6280 16108 6320
rect 16148 6280 16149 6320
rect 16107 6271 16149 6280
rect 16108 6186 16148 6271
rect 16305 6236 16345 6355
rect 16396 6329 16436 6364
rect 16588 6404 16628 6859
rect 16588 6355 16628 6364
rect 16396 6320 16438 6329
rect 16396 6280 16397 6320
rect 16437 6280 16438 6320
rect 16396 6271 16438 6280
rect 16300 6196 16345 6236
rect 16011 6068 16053 6077
rect 16011 6028 16012 6068
rect 16052 6028 16053 6068
rect 16011 6019 16053 6028
rect 15915 5984 15957 5993
rect 15915 5944 15916 5984
rect 15956 5944 15957 5984
rect 15915 5935 15957 5944
rect 15628 5860 15860 5900
rect 15532 5683 15572 5692
rect 15724 5732 15764 5743
rect 15820 5732 15860 5860
rect 15916 5732 15956 5741
rect 15820 5692 15916 5732
rect 15724 5657 15764 5692
rect 15916 5683 15956 5692
rect 15723 5648 15765 5657
rect 15723 5608 15724 5648
rect 15764 5608 15860 5648
rect 15723 5599 15765 5608
rect 15724 5480 15764 5489
rect 15724 5153 15764 5440
rect 15723 5144 15765 5153
rect 15436 5104 15572 5144
rect 15532 5069 15572 5104
rect 15723 5104 15724 5144
rect 15764 5104 15765 5144
rect 15723 5095 15765 5104
rect 15339 5060 15381 5069
rect 15339 5020 15340 5060
rect 15380 5020 15381 5060
rect 15532 5060 15576 5069
rect 15532 5020 15535 5060
rect 15575 5020 15576 5060
rect 15339 5011 15381 5020
rect 15534 5011 15576 5020
rect 15436 4976 15476 4987
rect 15436 4901 15476 4936
rect 15435 4892 15477 4901
rect 15435 4852 15436 4892
rect 15476 4852 15477 4892
rect 15435 4843 15477 4852
rect 15820 4892 15860 5608
rect 15820 4843 15860 4852
rect 16012 4892 16052 6019
rect 16107 5816 16149 5825
rect 16107 5776 16108 5816
rect 16148 5776 16149 5816
rect 16107 5767 16149 5776
rect 16108 5732 16148 5767
rect 16108 5681 16148 5692
rect 16300 5732 16340 6196
rect 16683 6068 16725 6077
rect 16683 6028 16684 6068
rect 16724 6028 16725 6068
rect 16683 6019 16725 6028
rect 16395 5984 16437 5993
rect 16395 5944 16396 5984
rect 16436 5944 16437 5984
rect 16395 5935 16437 5944
rect 16300 5683 16340 5692
rect 16108 5480 16148 5489
rect 16108 5321 16148 5440
rect 16107 5312 16149 5321
rect 16107 5272 16108 5312
rect 16148 5272 16149 5312
rect 16107 5263 16149 5272
rect 16299 5228 16341 5237
rect 16299 5188 16300 5228
rect 16340 5188 16341 5228
rect 16299 5179 16341 5188
rect 16107 5060 16149 5069
rect 16107 5020 16108 5060
rect 16148 5020 16149 5060
rect 16107 5011 16149 5020
rect 16012 4843 16052 4852
rect 15244 4724 15284 4733
rect 15627 4724 15669 4733
rect 15916 4724 15956 4733
rect 15284 4684 15476 4724
rect 15244 4675 15284 4684
rect 15340 4136 15380 4145
rect 15148 4096 15340 4136
rect 15340 4087 15380 4096
rect 15148 3968 15188 3977
rect 15188 3928 15380 3968
rect 15148 3919 15188 3928
rect 15051 3884 15093 3893
rect 15051 3844 15052 3884
rect 15092 3844 15093 3884
rect 15051 3835 15093 3844
rect 15147 3800 15189 3809
rect 15147 3760 15148 3800
rect 15188 3760 15189 3800
rect 15147 3751 15189 3760
rect 15051 3716 15093 3725
rect 15051 3676 15052 3716
rect 15092 3676 15093 3716
rect 15051 3667 15093 3676
rect 14860 3592 14996 3632
rect 14668 3415 14708 3424
rect 14763 3380 14805 3389
rect 14763 3340 14764 3380
rect 14804 3340 14805 3380
rect 14763 3331 14805 3340
rect 14572 2500 14708 2540
rect 14475 1700 14517 1709
rect 14475 1660 14476 1700
rect 14516 1660 14517 1700
rect 14475 1651 14517 1660
rect 14475 1532 14517 1541
rect 14475 1492 14476 1532
rect 14516 1492 14517 1532
rect 14475 1483 14517 1492
rect 14379 1112 14421 1121
rect 14379 1072 14380 1112
rect 14420 1072 14421 1112
rect 14379 1063 14421 1072
rect 14476 80 14516 1483
rect 14668 80 14708 2500
rect 14764 1289 14804 3331
rect 14860 3212 14900 3221
rect 14860 1541 14900 3172
rect 14956 2540 14996 3592
rect 15052 3464 15092 3667
rect 15052 3415 15092 3424
rect 15148 3305 15188 3751
rect 15147 3296 15189 3305
rect 15147 3256 15148 3296
rect 15188 3256 15189 3296
rect 15147 3247 15189 3256
rect 15244 3212 15284 3221
rect 14956 2500 15188 2540
rect 15051 1616 15093 1625
rect 15051 1576 15052 1616
rect 15092 1576 15093 1616
rect 15051 1567 15093 1576
rect 14859 1532 14901 1541
rect 14859 1492 14860 1532
rect 14900 1492 14901 1532
rect 14859 1483 14901 1492
rect 14859 1364 14901 1373
rect 14859 1324 14860 1364
rect 14900 1324 14901 1364
rect 14859 1315 14901 1324
rect 14763 1280 14805 1289
rect 14763 1240 14764 1280
rect 14804 1240 14805 1280
rect 14763 1231 14805 1240
rect 14860 80 14900 1315
rect 15052 80 15092 1567
rect 15148 1280 15188 2500
rect 15244 1625 15284 3172
rect 15243 1616 15285 1625
rect 15243 1576 15244 1616
rect 15284 1576 15285 1616
rect 15243 1567 15285 1576
rect 15148 1240 15284 1280
rect 15244 80 15284 1240
rect 15340 1205 15380 3928
rect 15436 3725 15476 4684
rect 15627 4684 15628 4724
rect 15668 4684 15669 4724
rect 15627 4675 15669 4684
rect 15724 4684 15916 4724
rect 15628 4590 15668 4675
rect 15724 4472 15764 4684
rect 15916 4675 15956 4684
rect 15628 4432 15764 4472
rect 15532 3968 15572 3977
rect 15435 3716 15477 3725
rect 15435 3676 15436 3716
rect 15476 3676 15477 3716
rect 15435 3667 15477 3676
rect 15436 3464 15476 3473
rect 15436 3221 15476 3424
rect 15435 3212 15477 3221
rect 15435 3172 15436 3212
rect 15476 3172 15477 3212
rect 15435 3163 15477 3172
rect 15532 2633 15572 3928
rect 15628 3809 15668 4432
rect 15723 4304 15765 4313
rect 15723 4264 15724 4304
rect 15764 4264 15765 4304
rect 15723 4255 15765 4264
rect 15724 4136 15764 4255
rect 15724 4087 15764 4096
rect 16108 4136 16148 5011
rect 16300 4472 16340 5179
rect 16396 4976 16436 5935
rect 16492 5741 16532 5826
rect 16491 5732 16533 5741
rect 16491 5692 16492 5732
rect 16532 5692 16533 5732
rect 16491 5683 16533 5692
rect 16684 5732 16724 6019
rect 16684 5683 16724 5692
rect 16491 5480 16533 5489
rect 16491 5440 16492 5480
rect 16532 5440 16533 5480
rect 16491 5431 16533 5440
rect 16492 5346 16532 5431
rect 16780 5228 16820 8791
rect 17164 7916 17204 7925
rect 17164 7253 17204 7876
rect 17163 7244 17205 7253
rect 17163 7204 17164 7244
rect 17204 7204 17205 7244
rect 17163 7195 17205 7204
rect 17259 6320 17301 6329
rect 17259 6280 17260 6320
rect 17300 6280 17301 6320
rect 17259 6271 17301 6280
rect 17067 5984 17109 5993
rect 17067 5944 17068 5984
rect 17108 5944 17109 5984
rect 17067 5935 17109 5944
rect 16971 5900 17013 5909
rect 16971 5860 16972 5900
rect 17012 5860 17013 5900
rect 16971 5851 17013 5860
rect 16875 5816 16917 5825
rect 16875 5776 16876 5816
rect 16916 5776 16917 5816
rect 16875 5767 16917 5776
rect 16684 5188 16820 5228
rect 16876 5732 16916 5767
rect 16972 5766 17012 5851
rect 16491 5144 16533 5153
rect 16491 5104 16492 5144
rect 16532 5104 16533 5144
rect 16491 5095 16533 5104
rect 16396 4927 16436 4936
rect 16108 4087 16148 4096
rect 16204 4432 16340 4472
rect 15916 3968 15956 3977
rect 15916 3809 15956 3928
rect 16107 3968 16149 3977
rect 16107 3928 16108 3968
rect 16148 3928 16149 3968
rect 16107 3919 16149 3928
rect 15627 3800 15669 3809
rect 15627 3760 15628 3800
rect 15668 3760 15669 3800
rect 15627 3751 15669 3760
rect 15915 3800 15957 3809
rect 15915 3760 15916 3800
rect 15956 3760 15957 3800
rect 15915 3751 15957 3760
rect 15723 3716 15765 3725
rect 15723 3676 15724 3716
rect 15764 3676 15765 3716
rect 15723 3667 15765 3676
rect 15628 3212 15668 3221
rect 15531 2624 15573 2633
rect 15531 2584 15532 2624
rect 15572 2584 15573 2624
rect 15531 2575 15573 2584
rect 15628 1373 15668 3172
rect 15724 2540 15764 3667
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 15820 3330 15860 3415
rect 15915 3380 15957 3389
rect 15915 3340 15916 3380
rect 15956 3340 15957 3380
rect 15915 3331 15957 3340
rect 15916 3221 15956 3331
rect 15915 3212 15957 3221
rect 15915 3172 15916 3212
rect 15956 3172 15957 3212
rect 15915 3163 15957 3172
rect 16012 3212 16052 3221
rect 16012 2540 16052 3172
rect 15724 2500 15860 2540
rect 15627 1364 15669 1373
rect 15627 1324 15628 1364
rect 15668 1324 15669 1364
rect 15627 1315 15669 1324
rect 15435 1280 15477 1289
rect 15435 1240 15436 1280
rect 15476 1240 15477 1280
rect 15435 1231 15477 1240
rect 15339 1196 15381 1205
rect 15339 1156 15340 1196
rect 15380 1156 15381 1196
rect 15339 1147 15381 1156
rect 15436 80 15476 1231
rect 15627 1028 15669 1037
rect 15627 988 15628 1028
rect 15668 988 15669 1028
rect 15627 979 15669 988
rect 15628 80 15668 979
rect 15820 80 15860 2500
rect 15916 2500 16052 2540
rect 15916 365 15956 2500
rect 16108 1280 16148 3919
rect 16204 3464 16244 4432
rect 16492 4136 16532 5095
rect 16492 4087 16532 4096
rect 16588 4724 16628 4733
rect 16588 3977 16628 4684
rect 16684 4136 16724 5188
rect 16779 5060 16821 5069
rect 16779 5020 16780 5060
rect 16820 5020 16821 5060
rect 16779 5011 16821 5020
rect 16780 4976 16820 5011
rect 16780 4925 16820 4936
rect 16876 4220 16916 5692
rect 17068 5732 17108 5935
rect 17163 5900 17205 5909
rect 17163 5860 17164 5900
rect 17204 5860 17205 5900
rect 17163 5851 17205 5860
rect 17068 5683 17108 5692
rect 17164 5564 17204 5851
rect 17260 5741 17300 6271
rect 17451 5984 17493 5993
rect 17451 5944 17452 5984
rect 17492 5944 17493 5984
rect 17451 5935 17493 5944
rect 17259 5732 17301 5741
rect 17259 5692 17260 5732
rect 17300 5692 17301 5732
rect 17259 5683 17301 5692
rect 17452 5732 17492 5935
rect 17452 5683 17492 5692
rect 17644 5648 17684 10135
rect 18988 10109 19028 10228
rect 19180 10268 19220 10471
rect 19180 10193 19220 10228
rect 19179 10184 19221 10193
rect 19179 10144 19180 10184
rect 19220 10144 19221 10184
rect 19179 10135 19221 10144
rect 18987 10100 19029 10109
rect 19180 10104 19220 10135
rect 18987 10060 18988 10100
rect 19028 10060 19029 10100
rect 18987 10051 19029 10060
rect 18700 10016 18740 10025
rect 18700 9521 18740 9976
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19179 9680 19221 9689
rect 19179 9640 19180 9680
rect 19220 9640 19221 9680
rect 19179 9631 19221 9640
rect 18699 9512 18741 9521
rect 18699 9472 18700 9512
rect 18740 9472 18741 9512
rect 18699 9463 18741 9472
rect 18987 9428 19029 9437
rect 18987 9388 18988 9428
rect 19028 9388 19029 9428
rect 18987 9379 19029 9388
rect 19180 9428 19220 9631
rect 19180 9379 19220 9388
rect 18988 9294 19028 9379
rect 19084 9344 19124 9353
rect 18411 9008 18453 9017
rect 18411 8968 18412 9008
rect 18452 8968 18453 9008
rect 18411 8959 18453 8968
rect 17835 8336 17877 8345
rect 17835 8296 17836 8336
rect 17876 8296 17877 8336
rect 17835 8287 17877 8296
rect 17836 8093 17876 8287
rect 17835 8084 17877 8093
rect 17835 8044 17836 8084
rect 17876 8044 17877 8084
rect 17835 8035 17877 8044
rect 17836 7916 17876 8035
rect 17836 7867 17876 7876
rect 18027 7916 18069 7925
rect 18027 7876 18028 7916
rect 18068 7876 18069 7916
rect 18027 7867 18069 7876
rect 18219 7916 18261 7925
rect 18219 7876 18220 7916
rect 18260 7876 18261 7916
rect 18219 7867 18261 7876
rect 18412 7916 18452 8959
rect 19084 8849 19124 9304
rect 19276 9092 19316 10975
rect 19564 10974 19604 11059
rect 19468 10940 19508 10949
rect 19372 10268 19412 10277
rect 19468 10268 19508 10900
rect 19660 10940 19700 10949
rect 19563 10856 19605 10865
rect 19563 10816 19564 10856
rect 19604 10816 19605 10856
rect 19563 10807 19605 10816
rect 19564 10688 19604 10807
rect 19660 10781 19700 10900
rect 19947 10940 19989 10949
rect 19947 10900 19948 10940
rect 19988 10900 19989 10940
rect 19947 10891 19989 10900
rect 19659 10772 19701 10781
rect 19659 10732 19660 10772
rect 19700 10732 19701 10772
rect 19659 10723 19701 10732
rect 19563 10648 19604 10688
rect 19563 10352 19603 10648
rect 19948 10613 19988 10891
rect 19947 10604 19989 10613
rect 19947 10564 19948 10604
rect 19988 10564 19989 10604
rect 19947 10555 19989 10564
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 19851 10520 19893 10529
rect 19851 10480 19852 10520
rect 19892 10480 19893 10520
rect 19851 10471 19893 10480
rect 19852 10352 19892 10471
rect 19948 10436 19988 10555
rect 19948 10396 20084 10436
rect 19563 10312 19604 10352
rect 19412 10228 19508 10268
rect 19564 10268 19604 10312
rect 19852 10303 19892 10312
rect 19372 10109 19412 10228
rect 19371 10100 19413 10109
rect 19371 10060 19372 10100
rect 19412 10060 19413 10100
rect 19371 10051 19413 10060
rect 19372 9437 19412 10051
rect 19468 10016 19508 10025
rect 19468 9521 19508 9976
rect 19564 9773 19604 10228
rect 19756 10268 19796 10277
rect 19756 10109 19796 10228
rect 19947 10268 19989 10277
rect 19947 10228 19948 10268
rect 19988 10228 19989 10268
rect 19947 10219 19989 10228
rect 19948 10134 19988 10219
rect 19755 10100 19797 10109
rect 19755 10060 19756 10100
rect 19796 10060 19797 10100
rect 19755 10051 19797 10060
rect 20044 9848 20084 10396
rect 20331 10352 20373 10361
rect 20331 10312 20332 10352
rect 20372 10312 20373 10352
rect 20331 10303 20373 10312
rect 20332 10268 20372 10303
rect 20131 10253 20171 10262
rect 20332 10217 20372 10228
rect 20131 10109 20171 10213
rect 20130 10100 20172 10109
rect 20130 10060 20131 10100
rect 20171 10060 20172 10100
rect 20130 10051 20172 10060
rect 20236 10016 20276 10025
rect 20276 9976 20564 10016
rect 20236 9967 20276 9976
rect 19756 9808 20084 9848
rect 19563 9764 19605 9773
rect 19563 9724 19564 9764
rect 19604 9724 19605 9764
rect 19563 9715 19605 9724
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19467 9463 19509 9472
rect 19371 9428 19413 9437
rect 19371 9388 19372 9428
rect 19412 9388 19413 9428
rect 19371 9379 19413 9388
rect 19564 9428 19604 9437
rect 19372 9294 19412 9379
rect 19467 9344 19509 9353
rect 19467 9304 19468 9344
rect 19508 9304 19509 9344
rect 19467 9295 19509 9304
rect 19468 9210 19508 9295
rect 19564 9092 19604 9388
rect 19756 9428 19796 9808
rect 19756 9379 19796 9388
rect 19947 9428 19989 9437
rect 19947 9388 19948 9428
rect 19988 9388 19989 9428
rect 19947 9379 19989 9388
rect 19276 9052 19604 9092
rect 19852 9344 19892 9353
rect 18699 8840 18741 8849
rect 18699 8800 18700 8840
rect 18740 8800 18741 8840
rect 18699 8791 18741 8800
rect 19083 8840 19125 8849
rect 19083 8800 19084 8840
rect 19124 8800 19125 8840
rect 19083 8791 19125 8800
rect 18603 8756 18645 8765
rect 18603 8716 18604 8756
rect 18644 8716 18645 8756
rect 18603 8707 18645 8716
rect 18604 8429 18644 8707
rect 18700 8706 18740 8791
rect 18796 8756 18836 8767
rect 18796 8681 18836 8716
rect 18795 8672 18837 8681
rect 18795 8632 18796 8672
rect 18836 8632 18837 8672
rect 18795 8623 18837 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 18603 8420 18645 8429
rect 18603 8380 18604 8420
rect 18644 8380 18645 8420
rect 18603 8371 18645 8380
rect 19275 8420 19317 8429
rect 19275 8380 19276 8420
rect 19316 8380 19317 8420
rect 19275 8371 19317 8380
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18795 8168 18837 8177
rect 18795 8128 18796 8168
rect 18836 8128 18837 8168
rect 18795 8119 18837 8128
rect 19179 8168 19221 8177
rect 19179 8128 19180 8168
rect 19220 8128 19221 8168
rect 19179 8119 19221 8128
rect 17931 7832 17973 7841
rect 17931 7792 17932 7832
rect 17972 7792 17973 7832
rect 17931 7783 17973 7792
rect 17932 7698 17972 7783
rect 18028 7782 18068 7867
rect 18220 7782 18260 7867
rect 18316 7832 18356 7841
rect 17739 6908 17781 6917
rect 17739 6868 17740 6908
rect 17780 6868 17781 6908
rect 17739 6859 17781 6868
rect 17740 6404 17780 6859
rect 18219 6656 18261 6665
rect 18219 6616 18220 6656
rect 18260 6616 18261 6656
rect 18219 6607 18261 6616
rect 17740 6355 17780 6364
rect 17932 6404 17972 6413
rect 18124 6404 18164 6413
rect 17972 6364 18124 6404
rect 18220 6404 18260 6607
rect 18316 6581 18356 7792
rect 18412 7505 18452 7876
rect 18603 7916 18645 7925
rect 18603 7876 18604 7916
rect 18644 7876 18645 7916
rect 18603 7867 18645 7876
rect 18796 7916 18836 8119
rect 18411 7496 18453 7505
rect 18411 7456 18412 7496
rect 18452 7456 18453 7496
rect 18411 7447 18453 7456
rect 18604 7244 18644 7867
rect 18796 7841 18836 7876
rect 18987 7916 19029 7925
rect 18987 7876 18988 7916
rect 19028 7876 19029 7916
rect 18987 7867 19029 7876
rect 19180 7916 19220 8119
rect 19180 7867 19220 7876
rect 18700 7832 18740 7841
rect 18700 7421 18740 7792
rect 18795 7832 18837 7841
rect 18795 7792 18796 7832
rect 18836 7792 18837 7832
rect 18795 7783 18837 7792
rect 18988 7782 19028 7867
rect 19276 7841 19316 8371
rect 19372 7925 19412 8623
rect 19563 8504 19605 8513
rect 19563 8464 19564 8504
rect 19604 8464 19605 8504
rect 19563 8455 19605 8464
rect 19564 8009 19604 8455
rect 19852 8084 19892 9304
rect 19948 9294 19988 9379
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19660 8044 19892 8084
rect 19563 8000 19605 8009
rect 19563 7960 19564 8000
rect 19604 7960 19605 8000
rect 19563 7951 19605 7960
rect 19371 7916 19413 7925
rect 19371 7876 19372 7916
rect 19412 7876 19413 7916
rect 19371 7867 19413 7876
rect 19564 7916 19604 7951
rect 19084 7832 19124 7841
rect 18891 7748 18933 7757
rect 18891 7708 18892 7748
rect 18932 7708 18933 7748
rect 18891 7699 18933 7708
rect 18892 7589 18932 7699
rect 18891 7580 18933 7589
rect 18891 7540 18892 7580
rect 18932 7540 18933 7580
rect 18891 7531 18933 7540
rect 18699 7412 18741 7421
rect 18699 7372 18700 7412
rect 18740 7372 18741 7412
rect 18699 7363 18741 7372
rect 18700 7244 18740 7253
rect 18604 7204 18700 7244
rect 18700 7195 18740 7204
rect 18892 7244 18932 7531
rect 18892 7195 18932 7204
rect 18796 7001 18836 7086
rect 19084 7085 19124 7792
rect 19275 7832 19317 7841
rect 19275 7792 19276 7832
rect 19316 7792 19317 7832
rect 19275 7783 19317 7792
rect 19372 7782 19412 7867
rect 19564 7866 19604 7876
rect 19468 7832 19508 7841
rect 19275 7496 19317 7505
rect 19275 7456 19276 7496
rect 19316 7456 19317 7496
rect 19275 7447 19317 7456
rect 19083 7076 19125 7085
rect 19083 7036 19084 7076
rect 19124 7036 19125 7076
rect 19083 7027 19125 7036
rect 18795 6992 18837 7001
rect 18795 6952 18796 6992
rect 18836 6952 18837 6992
rect 18795 6943 18837 6952
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18315 6572 18357 6581
rect 18508 6572 18548 6581
rect 18315 6532 18316 6572
rect 18356 6532 18357 6572
rect 18315 6523 18357 6532
rect 18412 6532 18508 6572
rect 18316 6404 18356 6413
rect 18220 6364 18316 6404
rect 17932 6355 17972 6364
rect 17836 6236 17876 6245
rect 17740 5648 17780 5657
rect 17644 5608 17740 5648
rect 17740 5599 17780 5608
rect 17068 5524 17204 5564
rect 17259 5564 17301 5573
rect 17259 5524 17260 5564
rect 17300 5524 17301 5564
rect 17068 4808 17108 5524
rect 17259 5515 17301 5524
rect 17260 5430 17300 5515
rect 17163 5396 17205 5405
rect 17163 5356 17164 5396
rect 17204 5356 17205 5396
rect 17163 5347 17205 5356
rect 17739 5396 17781 5405
rect 17739 5356 17740 5396
rect 17780 5356 17781 5396
rect 17739 5347 17781 5356
rect 17164 4905 17204 5347
rect 17356 4901 17396 4986
rect 17740 4976 17780 5347
rect 17836 5153 17876 6196
rect 18124 5741 18164 6364
rect 18316 6355 18356 6364
rect 18219 6236 18261 6245
rect 18219 6196 18220 6236
rect 18260 6196 18261 6236
rect 18219 6187 18261 6196
rect 18220 6102 18260 6187
rect 18315 5984 18357 5993
rect 18315 5944 18316 5984
rect 18356 5944 18357 5984
rect 18315 5935 18357 5944
rect 18123 5732 18165 5741
rect 18028 5692 18124 5732
rect 18164 5692 18165 5732
rect 17932 5480 17972 5489
rect 17835 5144 17877 5153
rect 17835 5104 17836 5144
rect 17876 5104 17877 5144
rect 17835 5095 17877 5104
rect 17740 4936 17876 4976
rect 17164 4856 17204 4865
rect 17355 4892 17397 4901
rect 17355 4852 17356 4892
rect 17396 4852 17397 4892
rect 17355 4843 17397 4852
rect 17547 4892 17589 4901
rect 17547 4852 17548 4892
rect 17588 4852 17589 4892
rect 17547 4843 17589 4852
rect 17740 4881 17780 4890
rect 17068 4768 17204 4808
rect 16972 4724 17012 4733
rect 17012 4684 17108 4724
rect 16972 4675 17012 4684
rect 16972 4220 17012 4229
rect 16876 4180 16972 4220
rect 16972 4171 17012 4180
rect 16684 4096 16820 4136
rect 16204 3415 16244 3424
rect 16300 3968 16340 3977
rect 16300 1289 16340 3928
rect 16587 3968 16629 3977
rect 16587 3928 16588 3968
rect 16628 3928 16629 3968
rect 16587 3919 16629 3928
rect 16684 3968 16724 3977
rect 16588 3464 16628 3473
rect 16396 3212 16436 3221
rect 16436 3172 16532 3212
rect 16396 3163 16436 3172
rect 16395 2456 16437 2465
rect 16395 2416 16396 2456
rect 16436 2416 16437 2456
rect 16395 2407 16437 2416
rect 16012 1240 16148 1280
rect 16299 1280 16341 1289
rect 16299 1240 16300 1280
rect 16340 1240 16341 1280
rect 15915 356 15957 365
rect 15915 316 15916 356
rect 15956 316 15957 356
rect 15915 307 15957 316
rect 16012 80 16052 1240
rect 16299 1231 16341 1240
rect 16203 1112 16245 1121
rect 16203 1072 16204 1112
rect 16244 1072 16245 1112
rect 16203 1063 16245 1072
rect 16204 80 16244 1063
rect 16396 80 16436 2407
rect 16492 1868 16532 3172
rect 16588 2717 16628 3424
rect 16587 2708 16629 2717
rect 16587 2668 16588 2708
rect 16628 2668 16629 2708
rect 16587 2659 16629 2668
rect 16684 2633 16724 3928
rect 16780 3473 16820 4096
rect 16875 3968 16917 3977
rect 16875 3928 16876 3968
rect 16916 3928 16917 3968
rect 16875 3919 16917 3928
rect 16779 3464 16821 3473
rect 16779 3424 16780 3464
rect 16820 3424 16821 3464
rect 16779 3415 16821 3424
rect 16780 3212 16820 3221
rect 16683 2624 16725 2633
rect 16683 2584 16684 2624
rect 16724 2584 16725 2624
rect 16683 2575 16725 2584
rect 16492 1828 16724 1868
rect 16491 1700 16533 1709
rect 16491 1660 16492 1700
rect 16532 1660 16533 1700
rect 16491 1651 16533 1660
rect 16492 449 16532 1651
rect 16587 1196 16629 1205
rect 16587 1156 16588 1196
rect 16628 1156 16629 1196
rect 16587 1147 16629 1156
rect 16491 440 16533 449
rect 16491 400 16492 440
rect 16532 400 16533 440
rect 16491 391 16533 400
rect 16588 80 16628 1147
rect 16684 953 16724 1828
rect 16683 944 16725 953
rect 16683 904 16684 944
rect 16724 904 16725 944
rect 16683 895 16725 904
rect 16780 617 16820 3172
rect 16876 1205 16916 3919
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 16972 3330 17012 3415
rect 16971 2456 17013 2465
rect 16971 2416 16972 2456
rect 17012 2416 17013 2456
rect 16971 2407 17013 2416
rect 16875 1196 16917 1205
rect 16875 1156 16876 1196
rect 16916 1156 16917 1196
rect 16875 1147 16917 1156
rect 16779 608 16821 617
rect 16779 568 16780 608
rect 16820 568 16821 608
rect 16779 559 16821 568
rect 16779 440 16821 449
rect 16779 400 16780 440
rect 16820 400 16821 440
rect 16779 391 16821 400
rect 16780 80 16820 391
rect 16972 80 17012 2407
rect 17068 869 17108 4684
rect 17164 4649 17204 4768
rect 17548 4758 17588 4843
rect 17260 4724 17300 4733
rect 17163 4640 17205 4649
rect 17163 4600 17164 4640
rect 17204 4600 17205 4640
rect 17163 4591 17205 4600
rect 17164 4220 17204 4591
rect 17164 4171 17204 4180
rect 17260 4052 17300 4684
rect 17644 4724 17684 4733
rect 17355 4640 17397 4649
rect 17355 4600 17356 4640
rect 17396 4600 17397 4640
rect 17355 4591 17397 4600
rect 17356 4220 17396 4591
rect 17547 4472 17589 4481
rect 17547 4432 17548 4472
rect 17588 4432 17589 4472
rect 17547 4423 17589 4432
rect 17548 4231 17588 4423
rect 17644 4229 17684 4684
rect 17740 4649 17780 4841
rect 17739 4640 17781 4649
rect 17739 4600 17740 4640
rect 17780 4600 17781 4640
rect 17739 4591 17781 4600
rect 17548 4182 17588 4191
rect 17643 4220 17685 4229
rect 17356 4171 17396 4180
rect 17643 4180 17644 4220
rect 17684 4180 17685 4220
rect 17643 4171 17685 4180
rect 17740 4136 17780 4145
rect 17164 4012 17300 4052
rect 17643 4052 17685 4061
rect 17643 4012 17644 4052
rect 17684 4012 17685 4052
rect 17164 3473 17204 4012
rect 17643 4003 17685 4012
rect 17356 3968 17396 3977
rect 17260 3928 17356 3968
rect 17163 3464 17205 3473
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 17163 3212 17205 3221
rect 17163 3172 17164 3212
rect 17204 3172 17205 3212
rect 17163 3163 17205 3172
rect 17164 3078 17204 3163
rect 17260 3137 17300 3928
rect 17356 3919 17396 3928
rect 17547 3800 17589 3809
rect 17547 3760 17548 3800
rect 17588 3760 17589 3800
rect 17547 3751 17589 3760
rect 17355 3464 17397 3473
rect 17355 3424 17356 3464
rect 17396 3424 17397 3464
rect 17355 3415 17397 3424
rect 17356 3330 17396 3415
rect 17548 3380 17588 3751
rect 17644 3716 17684 4003
rect 17740 3893 17780 4096
rect 17739 3884 17781 3893
rect 17739 3844 17740 3884
rect 17780 3844 17781 3884
rect 17739 3835 17781 3844
rect 17644 3676 17780 3716
rect 17740 3380 17780 3676
rect 17548 3340 17684 3380
rect 17548 3212 17588 3221
rect 17259 3128 17301 3137
rect 17259 3088 17260 3128
rect 17300 3088 17301 3128
rect 17259 3079 17301 3088
rect 17548 2633 17588 3172
rect 17547 2624 17589 2633
rect 17547 2584 17548 2624
rect 17588 2584 17589 2624
rect 17547 2575 17589 2584
rect 17644 2456 17684 3340
rect 17836 3380 17876 4936
rect 17932 4304 17972 5440
rect 18028 4892 18068 5692
rect 18123 5683 18165 5692
rect 18316 5732 18356 5935
rect 18316 5683 18356 5692
rect 18028 4843 18068 4852
rect 18124 5480 18164 5489
rect 18124 4565 18164 5440
rect 18219 5144 18261 5153
rect 18219 5104 18220 5144
rect 18260 5104 18261 5144
rect 18219 5095 18261 5104
rect 18220 4892 18260 5095
rect 18220 4843 18260 4852
rect 18315 4724 18357 4733
rect 18412 4724 18452 6532
rect 18508 6523 18548 6532
rect 18699 6488 18741 6497
rect 18699 6448 18700 6488
rect 18740 6448 18741 6488
rect 18699 6439 18741 6448
rect 18508 6404 18548 6413
rect 18508 6236 18548 6364
rect 18700 6404 18740 6439
rect 18700 6353 18740 6364
rect 18892 6404 18932 6413
rect 18892 6245 18932 6364
rect 19084 6404 19124 6413
rect 19276 6404 19316 7447
rect 19468 6749 19508 7792
rect 19467 6740 19509 6749
rect 19467 6700 19468 6740
rect 19508 6700 19509 6740
rect 19467 6691 19509 6700
rect 19660 6656 19700 8044
rect 20043 8000 20085 8009
rect 19756 7960 20044 8000
rect 20084 7960 20085 8000
rect 19756 7916 19796 7960
rect 20043 7951 20085 7960
rect 20427 7916 20469 7925
rect 19756 7673 19796 7876
rect 19948 7903 19988 7912
rect 20427 7876 20428 7916
rect 20468 7876 20469 7916
rect 20427 7867 20469 7876
rect 19948 7841 19988 7863
rect 19852 7832 19892 7841
rect 19755 7664 19797 7673
rect 19755 7624 19756 7664
rect 19796 7624 19797 7664
rect 19755 7615 19797 7624
rect 19852 7589 19892 7792
rect 19947 7832 19989 7841
rect 19947 7792 19948 7832
rect 19988 7792 19989 7832
rect 19947 7783 19989 7792
rect 19948 7768 19988 7783
rect 20428 7782 20468 7867
rect 19851 7580 19893 7589
rect 19851 7540 19852 7580
rect 19892 7540 19893 7580
rect 19851 7531 19893 7540
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19564 6616 19700 6656
rect 19467 6572 19509 6581
rect 19467 6532 19468 6572
rect 19508 6532 19509 6572
rect 19467 6523 19509 6532
rect 19468 6488 19508 6523
rect 19468 6437 19508 6448
rect 19124 6364 19316 6404
rect 18603 6236 18645 6245
rect 18508 6196 18604 6236
rect 18644 6196 18645 6236
rect 18603 6187 18645 6196
rect 18891 6236 18933 6245
rect 18891 6196 18892 6236
rect 18932 6196 18933 6236
rect 18891 6187 18933 6196
rect 18988 6236 19028 6245
rect 18604 5741 18644 6187
rect 18988 5900 19028 6196
rect 19084 6077 19124 6364
rect 19276 6236 19316 6245
rect 19179 6152 19221 6161
rect 19179 6112 19180 6152
rect 19220 6112 19221 6152
rect 19179 6103 19221 6112
rect 19083 6068 19125 6077
rect 19083 6028 19084 6068
rect 19124 6028 19125 6068
rect 19083 6019 19125 6028
rect 18892 5860 19028 5900
rect 18603 5732 18645 5741
rect 18603 5692 18604 5732
rect 18644 5692 18645 5732
rect 18603 5683 18645 5692
rect 18795 5732 18837 5741
rect 18795 5692 18796 5732
rect 18836 5692 18837 5732
rect 18795 5683 18837 5692
rect 18796 5598 18836 5683
rect 18892 5489 18932 5860
rect 19083 5816 19125 5825
rect 18988 5776 19084 5816
rect 19124 5776 19125 5816
rect 18988 5732 19028 5776
rect 19083 5767 19125 5776
rect 19180 5741 19220 6103
rect 18988 5683 19028 5692
rect 19179 5732 19221 5741
rect 19179 5692 19180 5732
rect 19220 5692 19221 5732
rect 19179 5683 19221 5692
rect 19084 5648 19124 5657
rect 19084 5489 19124 5608
rect 19180 5598 19220 5683
rect 18604 5480 18644 5489
rect 18507 5396 18549 5405
rect 18507 5356 18508 5396
rect 18548 5356 18549 5396
rect 18507 5347 18549 5356
rect 18508 4892 18548 5347
rect 18604 5069 18644 5440
rect 18891 5480 18933 5489
rect 18891 5440 18892 5480
rect 18932 5440 18933 5480
rect 18891 5431 18933 5440
rect 19083 5480 19125 5489
rect 19083 5440 19084 5480
rect 19124 5440 19125 5480
rect 19083 5431 19125 5440
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18891 5144 18933 5153
rect 18891 5104 18892 5144
rect 18932 5104 18933 5144
rect 18891 5095 18933 5104
rect 18603 5060 18645 5069
rect 18603 5020 18604 5060
rect 18644 5020 18645 5060
rect 18603 5011 18645 5020
rect 18604 4892 18644 4901
rect 18508 4852 18604 4892
rect 18604 4843 18644 4852
rect 18795 4892 18837 4901
rect 18795 4852 18796 4892
rect 18836 4852 18837 4892
rect 18795 4843 18837 4852
rect 18796 4758 18836 4843
rect 18315 4684 18316 4724
rect 18356 4684 18452 4724
rect 18507 4724 18549 4733
rect 18700 4724 18740 4733
rect 18507 4684 18508 4724
rect 18548 4684 18549 4724
rect 18315 4675 18357 4684
rect 18507 4675 18549 4684
rect 18604 4684 18700 4724
rect 18123 4556 18165 4565
rect 18123 4516 18124 4556
rect 18164 4516 18165 4556
rect 18123 4507 18165 4516
rect 17932 4264 18452 4304
rect 18123 4136 18165 4145
rect 18123 4096 18124 4136
rect 18164 4096 18165 4136
rect 18123 4087 18165 4096
rect 18124 4002 18164 4087
rect 17932 3968 17972 3977
rect 18316 3968 18356 3977
rect 17972 3928 18068 3968
rect 17932 3919 17972 3928
rect 17932 3380 17972 3389
rect 17836 3340 17932 3380
rect 17740 3331 17780 3340
rect 17932 3331 17972 3340
rect 17548 2416 17684 2456
rect 17163 1532 17205 1541
rect 17163 1492 17164 1532
rect 17204 1492 17205 1532
rect 17163 1483 17205 1492
rect 17067 860 17109 869
rect 17067 820 17068 860
rect 17108 820 17109 860
rect 17067 811 17109 820
rect 17164 80 17204 1483
rect 17355 1196 17397 1205
rect 17355 1156 17356 1196
rect 17396 1156 17397 1196
rect 17355 1147 17397 1156
rect 17356 80 17396 1147
rect 17548 80 17588 2416
rect 17739 1616 17781 1625
rect 17739 1576 17740 1616
rect 17780 1576 17781 1616
rect 17739 1567 17781 1576
rect 17740 80 17780 1567
rect 17931 860 17973 869
rect 17931 820 17932 860
rect 17972 820 17973 860
rect 17931 811 17973 820
rect 17932 80 17972 811
rect 18028 701 18068 3928
rect 18219 1364 18261 1373
rect 18219 1324 18220 1364
rect 18260 1324 18261 1364
rect 18219 1315 18261 1324
rect 18123 1280 18165 1289
rect 18123 1240 18124 1280
rect 18164 1240 18165 1280
rect 18123 1231 18165 1240
rect 18027 692 18069 701
rect 18027 652 18028 692
rect 18068 652 18069 692
rect 18027 643 18069 652
rect 18124 80 18164 1231
rect 18220 1112 18260 1315
rect 18316 1289 18356 3928
rect 18412 2540 18452 4264
rect 18508 4136 18548 4675
rect 18508 4087 18548 4096
rect 18604 3557 18644 4684
rect 18700 4675 18740 4684
rect 18892 4220 18932 5095
rect 19184 4976 19226 4985
rect 19180 4936 19185 4976
rect 19225 4936 19226 4976
rect 19180 4927 19226 4936
rect 18988 4892 19028 4901
rect 18988 4649 19028 4852
rect 19180 4892 19220 4927
rect 19083 4808 19125 4817
rect 19083 4768 19084 4808
rect 19124 4768 19125 4808
rect 19083 4759 19125 4768
rect 19084 4674 19124 4759
rect 18987 4640 19029 4649
rect 18987 4600 18988 4640
rect 19028 4600 19029 4640
rect 18987 4591 19029 4600
rect 18988 4220 19028 4591
rect 19180 4481 19220 4852
rect 19179 4472 19221 4481
rect 19179 4432 19180 4472
rect 19220 4432 19221 4472
rect 19179 4423 19221 4432
rect 19084 4220 19124 4229
rect 18988 4180 19084 4220
rect 18892 4171 18932 4180
rect 19084 4171 19124 4180
rect 18700 3968 18740 3977
rect 18603 3548 18645 3557
rect 18603 3508 18604 3548
rect 18644 3508 18645 3548
rect 18603 3499 18645 3508
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18508 3330 18548 3415
rect 18700 3380 18740 3928
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3632 19316 6196
rect 19371 6236 19413 6245
rect 19371 6196 19372 6236
rect 19412 6196 19413 6236
rect 19564 6236 19604 6616
rect 19660 6413 19700 6498
rect 19659 6404 19701 6413
rect 19659 6364 19660 6404
rect 19700 6364 19701 6404
rect 19659 6355 19701 6364
rect 19852 6404 19892 6413
rect 20524 6404 20564 9976
rect 20619 9428 20661 9437
rect 20619 9388 20620 9428
rect 20660 9388 20661 9428
rect 20619 9379 20661 9388
rect 20620 8756 20660 9379
rect 21196 8840 21236 11059
rect 24172 10940 24212 10949
rect 24075 10856 24117 10865
rect 24075 10816 24076 10856
rect 24116 10816 24117 10856
rect 24075 10807 24117 10816
rect 21291 10772 21333 10781
rect 21291 10732 21292 10772
rect 21332 10732 21333 10772
rect 21291 10723 21333 10732
rect 21483 10772 21525 10781
rect 21483 10732 21484 10772
rect 21524 10732 21525 10772
rect 21483 10723 21525 10732
rect 21292 10445 21332 10723
rect 21291 10436 21333 10445
rect 21291 10396 21292 10436
rect 21332 10396 21333 10436
rect 21291 10387 21333 10396
rect 21484 10361 21524 10723
rect 23403 10688 23445 10697
rect 23403 10648 23404 10688
rect 23444 10648 23445 10688
rect 23403 10639 23445 10648
rect 23883 10688 23925 10697
rect 23883 10648 23884 10688
rect 23924 10648 23925 10688
rect 23883 10639 23925 10648
rect 21675 10520 21717 10529
rect 21675 10480 21676 10520
rect 21716 10480 21717 10520
rect 21675 10471 21717 10480
rect 21483 10352 21525 10361
rect 21483 10312 21484 10352
rect 21524 10312 21525 10352
rect 21483 10303 21525 10312
rect 21484 10184 21524 10303
rect 21676 10268 21716 10471
rect 21676 10219 21716 10228
rect 21484 10135 21524 10144
rect 21580 10100 21620 10109
rect 21580 9941 21620 10060
rect 21579 9932 21621 9941
rect 21579 9892 21580 9932
rect 21620 9892 21621 9932
rect 21579 9883 21621 9892
rect 21963 9512 22005 9521
rect 21963 9472 21964 9512
rect 22004 9472 22005 9512
rect 21963 9463 22005 9472
rect 21196 8800 21332 8840
rect 20620 8707 20660 8716
rect 20812 8756 20852 8765
rect 20620 7916 20660 7927
rect 20620 7841 20660 7876
rect 20812 7841 20852 8716
rect 20619 7832 20661 7841
rect 20619 7792 20620 7832
rect 20660 7792 20661 7832
rect 20619 7783 20661 7792
rect 20811 7832 20853 7841
rect 20811 7792 20812 7832
rect 20852 7792 20853 7832
rect 20811 7783 20853 7792
rect 21003 7076 21045 7085
rect 21003 7036 21004 7076
rect 21044 7036 21045 7076
rect 21003 7027 21045 7036
rect 20715 6992 20757 7001
rect 20715 6952 20716 6992
rect 20756 6952 20757 6992
rect 20715 6943 20757 6952
rect 20716 6488 20756 6943
rect 20716 6439 20756 6448
rect 19755 6320 19797 6329
rect 19755 6280 19756 6320
rect 19796 6280 19797 6320
rect 19755 6271 19797 6280
rect 19564 6196 19700 6236
rect 19371 6187 19413 6196
rect 19372 5732 19412 6187
rect 19563 5900 19605 5909
rect 19563 5860 19564 5900
rect 19604 5860 19605 5900
rect 19563 5851 19605 5860
rect 19564 5732 19604 5851
rect 19412 5692 19508 5732
rect 19372 5683 19412 5692
rect 19372 5480 19412 5489
rect 19372 5237 19412 5440
rect 19371 5228 19413 5237
rect 19371 5188 19372 5228
rect 19412 5188 19413 5228
rect 19371 5179 19413 5188
rect 19372 4892 19412 4901
rect 19468 4892 19508 5692
rect 19564 5683 19604 5692
rect 19563 5480 19605 5489
rect 19563 5440 19564 5480
rect 19604 5440 19605 5480
rect 19563 5431 19605 5440
rect 19412 4852 19508 4892
rect 19564 4892 19604 5431
rect 19372 4843 19412 4852
rect 19564 4843 19604 4852
rect 19371 4724 19413 4733
rect 19371 4684 19372 4724
rect 19412 4684 19413 4724
rect 19371 4675 19413 4684
rect 19468 4724 19508 4733
rect 19180 3592 19316 3632
rect 18891 3548 18933 3557
rect 18891 3508 18892 3548
rect 18932 3508 18933 3548
rect 18891 3499 18933 3508
rect 18892 3464 18932 3499
rect 18892 3413 18932 3424
rect 18700 3340 18836 3380
rect 18700 3212 18740 3221
rect 18412 2500 18548 2540
rect 18315 1280 18357 1289
rect 18315 1240 18316 1280
rect 18356 1240 18357 1280
rect 18315 1231 18357 1240
rect 18220 1072 18356 1112
rect 18316 80 18356 1072
rect 18508 80 18548 2500
rect 18603 1952 18645 1961
rect 18603 1912 18604 1952
rect 18644 1912 18645 1952
rect 18603 1903 18645 1912
rect 18604 860 18644 1903
rect 18700 1037 18740 3172
rect 18796 1121 18836 3340
rect 19084 3212 19124 3221
rect 19084 1625 19124 3172
rect 19180 2540 19220 3592
rect 19372 3557 19412 4675
rect 19468 4313 19508 4684
rect 19467 4304 19509 4313
rect 19467 4264 19468 4304
rect 19508 4264 19509 4304
rect 19467 4255 19509 4264
rect 19563 4220 19605 4229
rect 19563 4180 19564 4220
rect 19604 4180 19605 4220
rect 19563 4171 19605 4180
rect 19564 4086 19604 4171
rect 19371 3548 19413 3557
rect 19371 3508 19372 3548
rect 19412 3508 19413 3548
rect 19371 3499 19413 3508
rect 19275 3464 19317 3473
rect 19275 3424 19276 3464
rect 19316 3424 19317 3464
rect 19275 3415 19317 3424
rect 19660 3464 19700 6196
rect 19756 6186 19796 6271
rect 19852 6245 19892 6364
rect 20428 6364 20564 6404
rect 20428 6245 20468 6364
rect 19851 6236 19893 6245
rect 19851 6196 19852 6236
rect 19892 6196 19893 6236
rect 19851 6187 19893 6196
rect 20427 6236 20469 6245
rect 20427 6196 20428 6236
rect 20468 6196 20469 6236
rect 20427 6187 20469 6196
rect 20524 6236 20564 6245
rect 20908 6236 20948 6245
rect 20564 6196 20660 6236
rect 20524 6187 20564 6196
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19947 5900 19989 5909
rect 19947 5860 19948 5900
rect 19988 5860 19989 5900
rect 19947 5851 19989 5860
rect 19756 5825 19796 5827
rect 19755 5816 19797 5825
rect 19755 5776 19756 5816
rect 19796 5776 19797 5816
rect 19755 5767 19797 5776
rect 19756 5732 19796 5767
rect 19756 5683 19796 5692
rect 19948 5732 19988 5851
rect 20331 5816 20373 5825
rect 20331 5776 20332 5816
rect 20372 5776 20373 5816
rect 20331 5767 20373 5776
rect 19948 5683 19988 5692
rect 20140 5732 20180 5741
rect 20140 5573 20180 5692
rect 20332 5732 20372 5767
rect 20524 5741 20564 5826
rect 20235 5648 20277 5657
rect 20235 5608 20236 5648
rect 20276 5608 20277 5648
rect 20235 5599 20277 5608
rect 19755 5564 19797 5573
rect 19755 5524 19756 5564
rect 19796 5524 19797 5564
rect 19755 5515 19797 5524
rect 20139 5564 20181 5573
rect 20139 5524 20140 5564
rect 20180 5524 20181 5564
rect 20139 5515 20181 5524
rect 19756 5430 19796 5515
rect 20236 5514 20276 5599
rect 20332 5489 20372 5692
rect 20523 5732 20565 5741
rect 20523 5692 20524 5732
rect 20564 5692 20565 5732
rect 20523 5683 20565 5692
rect 20331 5480 20373 5489
rect 20331 5440 20332 5480
rect 20372 5440 20373 5480
rect 20331 5431 20373 5440
rect 20523 5480 20565 5489
rect 20523 5440 20524 5480
rect 20564 5440 20565 5480
rect 20523 5431 20565 5440
rect 20524 5346 20564 5431
rect 19948 5069 19988 5154
rect 19947 5060 19989 5069
rect 19947 5020 19948 5060
rect 19988 5020 19989 5060
rect 19947 5011 19989 5020
rect 20121 4901 20161 4986
rect 20331 4976 20373 4985
rect 20331 4936 20332 4976
rect 20372 4936 20373 4976
rect 20331 4927 20373 4936
rect 19948 4892 19988 4901
rect 19852 4852 19948 4892
rect 19852 4649 19892 4852
rect 19948 4843 19988 4852
rect 20120 4892 20162 4901
rect 20120 4852 20121 4892
rect 20161 4852 20162 4892
rect 20120 4843 20162 4852
rect 20332 4842 20372 4927
rect 19947 4724 19989 4733
rect 19947 4684 19948 4724
rect 19988 4684 19989 4724
rect 19947 4675 19989 4684
rect 20524 4724 20564 4733
rect 19851 4640 19893 4649
rect 19851 4600 19852 4640
rect 19892 4600 19893 4640
rect 19851 4591 19893 4600
rect 19756 4220 19796 4229
rect 19948 4220 19988 4675
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20331 4304 20373 4313
rect 20331 4264 20332 4304
rect 20372 4264 20373 4304
rect 20331 4255 20373 4264
rect 19796 4180 19948 4220
rect 19756 4171 19796 4180
rect 19948 4171 19988 4180
rect 20144 4220 20186 4229
rect 20144 4180 20145 4220
rect 20185 4180 20186 4220
rect 20144 4171 20186 4180
rect 20145 4086 20185 4171
rect 20332 4136 20372 4255
rect 20524 4229 20564 4684
rect 20523 4220 20565 4229
rect 20523 4180 20524 4220
rect 20564 4180 20565 4220
rect 20523 4171 20565 4180
rect 20332 4087 20372 4096
rect 19755 3968 19797 3977
rect 19755 3928 19756 3968
rect 19796 3928 19797 3968
rect 19755 3919 19797 3928
rect 19947 3968 19989 3977
rect 19947 3928 19948 3968
rect 19988 3928 19989 3968
rect 19947 3919 19989 3928
rect 20524 3968 20564 3977
rect 19756 3834 19796 3919
rect 19948 3834 19988 3919
rect 20427 3884 20469 3893
rect 20427 3844 20428 3884
rect 20468 3844 20469 3884
rect 20427 3835 20469 3844
rect 19660 3415 19700 3424
rect 20043 3464 20085 3473
rect 20043 3424 20044 3464
rect 20084 3424 20085 3464
rect 20043 3415 20085 3424
rect 20428 3464 20468 3835
rect 20524 3557 20564 3928
rect 20523 3548 20565 3557
rect 20523 3508 20524 3548
rect 20564 3508 20565 3548
rect 20523 3499 20565 3508
rect 20428 3415 20468 3424
rect 19276 3330 19316 3415
rect 20044 3330 20084 3415
rect 20620 3380 20660 6196
rect 20715 5816 20757 5825
rect 20715 5776 20716 5816
rect 20756 5776 20757 5816
rect 20715 5767 20757 5776
rect 20716 5732 20756 5767
rect 20716 5681 20756 5692
rect 20715 5312 20757 5321
rect 20715 5272 20716 5312
rect 20756 5272 20757 5312
rect 20715 5263 20757 5272
rect 20716 5060 20756 5263
rect 20908 5237 20948 6196
rect 21004 5648 21044 7027
rect 21099 6740 21141 6749
rect 21099 6700 21100 6740
rect 21140 6700 21141 6740
rect 21099 6691 21141 6700
rect 21100 6488 21140 6691
rect 21100 6439 21140 6448
rect 21004 5599 21044 5608
rect 21196 5480 21236 5489
rect 21004 5440 21196 5480
rect 20907 5228 20949 5237
rect 20907 5188 20908 5228
rect 20948 5188 20949 5228
rect 20907 5179 20949 5188
rect 20715 5020 20756 5060
rect 20715 4963 20755 5020
rect 20715 4923 20756 4963
rect 20716 4905 20756 4923
rect 20716 4733 20756 4865
rect 20907 4892 20949 4901
rect 20907 4852 20908 4892
rect 20948 4852 20949 4892
rect 20907 4843 20949 4852
rect 20812 4808 20852 4817
rect 20715 4724 20757 4733
rect 20715 4684 20716 4724
rect 20756 4684 20757 4724
rect 20715 4675 20757 4684
rect 20715 4556 20757 4565
rect 20715 4516 20716 4556
rect 20756 4516 20757 4556
rect 20715 4507 20757 4516
rect 20716 4136 20756 4507
rect 20812 4481 20852 4768
rect 20908 4758 20948 4843
rect 20811 4472 20853 4481
rect 20811 4432 20812 4472
rect 20852 4432 20853 4472
rect 20811 4423 20853 4432
rect 20716 4087 20756 4096
rect 20908 3968 20948 3977
rect 20524 3340 20660 3380
rect 20716 3928 20908 3968
rect 20236 3221 20276 3306
rect 19468 3212 19508 3221
rect 19180 2500 19316 2540
rect 19083 1616 19125 1625
rect 19083 1576 19084 1616
rect 19124 1576 19125 1616
rect 19083 1567 19125 1576
rect 18795 1112 18837 1121
rect 18795 1072 18796 1112
rect 18836 1072 18837 1112
rect 18795 1063 18837 1072
rect 18699 1028 18741 1037
rect 18699 988 18700 1028
rect 18740 988 18741 1028
rect 18699 979 18741 988
rect 19083 944 19125 953
rect 19083 904 19084 944
rect 19124 904 19125 944
rect 19083 895 19125 904
rect 18604 820 18740 860
rect 18700 80 18740 820
rect 18891 356 18933 365
rect 18891 316 18892 356
rect 18932 316 18933 356
rect 18891 307 18933 316
rect 18892 80 18932 307
rect 19084 80 19124 895
rect 19276 80 19316 2500
rect 19468 1541 19508 3172
rect 19659 3212 19701 3221
rect 19659 3172 19660 3212
rect 19700 3172 19701 3212
rect 19659 3163 19701 3172
rect 19852 3212 19892 3221
rect 19467 1532 19509 1541
rect 19467 1492 19468 1532
rect 19508 1492 19509 1532
rect 19467 1483 19509 1492
rect 19467 608 19509 617
rect 19467 568 19468 608
rect 19508 568 19509 608
rect 19467 559 19509 568
rect 19468 80 19508 559
rect 19660 80 19700 3163
rect 19852 1373 19892 3172
rect 20235 3212 20277 3221
rect 20235 3172 20236 3212
rect 20276 3172 20277 3212
rect 20235 3163 20277 3172
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 20524 2540 20564 3340
rect 20428 2500 20564 2540
rect 20620 3212 20660 3221
rect 20043 2456 20085 2465
rect 20043 2416 20044 2456
rect 20084 2416 20085 2456
rect 20043 2407 20085 2416
rect 19851 1364 19893 1373
rect 19851 1324 19852 1364
rect 19892 1324 19893 1364
rect 19851 1315 19893 1324
rect 19851 692 19893 701
rect 19851 652 19852 692
rect 19892 652 19893 692
rect 19851 643 19893 652
rect 19852 80 19892 643
rect 20044 80 20084 2407
rect 20235 1280 20277 1289
rect 20235 1240 20236 1280
rect 20276 1240 20277 1280
rect 20235 1231 20277 1240
rect 20236 80 20276 1231
rect 20428 80 20468 2500
rect 20620 1877 20660 3172
rect 20619 1868 20661 1877
rect 20619 1828 20620 1868
rect 20660 1828 20661 1868
rect 20619 1819 20661 1828
rect 20619 1112 20661 1121
rect 20619 1072 20620 1112
rect 20660 1072 20661 1112
rect 20619 1063 20661 1072
rect 20620 80 20660 1063
rect 20716 953 20756 3928
rect 20908 3919 20948 3928
rect 20907 3716 20949 3725
rect 20907 3676 20908 3716
rect 20948 3676 20949 3716
rect 20907 3667 20949 3676
rect 20812 3464 20852 3473
rect 20908 3464 20948 3667
rect 20852 3424 20948 3464
rect 20812 3415 20852 3424
rect 21004 3380 21044 5440
rect 21196 5431 21236 5440
rect 21292 5060 21332 8800
rect 21483 6236 21525 6245
rect 21483 6196 21484 6236
rect 21524 6196 21525 6236
rect 21483 6187 21525 6196
rect 21388 5648 21428 5657
rect 21388 5237 21428 5608
rect 21387 5228 21429 5237
rect 21387 5188 21388 5228
rect 21428 5188 21429 5228
rect 21387 5179 21429 5188
rect 21292 5020 21428 5060
rect 21100 4892 21140 4901
rect 21100 4649 21140 4852
rect 21291 4892 21333 4901
rect 21291 4852 21292 4892
rect 21332 4852 21333 4892
rect 21291 4843 21333 4852
rect 21292 4758 21332 4843
rect 21196 4724 21236 4733
rect 21099 4640 21141 4649
rect 21099 4600 21100 4640
rect 21140 4600 21141 4640
rect 21099 4591 21141 4600
rect 21100 4220 21140 4591
rect 21196 4397 21236 4684
rect 21291 4556 21333 4565
rect 21291 4516 21292 4556
rect 21332 4516 21333 4556
rect 21291 4507 21333 4516
rect 21195 4388 21237 4397
rect 21195 4348 21196 4388
rect 21236 4348 21237 4388
rect 21195 4339 21237 4348
rect 21100 4171 21140 4180
rect 21195 4220 21237 4229
rect 21195 4180 21196 4220
rect 21236 4180 21237 4220
rect 21195 4171 21237 4180
rect 21292 4220 21332 4507
rect 21292 4171 21332 4180
rect 21099 4052 21141 4061
rect 21099 4012 21100 4052
rect 21140 4012 21141 4052
rect 21099 4003 21141 4012
rect 21100 3918 21140 4003
rect 21196 3632 21236 4171
rect 21388 3893 21428 5020
rect 21484 4976 21524 6187
rect 21484 4927 21524 4936
rect 21580 5480 21620 5489
rect 21483 4808 21525 4817
rect 21483 4768 21484 4808
rect 21524 4768 21525 4808
rect 21483 4759 21525 4768
rect 21484 4481 21524 4759
rect 21483 4472 21525 4481
rect 21483 4432 21484 4472
rect 21524 4432 21525 4472
rect 21483 4423 21525 4432
rect 21484 4229 21524 4423
rect 21483 4220 21525 4229
rect 21483 4180 21484 4220
rect 21524 4180 21525 4220
rect 21483 4171 21525 4180
rect 21484 3968 21524 3977
rect 21387 3884 21429 3893
rect 21387 3844 21388 3884
rect 21428 3844 21429 3884
rect 21387 3835 21429 3844
rect 21196 3592 21332 3632
rect 21195 3464 21237 3473
rect 21195 3424 21196 3464
rect 21236 3424 21237 3464
rect 21195 3415 21237 3424
rect 21004 3340 21140 3380
rect 20811 3296 20853 3305
rect 20811 3256 20812 3296
rect 20852 3256 20853 3296
rect 20811 3247 20853 3256
rect 20715 944 20757 953
rect 20715 904 20716 944
rect 20756 904 20757 944
rect 20715 895 20757 904
rect 20812 80 20852 3247
rect 21003 3212 21045 3221
rect 21003 3172 21004 3212
rect 21044 3172 21045 3212
rect 21003 3163 21045 3172
rect 20907 3128 20949 3137
rect 20907 3088 20908 3128
rect 20948 3088 20949 3128
rect 20907 3079 20949 3088
rect 20908 1205 20948 3079
rect 21004 3078 21044 3163
rect 21100 2540 21140 3340
rect 21196 3330 21236 3415
rect 21100 2500 21236 2540
rect 20907 1196 20949 1205
rect 20907 1156 20908 1196
rect 20948 1156 20949 1196
rect 20907 1147 20949 1156
rect 21003 1028 21045 1037
rect 21003 988 21004 1028
rect 21044 988 21045 1028
rect 21003 979 21045 988
rect 21004 80 21044 979
rect 21196 80 21236 2500
rect 21292 1280 21332 3592
rect 21388 3212 21428 3221
rect 21388 1364 21428 3172
rect 21484 2549 21524 3928
rect 21580 3800 21620 5440
rect 21964 5069 22004 9463
rect 22347 8588 22389 8597
rect 22347 8548 22348 8588
rect 22388 8548 22389 8588
rect 22347 8539 22389 8548
rect 22348 8084 22388 8539
rect 22348 8035 22388 8044
rect 22636 7925 22676 8010
rect 22540 7916 22580 7925
rect 22540 7673 22580 7876
rect 22635 7916 22677 7925
rect 22635 7876 22636 7916
rect 22676 7876 22677 7916
rect 22635 7867 22677 7876
rect 23212 7916 23252 7927
rect 23308 7925 23348 8010
rect 23212 7841 23252 7876
rect 23307 7916 23349 7925
rect 23307 7876 23308 7916
rect 23348 7876 23349 7916
rect 23307 7867 23349 7876
rect 23019 7832 23061 7841
rect 23019 7792 23020 7832
rect 23060 7792 23061 7832
rect 23019 7783 23061 7792
rect 23211 7832 23253 7841
rect 23211 7792 23212 7832
rect 23252 7792 23253 7832
rect 23211 7783 23253 7792
rect 22636 7748 22676 7757
rect 22539 7664 22581 7673
rect 22539 7624 22540 7664
rect 22580 7624 22581 7664
rect 22539 7615 22581 7624
rect 22636 7421 22676 7708
rect 23020 7698 23060 7783
rect 23308 7748 23348 7757
rect 23020 7421 23060 7506
rect 22635 7412 22677 7421
rect 22635 7372 22636 7412
rect 22676 7372 22677 7412
rect 22635 7363 22677 7372
rect 22827 7412 22869 7421
rect 22827 7372 22828 7412
rect 22868 7372 22869 7412
rect 22827 7363 22869 7372
rect 23019 7412 23061 7421
rect 23308 7412 23348 7708
rect 23019 7372 23020 7412
rect 23060 7372 23348 7412
rect 23019 7363 23061 7372
rect 22731 7244 22773 7253
rect 22731 7204 22732 7244
rect 22772 7204 22773 7244
rect 22731 7195 22773 7204
rect 22732 7110 22772 7195
rect 22732 5732 22772 5741
rect 22732 5573 22772 5692
rect 22828 5732 22868 7363
rect 22923 7244 22965 7253
rect 22923 7204 22924 7244
rect 22964 7204 22965 7244
rect 22923 7195 22965 7204
rect 23020 7244 23060 7253
rect 23115 7244 23157 7253
rect 23060 7204 23116 7244
rect 23156 7204 23157 7244
rect 23020 7195 23060 7204
rect 23115 7195 23157 7204
rect 22924 7110 22964 7195
rect 22923 6404 22965 6413
rect 22923 6364 22924 6404
rect 22964 6364 22965 6404
rect 22923 6355 22965 6364
rect 22924 5993 22964 6355
rect 23116 6152 23156 7195
rect 23211 7160 23253 7169
rect 23211 7120 23212 7160
rect 23252 7120 23253 7160
rect 23211 7111 23253 7120
rect 23212 6413 23252 7111
rect 23308 7085 23348 7372
rect 23307 7076 23349 7085
rect 23307 7036 23308 7076
rect 23348 7036 23349 7076
rect 23307 7027 23349 7036
rect 23404 6749 23444 10639
rect 23787 10604 23829 10613
rect 23787 10564 23788 10604
rect 23828 10564 23829 10604
rect 23787 10555 23829 10564
rect 23788 10268 23828 10555
rect 23884 10352 23924 10639
rect 23884 10303 23924 10312
rect 23788 9773 23828 10228
rect 23980 10268 24020 10277
rect 23980 10109 24020 10228
rect 23979 10100 24021 10109
rect 23979 10060 23980 10100
rect 24020 10060 24021 10100
rect 23979 10051 24021 10060
rect 23787 9764 23829 9773
rect 23787 9724 23788 9764
rect 23828 9724 23829 9764
rect 23787 9715 23829 9724
rect 24076 9689 24116 10807
rect 24172 10268 24212 10900
rect 24364 10940 24404 11059
rect 24459 11024 24501 11033
rect 24459 10984 24460 11024
rect 24500 10984 24501 11024
rect 24459 10975 24501 10984
rect 24364 10865 24404 10900
rect 24172 10109 24212 10228
rect 24268 10856 24308 10865
rect 24268 10184 24308 10816
rect 24363 10856 24405 10865
rect 24363 10816 24364 10856
rect 24404 10816 24405 10856
rect 24363 10807 24405 10816
rect 24460 10688 24500 10975
rect 24364 10648 24500 10688
rect 24556 10940 24596 11068
rect 24364 10289 24404 10648
rect 24364 10240 24404 10249
rect 24556 10268 24596 10900
rect 24747 10940 24789 10949
rect 24747 10900 24748 10940
rect 24788 10900 24789 10940
rect 24747 10891 24789 10900
rect 24940 10940 24980 11068
rect 25419 11068 25420 11108
rect 25460 11068 25461 11108
rect 25419 11059 25461 11068
rect 25420 10949 25460 11059
rect 24940 10891 24980 10900
rect 25132 10940 25172 10949
rect 24652 10856 24692 10865
rect 24652 10604 24692 10816
rect 24748 10806 24788 10891
rect 25036 10856 25076 10865
rect 24652 10564 24980 10604
rect 24843 10436 24885 10445
rect 24843 10396 24844 10436
rect 24884 10396 24885 10436
rect 24843 10387 24885 10396
rect 24268 10144 24500 10184
rect 24171 10100 24213 10109
rect 24171 10060 24172 10100
rect 24212 10060 24213 10100
rect 24171 10051 24213 10060
rect 24075 9680 24117 9689
rect 24075 9640 24076 9680
rect 24116 9640 24117 9680
rect 24075 9631 24117 9640
rect 24172 9437 24212 10051
rect 24268 10016 24308 10025
rect 24268 9605 24308 9976
rect 24363 9932 24405 9941
rect 24363 9892 24364 9932
rect 24404 9892 24405 9932
rect 24363 9883 24405 9892
rect 24267 9596 24309 9605
rect 24267 9556 24268 9596
rect 24308 9556 24309 9596
rect 24267 9547 24309 9556
rect 24171 9428 24213 9437
rect 24171 9388 24172 9428
rect 24212 9388 24213 9428
rect 24171 9379 24213 9388
rect 24364 9428 24404 9883
rect 24364 9379 24404 9388
rect 23499 9344 23541 9353
rect 23499 9304 23500 9344
rect 23540 9304 23541 9344
rect 23499 9295 23541 9304
rect 23403 6740 23445 6749
rect 23403 6700 23404 6740
rect 23444 6700 23445 6740
rect 23403 6691 23445 6700
rect 23211 6404 23253 6413
rect 23211 6364 23212 6404
rect 23252 6364 23253 6404
rect 23211 6355 23253 6364
rect 23403 6404 23445 6413
rect 23403 6364 23404 6404
rect 23444 6364 23445 6404
rect 23403 6355 23445 6364
rect 23212 6270 23252 6355
rect 23404 6270 23444 6355
rect 23308 6236 23348 6245
rect 23116 6112 23252 6152
rect 23019 6068 23061 6077
rect 23019 6028 23020 6068
rect 23060 6028 23061 6068
rect 23019 6019 23061 6028
rect 22923 5984 22965 5993
rect 22923 5944 22924 5984
rect 22964 5944 22965 5984
rect 22923 5935 22965 5944
rect 23020 5900 23060 6019
rect 23115 5984 23157 5993
rect 23115 5944 23116 5984
rect 23156 5944 23157 5984
rect 23115 5935 23157 5944
rect 23020 5851 23060 5860
rect 23020 5732 23060 5741
rect 22828 5692 23020 5732
rect 22731 5564 22773 5573
rect 22731 5524 22732 5564
rect 22772 5524 22773 5564
rect 22731 5515 22773 5524
rect 22444 5480 22484 5489
rect 22484 5440 22580 5480
rect 22444 5431 22484 5440
rect 21963 5060 22005 5069
rect 21963 5020 21964 5060
rect 22004 5020 22005 5060
rect 21963 5011 22005 5020
rect 22443 5060 22485 5069
rect 22443 5020 22444 5060
rect 22484 5020 22485 5060
rect 22443 5011 22485 5020
rect 22252 4901 22292 4986
rect 21867 4892 21909 4901
rect 21867 4852 21868 4892
rect 21908 4852 21909 4892
rect 21867 4843 21909 4852
rect 22060 4892 22100 4901
rect 22251 4892 22293 4901
rect 22100 4852 22196 4892
rect 22060 4843 22100 4852
rect 21868 4758 21908 4843
rect 21676 4724 21716 4733
rect 21964 4724 22004 4733
rect 21716 4684 21812 4724
rect 21676 4675 21716 4684
rect 21675 4472 21717 4481
rect 21675 4432 21676 4472
rect 21716 4432 21717 4472
rect 21675 4423 21717 4432
rect 21676 4220 21716 4423
rect 21676 4171 21716 4180
rect 21580 3760 21716 3800
rect 21579 3548 21621 3557
rect 21579 3508 21580 3548
rect 21620 3508 21621 3548
rect 21579 3499 21621 3508
rect 21580 3464 21620 3499
rect 21580 3413 21620 3424
rect 21483 2540 21525 2549
rect 21483 2500 21484 2540
rect 21524 2500 21525 2540
rect 21676 2540 21716 3760
rect 21772 3557 21812 4684
rect 21964 4472 22004 4684
rect 22156 4565 22196 4852
rect 22251 4852 22252 4892
rect 22292 4852 22293 4892
rect 22251 4843 22293 4852
rect 22444 4892 22484 5011
rect 22444 4843 22484 4852
rect 22540 4817 22580 5440
rect 22828 5396 22868 5692
rect 23020 5683 23060 5692
rect 22636 5356 22868 5396
rect 22636 4892 22676 5356
rect 22923 5312 22965 5321
rect 22923 5272 22924 5312
rect 22964 5272 22965 5312
rect 22923 5263 22965 5272
rect 22827 5144 22869 5153
rect 22827 5104 22828 5144
rect 22868 5104 22869 5144
rect 22827 5095 22869 5104
rect 22828 5010 22868 5095
rect 22636 4843 22676 4852
rect 22828 4892 22868 4901
rect 22539 4808 22581 4817
rect 22539 4768 22540 4808
rect 22580 4768 22581 4808
rect 22539 4759 22581 4768
rect 22828 4733 22868 4852
rect 22924 4892 22964 5263
rect 23019 5144 23061 5153
rect 23019 5104 23020 5144
rect 23060 5104 23061 5144
rect 23019 5095 23061 5104
rect 22924 4843 22964 4852
rect 22347 4724 22389 4733
rect 22347 4684 22348 4724
rect 22388 4684 22389 4724
rect 22347 4675 22389 4684
rect 22827 4724 22869 4733
rect 22827 4684 22828 4724
rect 22868 4684 22869 4724
rect 22827 4675 22869 4684
rect 22251 4640 22293 4649
rect 22251 4600 22252 4640
rect 22292 4600 22293 4640
rect 22251 4591 22293 4600
rect 22155 4556 22197 4565
rect 22155 4516 22156 4556
rect 22196 4516 22197 4556
rect 22155 4507 22197 4516
rect 21964 4432 22100 4472
rect 22060 4388 22100 4432
rect 22060 4348 22196 4388
rect 21868 4229 21908 4314
rect 21867 4220 21909 4229
rect 21867 4180 21868 4220
rect 21908 4180 21909 4220
rect 21867 4171 21909 4180
rect 22060 4220 22100 4229
rect 21868 3968 21908 3977
rect 21771 3548 21813 3557
rect 21771 3508 21772 3548
rect 21812 3508 21813 3548
rect 21771 3499 21813 3508
rect 21868 3296 21908 3928
rect 22060 3893 22100 4180
rect 22059 3884 22101 3893
rect 22059 3844 22060 3884
rect 22100 3844 22101 3884
rect 22059 3835 22101 3844
rect 22156 3632 22196 4348
rect 22252 4229 22292 4591
rect 22348 4590 22388 4675
rect 22827 4472 22869 4481
rect 22827 4432 22828 4472
rect 22868 4432 22869 4472
rect 22827 4423 22869 4432
rect 22731 4304 22773 4313
rect 22731 4264 22732 4304
rect 22772 4264 22773 4304
rect 22731 4255 22773 4264
rect 22251 4220 22293 4229
rect 22251 4180 22252 4220
rect 22292 4180 22293 4220
rect 22251 4171 22293 4180
rect 22444 4220 22484 4229
rect 22635 4220 22677 4229
rect 22484 4180 22580 4220
rect 22444 4171 22484 4180
rect 22252 4086 22292 4171
rect 22348 4136 22388 4145
rect 22348 3641 22388 4096
rect 22540 3893 22580 4180
rect 22635 4180 22636 4220
rect 22676 4180 22677 4220
rect 22635 4171 22677 4180
rect 22636 4086 22676 4171
rect 22732 4170 22772 4255
rect 22828 4220 22868 4423
rect 22828 4171 22868 4180
rect 22923 4220 22965 4229
rect 22923 4180 22924 4220
rect 22964 4180 22965 4220
rect 22923 4171 22965 4180
rect 22539 3884 22581 3893
rect 22539 3844 22540 3884
rect 22580 3844 22581 3884
rect 22539 3835 22581 3844
rect 22443 3800 22485 3809
rect 22443 3760 22444 3800
rect 22484 3760 22485 3800
rect 22443 3751 22485 3760
rect 22347 3632 22389 3641
rect 22156 3592 22292 3632
rect 21964 3473 22004 3558
rect 21963 3464 22005 3473
rect 21963 3424 21964 3464
rect 22004 3424 22005 3464
rect 21963 3415 22005 3424
rect 21868 3256 22004 3296
rect 21772 3212 21812 3221
rect 21812 3172 21908 3212
rect 21772 3163 21812 3172
rect 21676 2500 21812 2540
rect 21483 2491 21525 2500
rect 21579 1616 21621 1625
rect 21579 1576 21580 1616
rect 21620 1576 21621 1616
rect 21579 1567 21621 1576
rect 21388 1324 21524 1364
rect 21292 1240 21428 1280
rect 21388 80 21428 1240
rect 21484 1037 21524 1324
rect 21483 1028 21525 1037
rect 21483 988 21484 1028
rect 21524 988 21525 1028
rect 21483 979 21525 988
rect 21580 80 21620 1567
rect 21772 80 21812 2500
rect 21868 1709 21908 3172
rect 21964 2213 22004 3256
rect 22156 3212 22196 3221
rect 21963 2204 22005 2213
rect 21963 2164 21964 2204
rect 22004 2164 22005 2204
rect 21963 2155 22005 2164
rect 21867 1700 21909 1709
rect 21867 1660 21868 1700
rect 21908 1660 21909 1700
rect 21867 1651 21909 1660
rect 22156 1541 22196 3172
rect 22252 2045 22292 3592
rect 22347 3592 22348 3632
rect 22388 3592 22389 3632
rect 22347 3583 22389 3592
rect 22348 3464 22388 3473
rect 22444 3464 22484 3751
rect 22731 3632 22773 3641
rect 22924 3632 22964 4171
rect 23020 4136 23060 5095
rect 23020 4087 23060 4096
rect 23116 3725 23156 5935
rect 23212 5732 23252 6112
rect 23308 6077 23348 6196
rect 23307 6068 23349 6077
rect 23307 6028 23308 6068
rect 23348 6028 23349 6068
rect 23307 6019 23349 6028
rect 23403 5900 23445 5909
rect 23403 5860 23404 5900
rect 23444 5860 23445 5900
rect 23403 5851 23445 5860
rect 23212 4733 23252 5692
rect 23307 5732 23349 5741
rect 23307 5692 23308 5732
rect 23348 5692 23349 5732
rect 23307 5683 23349 5692
rect 23308 5598 23348 5683
rect 23404 5144 23444 5851
rect 23500 5228 23540 9295
rect 24172 9294 24212 9379
rect 24267 9344 24309 9353
rect 24267 9304 24268 9344
rect 24308 9304 24309 9344
rect 24267 9295 24309 9304
rect 24268 9210 24308 9295
rect 24460 9101 24500 10144
rect 24556 9437 24596 10228
rect 24747 10268 24789 10277
rect 24747 10228 24748 10268
rect 24788 10228 24789 10268
rect 24747 10219 24789 10228
rect 24748 10134 24788 10219
rect 24652 10016 24692 10025
rect 24652 9521 24692 9976
rect 24651 9512 24693 9521
rect 24651 9472 24652 9512
rect 24692 9472 24693 9512
rect 24651 9463 24693 9472
rect 24555 9428 24597 9437
rect 24555 9388 24556 9428
rect 24596 9388 24597 9428
rect 24555 9379 24597 9388
rect 24748 9428 24788 9437
rect 24844 9428 24884 10387
rect 24788 9388 24884 9428
rect 24748 9379 24788 9388
rect 24556 9294 24596 9379
rect 24652 9344 24692 9353
rect 24459 9092 24501 9101
rect 24459 9052 24460 9092
rect 24500 9052 24501 9092
rect 24459 9043 24501 9052
rect 24652 8924 24692 9304
rect 24940 8933 24980 10564
rect 25036 9017 25076 10816
rect 25132 10781 25172 10900
rect 25227 10940 25269 10949
rect 25227 10900 25228 10940
rect 25268 10900 25269 10940
rect 25227 10891 25269 10900
rect 25419 10940 25461 10949
rect 25419 10900 25420 10940
rect 25460 10900 25461 10940
rect 25419 10891 25461 10900
rect 28204 10940 28244 11320
rect 28204 10891 28244 10900
rect 28396 10940 28436 11395
rect 33928 11360 34296 11369
rect 33968 11320 34010 11360
rect 34050 11320 34092 11360
rect 34132 11320 34174 11360
rect 34214 11320 34256 11360
rect 33928 11311 34296 11320
rect 28396 10891 28436 10900
rect 30316 11236 30932 11276
rect 25131 10772 25173 10781
rect 25131 10732 25132 10772
rect 25172 10732 25173 10772
rect 25131 10723 25173 10732
rect 25228 10184 25268 10891
rect 29259 10688 29301 10697
rect 29259 10648 29260 10688
rect 29300 10648 29301 10688
rect 29259 10639 29301 10648
rect 25419 10520 25461 10529
rect 25419 10480 25420 10520
rect 25460 10480 25461 10520
rect 25419 10471 25461 10480
rect 25420 10268 25460 10471
rect 25420 10219 25460 10228
rect 25228 10135 25268 10144
rect 25324 10100 25364 10109
rect 25324 9857 25364 10060
rect 25323 9848 25365 9857
rect 25323 9808 25324 9848
rect 25364 9808 25365 9848
rect 25323 9799 25365 9808
rect 27723 9596 27765 9605
rect 27723 9556 27724 9596
rect 27764 9556 27765 9596
rect 27723 9547 27765 9556
rect 25227 9428 25269 9437
rect 25227 9388 25228 9428
rect 25268 9388 25269 9428
rect 25227 9379 25269 9388
rect 25420 9428 25460 9437
rect 25460 9388 25556 9428
rect 25420 9379 25460 9388
rect 25228 9294 25268 9379
rect 25323 9092 25365 9101
rect 25323 9052 25324 9092
rect 25364 9052 25365 9092
rect 25323 9043 25365 9052
rect 25035 9008 25077 9017
rect 25035 8968 25036 9008
rect 25076 8968 25077 9008
rect 25035 8959 25077 8968
rect 24460 8884 24692 8924
rect 24939 8924 24981 8933
rect 24939 8884 24940 8924
rect 24980 8884 24981 8924
rect 24075 8756 24117 8765
rect 24075 8716 24076 8756
rect 24116 8716 24117 8756
rect 24075 8707 24117 8716
rect 24172 8756 24212 8765
rect 24076 7925 24116 8707
rect 24172 8429 24212 8716
rect 24363 8756 24405 8765
rect 24363 8716 24364 8756
rect 24404 8716 24405 8756
rect 24363 8707 24405 8716
rect 24364 8622 24404 8707
rect 24268 8504 24308 8513
rect 24171 8420 24213 8429
rect 24171 8380 24172 8420
rect 24212 8380 24213 8420
rect 24171 8371 24213 8380
rect 23595 7916 23637 7925
rect 23595 7876 23596 7916
rect 23636 7876 23637 7916
rect 23595 7867 23637 7876
rect 24075 7916 24117 7925
rect 24075 7876 24076 7916
rect 24116 7876 24117 7916
rect 24075 7867 24117 7876
rect 23596 7337 23636 7867
rect 24268 7589 24308 8464
rect 24267 7580 24309 7589
rect 24267 7540 24268 7580
rect 24308 7540 24309 7580
rect 24267 7531 24309 7540
rect 24171 7496 24213 7505
rect 24171 7456 24172 7496
rect 24212 7456 24213 7496
rect 24171 7447 24213 7456
rect 23595 7328 23637 7337
rect 23595 7288 23596 7328
rect 23636 7288 23637 7328
rect 23595 7279 23637 7288
rect 23980 7244 24020 7253
rect 24075 7244 24117 7253
rect 24020 7204 24076 7244
rect 24116 7204 24117 7244
rect 23980 7195 24020 7204
rect 24075 7195 24117 7204
rect 24172 7244 24212 7447
rect 24460 7421 24500 8884
rect 24939 8875 24981 8884
rect 25035 8840 25077 8849
rect 25035 8800 25036 8840
rect 25076 8800 25077 8840
rect 25035 8791 25077 8800
rect 24555 8756 24597 8765
rect 24555 8716 24556 8756
rect 24596 8716 24597 8756
rect 24555 8707 24597 8716
rect 24748 8756 24788 8767
rect 24556 8622 24596 8707
rect 24748 8681 24788 8716
rect 24939 8756 24981 8765
rect 24939 8716 24940 8756
rect 24980 8716 24981 8756
rect 24939 8707 24981 8716
rect 24747 8672 24789 8681
rect 24747 8632 24748 8672
rect 24788 8632 24789 8672
rect 24747 8623 24789 8632
rect 24652 8504 24692 8513
rect 24692 8464 24884 8504
rect 24652 8455 24692 8464
rect 24555 8168 24597 8177
rect 24555 8128 24556 8168
rect 24596 8128 24597 8168
rect 24555 8119 24597 8128
rect 24556 7925 24596 8119
rect 24555 7916 24597 7925
rect 24555 7876 24556 7916
rect 24596 7876 24597 7916
rect 24555 7867 24597 7876
rect 24747 7916 24789 7925
rect 24747 7876 24748 7916
rect 24788 7876 24789 7916
rect 24747 7867 24789 7876
rect 24556 7782 24596 7867
rect 24652 7832 24692 7841
rect 24459 7412 24501 7421
rect 24459 7372 24460 7412
rect 24500 7372 24501 7412
rect 24459 7363 24501 7372
rect 24364 7253 24404 7338
rect 23980 6992 24020 7001
rect 23787 6656 23829 6665
rect 23787 6616 23788 6656
rect 23828 6616 23829 6656
rect 23787 6607 23829 6616
rect 23788 6497 23828 6607
rect 23787 6488 23829 6497
rect 23787 6448 23788 6488
rect 23828 6448 23829 6488
rect 23787 6439 23829 6448
rect 23595 6404 23637 6413
rect 23595 6364 23596 6404
rect 23636 6364 23637 6404
rect 23595 6355 23637 6364
rect 23788 6404 23828 6439
rect 23596 5732 23636 6355
rect 23788 6353 23828 6364
rect 23692 6236 23732 6245
rect 23692 5909 23732 6196
rect 23980 5909 24020 6952
rect 24076 6413 24116 7195
rect 24172 6833 24212 7204
rect 24363 7244 24405 7253
rect 24363 7204 24364 7244
rect 24404 7204 24405 7244
rect 24363 7195 24405 7204
rect 24556 7244 24596 7253
rect 24459 7076 24501 7085
rect 24459 7036 24460 7076
rect 24500 7036 24501 7076
rect 24459 7027 24501 7036
rect 24363 6992 24405 7001
rect 24363 6952 24364 6992
rect 24404 6952 24405 6992
rect 24363 6943 24405 6952
rect 24267 6908 24309 6917
rect 24267 6868 24268 6908
rect 24308 6868 24309 6908
rect 24267 6859 24309 6868
rect 24171 6824 24213 6833
rect 24171 6784 24172 6824
rect 24212 6784 24213 6824
rect 24171 6775 24213 6784
rect 24268 6572 24308 6859
rect 24364 6858 24404 6943
rect 24268 6532 24404 6572
rect 24075 6404 24117 6413
rect 24075 6364 24076 6404
rect 24116 6364 24117 6404
rect 24075 6355 24117 6364
rect 24268 6404 24308 6413
rect 23691 5900 23733 5909
rect 23691 5860 23692 5900
rect 23732 5860 23733 5900
rect 23691 5851 23733 5860
rect 23979 5900 24021 5909
rect 23979 5860 23980 5900
rect 24020 5860 24021 5900
rect 23979 5851 24021 5860
rect 23788 5732 23828 5741
rect 23596 5692 23788 5732
rect 23788 5683 23828 5692
rect 23979 5732 24021 5741
rect 23979 5692 23980 5732
rect 24020 5692 24021 5732
rect 24076 5732 24116 6355
rect 24268 6245 24308 6364
rect 24267 6236 24309 6245
rect 24267 6196 24268 6236
rect 24308 6196 24309 6236
rect 24267 6187 24309 6196
rect 24172 5732 24212 5741
rect 24076 5692 24172 5732
rect 23979 5683 24021 5692
rect 24172 5683 24212 5692
rect 24364 5732 24404 6532
rect 24460 6404 24500 7027
rect 24556 6749 24596 7204
rect 24555 6740 24597 6749
rect 24555 6700 24556 6740
rect 24596 6700 24597 6740
rect 24555 6691 24597 6700
rect 24652 6572 24692 7792
rect 24748 7782 24788 7867
rect 24747 7328 24789 7337
rect 24747 7288 24748 7328
rect 24788 7288 24789 7328
rect 24747 7279 24789 7288
rect 24748 7001 24788 7279
rect 24747 6992 24789 7001
rect 24747 6952 24748 6992
rect 24788 6952 24789 6992
rect 24747 6943 24789 6952
rect 24460 6355 24500 6364
rect 24556 6532 24692 6572
rect 24459 6236 24501 6245
rect 24459 6196 24460 6236
rect 24500 6196 24501 6236
rect 24459 6187 24501 6196
rect 24460 6102 24500 6187
rect 24364 5683 24404 5692
rect 23980 5598 24020 5683
rect 23787 5480 23829 5489
rect 24172 5480 24212 5489
rect 23787 5440 23788 5480
rect 23828 5440 23829 5480
rect 23787 5431 23829 5440
rect 23980 5440 24172 5480
rect 23788 5346 23828 5431
rect 23500 5188 23828 5228
rect 23308 5104 23444 5144
rect 23788 5144 23828 5188
rect 23788 5104 23833 5144
rect 23211 4724 23253 4733
rect 23211 4684 23212 4724
rect 23252 4684 23253 4724
rect 23211 4675 23253 4684
rect 23212 3968 23252 3977
rect 23115 3716 23157 3725
rect 23115 3676 23116 3716
rect 23156 3676 23157 3716
rect 23115 3667 23157 3676
rect 22731 3592 22732 3632
rect 22772 3592 22773 3632
rect 22731 3583 22773 3592
rect 22828 3592 22964 3632
rect 22635 3548 22677 3557
rect 22635 3508 22636 3548
rect 22676 3508 22677 3548
rect 22635 3499 22677 3508
rect 22388 3424 22484 3464
rect 22348 3415 22388 3424
rect 22540 3212 22580 3221
rect 22251 2036 22293 2045
rect 22251 1996 22252 2036
rect 22292 1996 22293 2036
rect 22251 1987 22293 1996
rect 21963 1532 22005 1541
rect 21963 1492 21964 1532
rect 22004 1492 22005 1532
rect 21963 1483 22005 1492
rect 22155 1532 22197 1541
rect 22155 1492 22156 1532
rect 22196 1492 22197 1532
rect 22155 1483 22197 1492
rect 21964 80 22004 1483
rect 22347 1364 22389 1373
rect 22347 1324 22348 1364
rect 22388 1324 22389 1364
rect 22347 1315 22389 1324
rect 22155 1196 22197 1205
rect 22155 1156 22156 1196
rect 22196 1156 22197 1196
rect 22155 1147 22197 1156
rect 22156 80 22196 1147
rect 22348 80 22388 1315
rect 22540 1121 22580 3172
rect 22636 2372 22676 3499
rect 22732 3464 22772 3583
rect 22732 3415 22772 3424
rect 22636 2332 22772 2372
rect 22539 1112 22581 1121
rect 22539 1072 22540 1112
rect 22580 1072 22581 1112
rect 22539 1063 22581 1072
rect 22539 944 22581 953
rect 22539 904 22540 944
rect 22580 904 22581 944
rect 22539 895 22581 904
rect 22540 80 22580 895
rect 22732 80 22772 2332
rect 22828 785 22868 3592
rect 23116 3473 23156 3558
rect 23115 3464 23157 3473
rect 23115 3424 23116 3464
rect 23156 3424 23157 3464
rect 23115 3415 23157 3424
rect 22924 3212 22964 3221
rect 22924 1793 22964 3172
rect 23115 3212 23157 3221
rect 23115 3172 23116 3212
rect 23156 3172 23157 3212
rect 23115 3163 23157 3172
rect 23019 1868 23061 1877
rect 23019 1828 23020 1868
rect 23060 1828 23061 1868
rect 23019 1819 23061 1828
rect 22923 1784 22965 1793
rect 22923 1744 22924 1784
rect 22964 1744 22965 1784
rect 22923 1735 22965 1744
rect 23020 1196 23060 1819
rect 23116 1280 23156 3163
rect 23212 1364 23252 3928
rect 23308 3389 23348 5104
rect 23595 5060 23637 5069
rect 23595 5020 23596 5060
rect 23636 5020 23637 5060
rect 23595 5011 23637 5020
rect 23404 4892 23444 4903
rect 23404 4817 23444 4852
rect 23596 4892 23636 5011
rect 23793 4976 23833 5104
rect 23788 4963 23833 4976
rect 23828 4936 23833 4963
rect 23788 4914 23828 4923
rect 23980 4892 24020 5440
rect 24172 5431 24212 5440
rect 24363 5228 24405 5237
rect 24363 5188 24364 5228
rect 24404 5188 24405 5228
rect 24363 5179 24405 5188
rect 23596 4843 23636 4852
rect 23884 4852 24020 4892
rect 24171 4892 24213 4901
rect 24171 4852 24172 4892
rect 24212 4852 24213 4892
rect 23403 4808 23445 4817
rect 23403 4768 23404 4808
rect 23444 4768 23445 4808
rect 23403 4759 23445 4768
rect 23787 4808 23829 4817
rect 23787 4768 23788 4808
rect 23828 4768 23829 4808
rect 23787 4759 23829 4768
rect 23500 4724 23540 4733
rect 23500 4640 23540 4684
rect 23500 4600 23636 4640
rect 23403 4304 23445 4313
rect 23403 4264 23404 4304
rect 23444 4264 23445 4304
rect 23403 4255 23445 4264
rect 23404 4136 23444 4255
rect 23596 4229 23636 4600
rect 23788 4388 23828 4759
rect 23692 4348 23828 4388
rect 23595 4220 23637 4229
rect 23595 4180 23596 4220
rect 23636 4180 23637 4220
rect 23595 4171 23637 4180
rect 23404 4087 23444 4096
rect 23596 3968 23636 3977
rect 23499 3464 23541 3473
rect 23499 3424 23500 3464
rect 23540 3424 23541 3464
rect 23499 3415 23541 3424
rect 23307 3380 23349 3389
rect 23307 3340 23308 3380
rect 23348 3340 23349 3380
rect 23307 3331 23349 3340
rect 23500 3330 23540 3415
rect 23308 3212 23348 3221
rect 23308 1625 23348 3172
rect 23596 2540 23636 3928
rect 23692 3464 23732 4348
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23829 4220
rect 23787 4171 23829 4180
rect 23788 4086 23828 4171
rect 23884 3641 23924 4852
rect 24171 4843 24213 4852
rect 24364 4892 24404 5179
rect 24556 5060 24596 6532
rect 24748 6488 24788 6943
rect 24652 6448 24788 6488
rect 24652 6446 24692 6448
rect 24652 6397 24692 6406
rect 24748 6390 24788 6399
rect 24748 6320 24788 6350
rect 24652 6280 24788 6320
rect 24652 6161 24692 6280
rect 24651 6152 24693 6161
rect 24651 6112 24652 6152
rect 24692 6112 24693 6152
rect 24651 6103 24693 6112
rect 24747 6068 24789 6077
rect 24747 6028 24748 6068
rect 24788 6028 24789 6068
rect 24747 6019 24789 6028
rect 24748 5732 24788 6019
rect 24748 5683 24788 5692
rect 24364 4843 24404 4852
rect 24460 5020 24596 5060
rect 23980 4724 24020 4733
rect 24020 4684 24116 4724
rect 23980 4675 24020 4684
rect 23980 4229 24020 4314
rect 23979 4220 24021 4229
rect 23979 4180 23980 4220
rect 24020 4180 24021 4220
rect 23979 4171 24021 4180
rect 23979 4052 24021 4061
rect 23979 4012 23980 4052
rect 24020 4012 24021 4052
rect 23979 4003 24021 4012
rect 23980 3918 24020 4003
rect 23883 3632 23925 3641
rect 23883 3592 23884 3632
rect 23924 3592 23925 3632
rect 23883 3583 23925 3592
rect 23884 3464 23924 3473
rect 23692 3424 23884 3464
rect 23884 3415 23924 3424
rect 24076 3380 24116 4684
rect 24172 4229 24212 4843
rect 24268 4724 24308 4733
rect 24268 4397 24308 4684
rect 24363 4640 24405 4649
rect 24363 4600 24364 4640
rect 24404 4600 24405 4640
rect 24363 4591 24405 4600
rect 24267 4388 24309 4397
rect 24267 4348 24268 4388
rect 24308 4348 24309 4388
rect 24267 4339 24309 4348
rect 24171 4220 24213 4229
rect 24171 4180 24172 4220
rect 24212 4180 24213 4220
rect 24171 4171 24213 4180
rect 24364 4220 24404 4591
rect 24364 4171 24404 4180
rect 24172 4086 24212 4171
rect 24267 4136 24309 4145
rect 24267 4096 24268 4136
rect 24308 4096 24309 4136
rect 24267 4087 24309 4096
rect 24268 4002 24308 4087
rect 24268 3464 24308 3473
rect 24460 3464 24500 5020
rect 24651 4976 24693 4985
rect 24651 4936 24652 4976
rect 24692 4936 24693 4976
rect 24651 4927 24693 4936
rect 24555 4892 24597 4901
rect 24555 4852 24556 4892
rect 24596 4852 24597 4892
rect 24555 4843 24597 4852
rect 24556 4220 24596 4843
rect 24652 4842 24692 4927
rect 24748 4892 24788 4901
rect 24748 4724 24788 4852
rect 24652 4684 24788 4724
rect 24652 4397 24692 4684
rect 24747 4556 24789 4565
rect 24747 4516 24748 4556
rect 24788 4516 24789 4556
rect 24747 4507 24789 4516
rect 24651 4388 24693 4397
rect 24651 4348 24652 4388
rect 24692 4348 24693 4388
rect 24651 4339 24693 4348
rect 24556 4171 24596 4180
rect 24748 4220 24788 4507
rect 24748 4171 24788 4180
rect 24555 3968 24597 3977
rect 24555 3928 24556 3968
rect 24596 3928 24597 3968
rect 24555 3919 24597 3928
rect 24556 3834 24596 3919
rect 24651 3800 24693 3809
rect 24651 3760 24652 3800
rect 24692 3760 24693 3800
rect 24651 3751 24693 3760
rect 24308 3424 24500 3464
rect 24652 3464 24692 3751
rect 24844 3464 24884 8464
rect 24940 7925 24980 8707
rect 25036 8706 25076 8791
rect 25132 8756 25172 8765
rect 25132 8261 25172 8716
rect 25324 8345 25364 9043
rect 25419 8756 25461 8765
rect 25419 8716 25420 8756
rect 25460 8716 25461 8756
rect 25516 8756 25556 9388
rect 26859 8840 26901 8849
rect 26859 8800 26860 8840
rect 26900 8800 26901 8840
rect 26859 8791 26901 8800
rect 25612 8756 25652 8765
rect 25516 8716 25612 8756
rect 25419 8707 25461 8716
rect 25420 8622 25460 8707
rect 25612 8513 25652 8716
rect 25611 8504 25653 8513
rect 25611 8464 25612 8504
rect 25652 8464 25653 8504
rect 25611 8455 25653 8464
rect 25323 8336 25365 8345
rect 25323 8296 25324 8336
rect 25364 8296 25365 8336
rect 25323 8287 25365 8296
rect 25131 8252 25173 8261
rect 25131 8212 25132 8252
rect 25172 8212 25173 8252
rect 25131 8203 25173 8212
rect 25131 8000 25173 8009
rect 25131 7960 25132 8000
rect 25172 7960 25173 8000
rect 25131 7951 25173 7960
rect 24939 7916 24981 7925
rect 24939 7876 24940 7916
rect 24980 7876 24981 7916
rect 24939 7867 24981 7876
rect 25132 7916 25172 7951
rect 24940 7244 24980 7867
rect 25132 7865 25172 7876
rect 25324 7916 25364 8287
rect 25899 8084 25941 8093
rect 25899 8044 25900 8084
rect 25940 8044 25941 8084
rect 25899 8035 25941 8044
rect 25324 7867 25364 7876
rect 25515 7916 25557 7925
rect 25515 7876 25516 7916
rect 25556 7876 25557 7916
rect 25515 7867 25557 7876
rect 25707 7916 25749 7925
rect 25707 7876 25708 7916
rect 25748 7876 25749 7916
rect 25707 7867 25749 7876
rect 25900 7916 25940 8035
rect 25900 7867 25940 7876
rect 25035 7832 25077 7841
rect 25035 7792 25036 7832
rect 25076 7792 25077 7832
rect 25035 7783 25077 7792
rect 25420 7832 25460 7841
rect 25036 7698 25076 7783
rect 25227 7748 25269 7757
rect 25227 7708 25228 7748
rect 25268 7708 25269 7748
rect 25227 7699 25269 7708
rect 25036 7244 25076 7253
rect 24940 7204 25036 7244
rect 25036 7195 25076 7204
rect 25131 7244 25173 7253
rect 25131 7204 25132 7244
rect 25172 7204 25173 7244
rect 25131 7195 25173 7204
rect 25228 7244 25268 7699
rect 25228 7195 25268 7204
rect 25132 7110 25172 7195
rect 25035 7076 25077 7085
rect 25035 7036 25036 7076
rect 25076 7036 25077 7076
rect 25035 7027 25077 7036
rect 25036 6749 25076 7027
rect 25035 6740 25077 6749
rect 25035 6700 25036 6740
rect 25076 6700 25077 6740
rect 25035 6691 25077 6700
rect 25131 6656 25173 6665
rect 25131 6616 25132 6656
rect 25172 6616 25173 6656
rect 25131 6607 25173 6616
rect 24950 6405 24990 6414
rect 25035 6404 25077 6413
rect 24990 6365 25036 6404
rect 24950 6364 25036 6365
rect 25076 6364 25077 6404
rect 24950 6356 24990 6364
rect 25035 6355 25077 6364
rect 25132 6404 25172 6607
rect 25420 6572 25460 7792
rect 25516 7782 25556 7867
rect 25708 7782 25748 7867
rect 25804 7832 25844 7841
rect 25707 7580 25749 7589
rect 25707 7540 25708 7580
rect 25748 7540 25749 7580
rect 25707 7531 25749 7540
rect 25132 6355 25172 6364
rect 25228 6532 25460 6572
rect 25036 6236 25076 6245
rect 24940 5732 24980 5741
rect 24940 4901 24980 5692
rect 25036 5405 25076 6196
rect 25035 5396 25077 5405
rect 25035 5356 25036 5396
rect 25076 5356 25077 5396
rect 25035 5347 25077 5356
rect 25131 5228 25173 5237
rect 25131 5188 25132 5228
rect 25172 5188 25173 5228
rect 25131 5179 25173 5188
rect 25132 5069 25172 5179
rect 25131 5060 25173 5069
rect 25131 5020 25132 5060
rect 25172 5020 25173 5060
rect 25131 5011 25173 5020
rect 24939 4892 24981 4901
rect 24939 4852 24940 4892
rect 24980 4852 24981 4892
rect 24939 4843 24981 4852
rect 25132 4892 25172 5011
rect 25132 4843 25172 4852
rect 24940 4220 24980 4843
rect 25228 4817 25268 6532
rect 25323 6404 25365 6413
rect 25323 6364 25324 6404
rect 25364 6364 25365 6404
rect 25323 6355 25365 6364
rect 25515 6404 25557 6413
rect 25515 6364 25516 6404
rect 25556 6364 25557 6404
rect 25515 6355 25557 6364
rect 25324 6270 25364 6355
rect 25516 6270 25556 6355
rect 25420 6236 25460 6245
rect 25420 5153 25460 6196
rect 25708 5984 25748 7531
rect 25804 6404 25844 7792
rect 26475 7832 26517 7841
rect 26475 7792 26476 7832
rect 26516 7792 26517 7832
rect 26475 7783 26517 7792
rect 26380 6413 26420 6498
rect 26187 6404 26229 6413
rect 25804 6364 26132 6404
rect 25708 5944 25844 5984
rect 25419 5144 25461 5153
rect 25419 5104 25420 5144
rect 25460 5104 25461 5144
rect 25419 5095 25461 5104
rect 25324 4901 25364 4986
rect 25323 4892 25365 4901
rect 25323 4852 25324 4892
rect 25364 4852 25365 4892
rect 25323 4843 25365 4852
rect 25516 4892 25556 4901
rect 25516 4817 25556 4852
rect 25227 4808 25269 4817
rect 25227 4768 25228 4808
rect 25268 4768 25269 4808
rect 25227 4759 25269 4768
rect 25515 4808 25557 4817
rect 25515 4768 25516 4808
rect 25556 4768 25557 4808
rect 25515 4759 25557 4768
rect 25035 4724 25077 4733
rect 25035 4684 25036 4724
rect 25076 4684 25077 4724
rect 25035 4675 25077 4684
rect 25323 4724 25365 4733
rect 25323 4684 25324 4724
rect 25364 4684 25365 4724
rect 25323 4675 25365 4684
rect 25420 4724 25460 4733
rect 25036 4590 25076 4675
rect 24940 4171 24980 4180
rect 25132 4220 25172 4229
rect 25036 4136 25076 4145
rect 25036 3632 25076 4096
rect 25132 3893 25172 4180
rect 25324 4136 25364 4675
rect 25324 4087 25364 4096
rect 25131 3884 25173 3893
rect 25131 3844 25132 3884
rect 25172 3844 25173 3884
rect 25131 3835 25173 3844
rect 25420 3641 25460 4684
rect 25516 4313 25556 4759
rect 25708 4724 25748 4733
rect 25515 4304 25557 4313
rect 25515 4264 25516 4304
rect 25556 4264 25557 4304
rect 25515 4255 25557 4264
rect 25708 4231 25748 4684
rect 25612 4191 25748 4231
rect 25804 4219 25844 5944
rect 25899 5060 25941 5069
rect 25899 5020 25900 5060
rect 25940 5020 25941 5060
rect 25899 5011 25941 5020
rect 25900 4976 25940 5011
rect 25900 4925 25940 4936
rect 26092 4976 26132 6364
rect 26187 6364 26188 6404
rect 26228 6364 26229 6404
rect 26187 6355 26229 6364
rect 26379 6404 26421 6413
rect 26379 6364 26380 6404
rect 26420 6364 26421 6404
rect 26379 6355 26421 6364
rect 26188 5993 26228 6355
rect 26284 6236 26324 6245
rect 26187 5984 26229 5993
rect 26187 5944 26188 5984
rect 26228 5944 26229 5984
rect 26187 5935 26229 5944
rect 26092 4927 26132 4936
rect 26284 4892 26324 6196
rect 26379 6236 26421 6245
rect 26379 6196 26380 6236
rect 26420 6196 26421 6236
rect 26379 6187 26421 6196
rect 26188 4852 26324 4892
rect 26188 4808 26228 4852
rect 25996 4768 26228 4808
rect 25516 3968 25556 3977
rect 25419 3632 25461 3641
rect 25036 3592 25172 3632
rect 25036 3464 25076 3473
rect 24844 3424 25036 3464
rect 24268 3415 24308 3424
rect 24652 3415 24692 3424
rect 25036 3415 25076 3424
rect 24076 3340 24212 3380
rect 23692 3212 23732 3221
rect 23692 2549 23732 3172
rect 24076 3212 24116 3221
rect 23500 2500 23636 2540
rect 23691 2540 23733 2549
rect 23691 2500 23692 2540
rect 23732 2500 23733 2540
rect 23307 1616 23349 1625
rect 23307 1576 23308 1616
rect 23348 1576 23349 1616
rect 23307 1567 23349 1576
rect 23212 1324 23444 1364
rect 23116 1240 23348 1280
rect 23020 1156 23156 1196
rect 22923 860 22965 869
rect 22923 820 22924 860
rect 22964 820 22965 860
rect 22923 811 22965 820
rect 22827 776 22869 785
rect 22827 736 22828 776
rect 22868 736 22869 776
rect 22827 727 22869 736
rect 22924 80 22964 811
rect 23116 80 23156 1156
rect 23308 80 23348 1240
rect 23404 1205 23444 1324
rect 23500 1289 23540 2500
rect 23691 2491 23733 2500
rect 23691 1700 23733 1709
rect 23691 1660 23692 1700
rect 23732 1660 23733 1700
rect 23691 1651 23733 1660
rect 23499 1280 23541 1289
rect 23499 1240 23500 1280
rect 23540 1240 23541 1280
rect 23499 1231 23541 1240
rect 23403 1196 23445 1205
rect 23403 1156 23404 1196
rect 23444 1156 23445 1196
rect 23403 1147 23445 1156
rect 23499 1028 23541 1037
rect 23499 988 23500 1028
rect 23540 988 23541 1028
rect 23499 979 23541 988
rect 23500 80 23540 979
rect 23692 80 23732 1651
rect 23883 1532 23925 1541
rect 23883 1492 23884 1532
rect 23924 1492 23925 1532
rect 23883 1483 23925 1492
rect 23884 80 23924 1483
rect 24076 1373 24116 3172
rect 24172 2540 24212 3340
rect 24460 3212 24500 3221
rect 24172 2500 24308 2540
rect 24075 1364 24117 1373
rect 24075 1324 24076 1364
rect 24116 1324 24117 1364
rect 24075 1315 24117 1324
rect 24075 1196 24117 1205
rect 24075 1156 24076 1196
rect 24116 1156 24117 1196
rect 24075 1147 24117 1156
rect 24076 80 24116 1147
rect 24268 80 24308 2500
rect 24460 1541 24500 3172
rect 24844 3212 24884 3221
rect 24747 1784 24789 1793
rect 24747 1744 24748 1784
rect 24788 1744 24789 1784
rect 24747 1735 24789 1744
rect 24459 1532 24501 1541
rect 24459 1492 24460 1532
rect 24500 1492 24501 1532
rect 24459 1483 24501 1492
rect 24651 1280 24693 1289
rect 24651 1240 24652 1280
rect 24692 1240 24693 1280
rect 24748 1280 24788 1735
rect 24844 1709 24884 3172
rect 25132 2297 25172 3592
rect 25419 3592 25420 3632
rect 25460 3592 25461 3632
rect 25419 3583 25461 3592
rect 25419 3464 25461 3473
rect 25419 3424 25420 3464
rect 25460 3424 25461 3464
rect 25419 3415 25461 3424
rect 25420 3330 25460 3415
rect 25227 3212 25269 3221
rect 25227 3172 25228 3212
rect 25268 3172 25269 3212
rect 25227 3163 25269 3172
rect 25228 3078 25268 3163
rect 25227 2456 25269 2465
rect 25227 2416 25228 2456
rect 25268 2416 25269 2456
rect 25227 2407 25269 2416
rect 25131 2288 25173 2297
rect 25131 2248 25132 2288
rect 25172 2248 25173 2288
rect 25131 2239 25173 2248
rect 24843 1700 24885 1709
rect 24843 1660 24844 1700
rect 24884 1660 24885 1700
rect 24843 1651 24885 1660
rect 25035 1616 25077 1625
rect 25035 1576 25036 1616
rect 25076 1576 25077 1616
rect 25035 1567 25077 1576
rect 24748 1240 24884 1280
rect 24651 1231 24693 1240
rect 24459 1112 24501 1121
rect 24459 1072 24460 1112
rect 24500 1072 24501 1112
rect 24459 1063 24501 1072
rect 24460 80 24500 1063
rect 24652 80 24692 1231
rect 24844 80 24884 1240
rect 25036 80 25076 1567
rect 25228 80 25268 2407
rect 25419 1364 25461 1373
rect 25419 1324 25420 1364
rect 25460 1324 25461 1364
rect 25419 1315 25461 1324
rect 25420 80 25460 1315
rect 25516 1289 25556 3928
rect 25612 3380 25652 4191
rect 25804 4179 25855 4219
rect 25707 4136 25749 4145
rect 25707 4096 25708 4136
rect 25748 4096 25749 4136
rect 25707 4087 25749 4096
rect 25708 4002 25748 4087
rect 25815 4052 25855 4179
rect 25804 4012 25855 4052
rect 25804 3464 25844 4012
rect 25804 3415 25844 3424
rect 25900 3968 25940 3977
rect 25612 3340 25748 3380
rect 25612 3212 25652 3221
rect 25612 2549 25652 3172
rect 25611 2540 25653 2549
rect 25611 2500 25612 2540
rect 25652 2500 25653 2540
rect 25611 2491 25653 2500
rect 25708 2372 25748 3340
rect 25612 2332 25748 2372
rect 25515 1280 25557 1289
rect 25515 1240 25516 1280
rect 25556 1240 25557 1280
rect 25515 1231 25557 1240
rect 25612 80 25652 2332
rect 25803 1532 25845 1541
rect 25803 1492 25804 1532
rect 25844 1492 25845 1532
rect 25803 1483 25845 1492
rect 25804 80 25844 1483
rect 25900 1205 25940 3928
rect 25996 3389 26036 4768
rect 26284 4724 26324 4733
rect 26188 4684 26284 4724
rect 26092 4136 26132 4147
rect 26092 4061 26132 4096
rect 26091 4052 26133 4061
rect 26091 4012 26092 4052
rect 26132 4012 26133 4052
rect 26091 4003 26133 4012
rect 26188 3632 26228 4684
rect 26284 4675 26324 4684
rect 26092 3592 26228 3632
rect 26284 3968 26324 3977
rect 25995 3380 26037 3389
rect 25995 3340 25996 3380
rect 26036 3340 26037 3380
rect 25995 3331 26037 3340
rect 25996 3212 26036 3221
rect 25996 1793 26036 3172
rect 26092 2540 26132 3592
rect 26188 3464 26228 3475
rect 26188 3389 26228 3424
rect 26187 3380 26229 3389
rect 26187 3340 26188 3380
rect 26228 3340 26229 3380
rect 26187 3331 26229 3340
rect 26092 2500 26228 2540
rect 25995 1784 26037 1793
rect 25995 1744 25996 1784
rect 26036 1744 26037 1784
rect 25995 1735 26037 1744
rect 25995 1280 26037 1289
rect 25995 1240 25996 1280
rect 26036 1240 26037 1280
rect 25995 1231 26037 1240
rect 25899 1196 25941 1205
rect 25899 1156 25900 1196
rect 25940 1156 25941 1196
rect 25899 1147 25941 1156
rect 25996 80 26036 1231
rect 26188 80 26228 2500
rect 26284 1037 26324 3928
rect 26380 3389 26420 6187
rect 26476 5144 26516 7783
rect 26571 6488 26613 6497
rect 26571 6448 26572 6488
rect 26612 6448 26613 6488
rect 26571 6439 26613 6448
rect 26572 6404 26612 6439
rect 26572 6353 26612 6364
rect 26763 6404 26805 6413
rect 26763 6364 26764 6404
rect 26804 6364 26805 6404
rect 26763 6355 26805 6364
rect 26571 6236 26613 6245
rect 26571 6196 26572 6236
rect 26612 6196 26613 6236
rect 26571 6187 26613 6196
rect 26668 6236 26708 6245
rect 26572 5909 26612 6187
rect 26571 5900 26613 5909
rect 26571 5860 26572 5900
rect 26612 5860 26613 5900
rect 26571 5851 26613 5860
rect 26572 5732 26612 5851
rect 26572 5683 26612 5692
rect 26476 5104 26612 5144
rect 26476 4976 26516 4985
rect 26476 4817 26516 4936
rect 26475 4808 26517 4817
rect 26475 4768 26476 4808
rect 26516 4768 26517 4808
rect 26475 4759 26517 4768
rect 26476 4136 26516 4145
rect 26572 4136 26612 5104
rect 26668 4901 26708 6196
rect 26764 5732 26804 6355
rect 26764 5683 26804 5692
rect 26764 5480 26804 5489
rect 26667 4892 26709 4901
rect 26667 4852 26668 4892
rect 26708 4852 26709 4892
rect 26667 4843 26709 4852
rect 26764 4808 26804 5440
rect 26860 4976 26900 8791
rect 27436 8756 27476 8765
rect 27436 8429 27476 8716
rect 27627 8756 27669 8765
rect 27627 8716 27628 8756
rect 27668 8716 27669 8756
rect 27627 8707 27669 8716
rect 27532 8504 27572 8513
rect 27435 8420 27477 8429
rect 27435 8380 27436 8420
rect 27476 8380 27477 8420
rect 27435 8371 27477 8380
rect 26956 7253 26996 7338
rect 26955 7244 26997 7253
rect 27148 7244 27188 7253
rect 26955 7204 26956 7244
rect 26996 7204 26997 7244
rect 26955 7195 26997 7204
rect 27052 7204 27148 7244
rect 27052 7076 27092 7204
rect 27148 7195 27188 7204
rect 26956 7036 27092 7076
rect 26956 6413 26996 7036
rect 27148 6992 27188 7001
rect 27188 6952 27284 6992
rect 27148 6943 27188 6952
rect 27147 6656 27189 6665
rect 27147 6616 27148 6656
rect 27188 6616 27189 6656
rect 27147 6607 27189 6616
rect 26955 6404 26997 6413
rect 26955 6364 26956 6404
rect 26996 6364 26997 6404
rect 26955 6355 26997 6364
rect 27148 6404 27188 6607
rect 27148 6355 27188 6364
rect 26956 6068 26996 6355
rect 27051 6320 27093 6329
rect 27051 6280 27052 6320
rect 27092 6280 27093 6320
rect 27051 6271 27093 6280
rect 27052 6186 27092 6271
rect 26956 6028 27188 6068
rect 26955 5900 26997 5909
rect 26955 5860 26956 5900
rect 26996 5860 26997 5900
rect 26955 5851 26997 5860
rect 26956 5732 26996 5851
rect 26956 5683 26996 5692
rect 27148 5732 27188 6028
rect 27148 5683 27188 5692
rect 27244 5648 27284 6952
rect 27339 6908 27381 6917
rect 27339 6868 27340 6908
rect 27380 6868 27381 6908
rect 27339 6859 27381 6868
rect 27340 6404 27380 6859
rect 27532 6572 27572 8464
rect 27628 7925 27668 8707
rect 27724 8084 27764 9547
rect 28107 9344 28149 9353
rect 28107 9304 28108 9344
rect 28148 9304 28149 9344
rect 28107 9295 28149 9304
rect 27915 8840 27957 8849
rect 27915 8800 27916 8840
rect 27956 8800 27957 8840
rect 27915 8791 27957 8800
rect 27819 8756 27861 8765
rect 27819 8716 27820 8756
rect 27860 8716 27861 8756
rect 27819 8707 27861 8716
rect 27820 8622 27860 8707
rect 27916 8706 27956 8791
rect 28012 8756 28052 8765
rect 28012 8261 28052 8716
rect 28108 8597 28148 9295
rect 28683 9176 28725 9185
rect 28683 9136 28684 9176
rect 28724 9136 28725 9176
rect 28683 9127 28725 9136
rect 28299 8924 28341 8933
rect 28299 8884 28300 8924
rect 28340 8884 28341 8924
rect 28299 8875 28341 8884
rect 28300 8840 28340 8875
rect 28300 8789 28340 8800
rect 28684 8840 28724 9127
rect 28684 8791 28724 8800
rect 28203 8756 28245 8765
rect 28203 8716 28204 8756
rect 28244 8716 28245 8756
rect 28203 8707 28245 8716
rect 28396 8756 28436 8767
rect 28204 8622 28244 8707
rect 28396 8681 28436 8716
rect 28587 8756 28629 8765
rect 28587 8716 28588 8756
rect 28628 8716 28629 8756
rect 28587 8707 28629 8716
rect 28780 8756 28820 8765
rect 28820 8716 28916 8756
rect 28780 8707 28820 8716
rect 28395 8672 28437 8681
rect 28395 8632 28396 8672
rect 28436 8632 28437 8672
rect 28395 8623 28437 8632
rect 28588 8622 28628 8707
rect 28683 8672 28725 8681
rect 28683 8632 28684 8672
rect 28724 8632 28725 8672
rect 28683 8623 28725 8632
rect 28107 8588 28149 8597
rect 28107 8548 28108 8588
rect 28148 8548 28149 8588
rect 28107 8539 28149 8548
rect 28587 8336 28629 8345
rect 28587 8296 28588 8336
rect 28628 8296 28629 8336
rect 28587 8287 28629 8296
rect 28011 8252 28053 8261
rect 28011 8212 28012 8252
rect 28052 8212 28053 8252
rect 28011 8203 28053 8212
rect 28203 8168 28245 8177
rect 28203 8128 28204 8168
rect 28244 8128 28245 8168
rect 28203 8119 28245 8128
rect 27724 8044 27956 8084
rect 27627 7916 27669 7925
rect 27627 7876 27628 7916
rect 27668 7876 27669 7916
rect 27627 7867 27669 7876
rect 27820 7916 27860 7925
rect 27628 7782 27668 7867
rect 27724 7832 27764 7841
rect 27724 6656 27764 7792
rect 27820 7757 27860 7876
rect 27819 7748 27861 7757
rect 27819 7708 27820 7748
rect 27860 7708 27861 7748
rect 27819 7699 27861 7708
rect 27916 6833 27956 8044
rect 28011 7916 28053 7925
rect 28011 7876 28012 7916
rect 28052 7876 28053 7916
rect 28011 7867 28053 7876
rect 28204 7916 28244 8119
rect 28012 7782 28052 7867
rect 28108 7832 28148 7841
rect 27915 6824 27957 6833
rect 27915 6784 27916 6824
rect 27956 6784 27957 6824
rect 27915 6775 27957 6784
rect 27724 6616 28052 6656
rect 27532 6532 27668 6572
rect 27340 6355 27380 6364
rect 27531 6404 27573 6413
rect 27531 6364 27532 6404
rect 27572 6364 27573 6404
rect 27531 6355 27573 6364
rect 27435 6320 27477 6329
rect 27435 6280 27436 6320
rect 27476 6280 27477 6320
rect 27435 6271 27477 6280
rect 27436 6186 27476 6271
rect 27532 6270 27572 6355
rect 27628 5657 27668 6532
rect 27916 6497 27956 6512
rect 27915 6488 27957 6497
rect 27915 6448 27916 6488
rect 27956 6448 27957 6488
rect 27915 6439 27957 6448
rect 27916 6417 27956 6439
rect 27724 6404 27764 6413
rect 27916 6368 27956 6377
rect 27724 6077 27764 6364
rect 27820 6320 27860 6329
rect 27723 6068 27765 6077
rect 27723 6028 27724 6068
rect 27764 6028 27765 6068
rect 27723 6019 27765 6028
rect 27724 5741 27764 6019
rect 27723 5732 27765 5741
rect 27723 5692 27724 5732
rect 27764 5692 27765 5732
rect 27723 5683 27765 5692
rect 27627 5648 27669 5657
rect 27244 5608 27380 5648
rect 27148 5480 27188 5489
rect 27148 5153 27188 5440
rect 27243 5480 27285 5489
rect 27243 5440 27244 5480
rect 27284 5440 27285 5480
rect 27243 5431 27285 5440
rect 27147 5144 27189 5153
rect 27147 5104 27148 5144
rect 27188 5104 27189 5144
rect 27147 5095 27189 5104
rect 26860 4927 26900 4936
rect 27244 4976 27284 5431
rect 27244 4927 27284 4936
rect 26955 4892 26997 4901
rect 26955 4852 26956 4892
rect 26996 4852 26997 4892
rect 26955 4843 26997 4852
rect 26764 4768 26900 4808
rect 26668 4724 26708 4733
rect 26708 4684 26804 4724
rect 26668 4675 26708 4684
rect 26516 4096 26612 4136
rect 26476 4087 26516 4096
rect 26668 3968 26708 3977
rect 26571 3632 26613 3641
rect 26571 3592 26572 3632
rect 26612 3592 26613 3632
rect 26571 3583 26613 3592
rect 26572 3464 26612 3583
rect 26668 3557 26708 3928
rect 26667 3548 26709 3557
rect 26667 3508 26668 3548
rect 26708 3508 26709 3548
rect 26667 3499 26709 3508
rect 26572 3415 26612 3424
rect 26379 3380 26421 3389
rect 26764 3380 26804 4684
rect 26860 4397 26900 4768
rect 26859 4388 26901 4397
rect 26859 4348 26860 4388
rect 26900 4348 26901 4388
rect 26859 4339 26901 4348
rect 26859 4220 26901 4229
rect 26859 4180 26860 4220
rect 26900 4180 26901 4220
rect 26859 4171 26901 4180
rect 26860 4136 26900 4171
rect 26860 4085 26900 4096
rect 26956 3464 26996 4843
rect 27052 4724 27092 4733
rect 27092 4684 27188 4724
rect 27052 4675 27092 4684
rect 26956 3415 26996 3424
rect 27052 3968 27092 3977
rect 26379 3340 26380 3380
rect 26420 3340 26421 3380
rect 26379 3331 26421 3340
rect 26668 3340 26804 3380
rect 26380 3212 26420 3221
rect 26380 1877 26420 3172
rect 26668 2540 26708 3340
rect 26764 3212 26804 3221
rect 26955 3212 26997 3221
rect 26804 3172 26900 3212
rect 26764 3163 26804 3172
rect 26668 2500 26804 2540
rect 26379 1868 26421 1877
rect 26379 1828 26380 1868
rect 26420 1828 26421 1868
rect 26379 1819 26421 1828
rect 26379 1700 26421 1709
rect 26379 1660 26380 1700
rect 26420 1660 26421 1700
rect 26379 1651 26421 1660
rect 26283 1028 26325 1037
rect 26283 988 26284 1028
rect 26324 988 26325 1028
rect 26283 979 26325 988
rect 26380 80 26420 1651
rect 26571 1196 26613 1205
rect 26571 1156 26572 1196
rect 26612 1156 26613 1196
rect 26571 1147 26613 1156
rect 26572 80 26612 1147
rect 26764 80 26804 2500
rect 26860 1541 26900 3172
rect 26955 3172 26956 3212
rect 26996 3172 26997 3212
rect 26955 3163 26997 3172
rect 26859 1532 26901 1541
rect 26859 1492 26860 1532
rect 26900 1492 26901 1532
rect 26859 1483 26901 1492
rect 26956 80 26996 3163
rect 27052 2717 27092 3928
rect 27148 3380 27188 4684
rect 27243 4472 27285 4481
rect 27243 4432 27244 4472
rect 27284 4432 27285 4472
rect 27243 4423 27285 4432
rect 27244 4220 27284 4423
rect 27244 3977 27284 4180
rect 27243 3968 27285 3977
rect 27243 3928 27244 3968
rect 27284 3928 27285 3968
rect 27243 3919 27285 3928
rect 27340 3464 27380 5608
rect 27627 5608 27628 5648
rect 27668 5608 27669 5648
rect 27627 5599 27669 5608
rect 27820 5480 27860 6280
rect 27724 5440 27860 5480
rect 27627 4892 27669 4901
rect 27627 4852 27628 4892
rect 27668 4852 27669 4892
rect 27627 4843 27669 4852
rect 27628 4758 27668 4843
rect 27436 4724 27476 4733
rect 27476 4684 27572 4724
rect 27436 4675 27476 4684
rect 27435 4220 27477 4229
rect 27435 4180 27436 4220
rect 27476 4180 27477 4220
rect 27435 4171 27477 4180
rect 27436 4086 27476 4171
rect 27436 3968 27476 3977
rect 27436 3473 27476 3928
rect 27532 3632 27572 4684
rect 27627 4220 27669 4229
rect 27627 4180 27628 4220
rect 27668 4180 27669 4220
rect 27627 4171 27669 4180
rect 27628 4086 27668 4171
rect 27724 4145 27764 5440
rect 27819 5312 27861 5321
rect 27819 5272 27820 5312
rect 27860 5272 27861 5312
rect 27819 5263 27861 5272
rect 27820 5144 27860 5263
rect 28012 5228 28052 6616
rect 28108 5909 28148 7792
rect 28204 7589 28244 7876
rect 28395 7916 28437 7925
rect 28395 7876 28396 7916
rect 28436 7876 28437 7916
rect 28395 7867 28437 7876
rect 28588 7916 28628 8287
rect 28684 8261 28724 8623
rect 28683 8252 28725 8261
rect 28683 8212 28684 8252
rect 28724 8212 28725 8252
rect 28683 8203 28725 8212
rect 28876 8009 28916 8716
rect 28971 8084 29013 8093
rect 28971 8044 28972 8084
rect 29012 8044 29013 8084
rect 28971 8035 29013 8044
rect 28875 8000 28917 8009
rect 28875 7960 28876 8000
rect 28916 7960 28917 8000
rect 28875 7951 28917 7960
rect 28972 7925 29012 8035
rect 28396 7782 28436 7867
rect 28492 7832 28532 7841
rect 28203 7580 28245 7589
rect 28203 7540 28204 7580
rect 28244 7540 28245 7580
rect 28203 7531 28245 7540
rect 28395 6824 28437 6833
rect 28395 6784 28396 6824
rect 28436 6784 28437 6824
rect 28395 6775 28437 6784
rect 28107 5900 28149 5909
rect 28107 5860 28108 5900
rect 28148 5860 28149 5900
rect 28107 5851 28149 5860
rect 28108 5648 28148 5657
rect 28108 5321 28148 5608
rect 28300 5480 28340 5489
rect 28107 5312 28149 5321
rect 28107 5272 28108 5312
rect 28148 5272 28149 5312
rect 28107 5263 28149 5272
rect 27820 5095 27860 5104
rect 27916 5188 28052 5228
rect 27819 4892 27861 4901
rect 27819 4852 27820 4892
rect 27860 4852 27861 4892
rect 27819 4843 27861 4852
rect 27820 4758 27860 4843
rect 27819 4640 27861 4649
rect 27819 4600 27820 4640
rect 27860 4600 27861 4640
rect 27819 4591 27861 4600
rect 27820 4220 27860 4591
rect 27916 4481 27956 5188
rect 28012 4901 28052 4986
rect 28011 4892 28053 4901
rect 28011 4852 28012 4892
rect 28052 4852 28053 4892
rect 28011 4843 28053 4852
rect 28204 4892 28244 4901
rect 28011 4841 28052 4843
rect 27915 4472 27957 4481
rect 27915 4432 27916 4472
rect 27956 4432 27957 4472
rect 27915 4423 27957 4432
rect 28012 4229 28052 4841
rect 28107 4724 28149 4733
rect 28107 4684 28108 4724
rect 28148 4684 28149 4724
rect 28107 4675 28149 4684
rect 28108 4590 28148 4675
rect 28204 4565 28244 4852
rect 28203 4556 28245 4565
rect 28203 4516 28204 4556
rect 28244 4516 28245 4556
rect 28203 4507 28245 4516
rect 28203 4304 28245 4313
rect 28203 4264 28204 4304
rect 28244 4264 28245 4304
rect 28203 4255 28245 4264
rect 27820 4171 27860 4180
rect 28011 4220 28053 4229
rect 28011 4180 28012 4220
rect 28052 4180 28053 4220
rect 28011 4171 28053 4180
rect 28204 4220 28244 4255
rect 28204 4169 28244 4180
rect 27723 4136 27765 4145
rect 27723 4096 27724 4136
rect 27764 4096 27765 4136
rect 27723 4087 27765 4096
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 27628 3968 27668 3977
rect 27628 3809 27668 3928
rect 28012 3918 28052 4003
rect 28300 3968 28340 5440
rect 28396 5321 28436 6775
rect 28492 6572 28532 7792
rect 28588 7757 28628 7876
rect 28779 7916 28821 7925
rect 28779 7876 28780 7916
rect 28820 7876 28821 7916
rect 28779 7867 28821 7876
rect 28971 7916 29013 7925
rect 28971 7876 28972 7916
rect 29012 7876 29013 7916
rect 28971 7867 29013 7876
rect 28780 7782 28820 7867
rect 28876 7832 28916 7841
rect 28587 7748 28629 7757
rect 28587 7708 28588 7748
rect 28628 7708 28629 7748
rect 28587 7699 28629 7708
rect 28492 6532 28628 6572
rect 28491 6404 28533 6413
rect 28491 6364 28492 6404
rect 28532 6364 28533 6404
rect 28491 6355 28533 6364
rect 28492 6270 28532 6355
rect 28492 5741 28532 5826
rect 28491 5732 28533 5741
rect 28491 5692 28492 5732
rect 28532 5692 28533 5732
rect 28491 5683 28533 5692
rect 28491 5480 28533 5489
rect 28491 5440 28492 5480
rect 28532 5440 28533 5480
rect 28491 5431 28533 5440
rect 28492 5346 28532 5431
rect 28395 5312 28437 5321
rect 28395 5272 28396 5312
rect 28436 5272 28437 5312
rect 28395 5263 28437 5272
rect 28396 5069 28436 5154
rect 28588 5144 28628 6532
rect 28683 6404 28725 6413
rect 28683 6364 28684 6404
rect 28724 6364 28725 6404
rect 28683 6355 28725 6364
rect 28684 6270 28724 6355
rect 28684 5732 28724 5741
rect 28684 5321 28724 5692
rect 28779 5732 28821 5741
rect 28779 5692 28780 5732
rect 28820 5692 28821 5732
rect 28779 5683 28821 5692
rect 28683 5312 28725 5321
rect 28683 5272 28684 5312
rect 28724 5272 28725 5312
rect 28683 5263 28725 5272
rect 28588 5104 28724 5144
rect 28395 5060 28437 5069
rect 28395 5020 28396 5060
rect 28436 5020 28437 5060
rect 28395 5011 28437 5020
rect 28396 4892 28436 4903
rect 28396 4817 28436 4852
rect 28588 4892 28628 4901
rect 28395 4808 28437 4817
rect 28395 4768 28396 4808
rect 28436 4768 28437 4808
rect 28395 4759 28437 4768
rect 28588 4724 28628 4852
rect 28492 4684 28628 4724
rect 28395 4136 28437 4145
rect 28395 4096 28396 4136
rect 28436 4096 28437 4136
rect 28395 4087 28437 4096
rect 28396 4002 28436 4087
rect 28204 3928 28340 3968
rect 27627 3800 27669 3809
rect 27627 3760 27628 3800
rect 27668 3760 27669 3800
rect 27627 3751 27669 3760
rect 27532 3592 27860 3632
rect 27340 3415 27380 3424
rect 27435 3464 27477 3473
rect 27435 3424 27436 3464
rect 27476 3424 27477 3464
rect 27435 3415 27477 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 27724 3464 27764 3473
rect 27148 3340 27284 3380
rect 27148 3212 27188 3221
rect 27051 2708 27093 2717
rect 27051 2668 27052 2708
rect 27092 2668 27093 2708
rect 27051 2659 27093 2668
rect 27148 1373 27188 3172
rect 27244 2540 27284 3340
rect 27532 3212 27572 3221
rect 27436 3172 27532 3212
rect 27244 2500 27380 2540
rect 27147 1364 27189 1373
rect 27147 1324 27148 1364
rect 27188 1324 27189 1364
rect 27147 1315 27189 1324
rect 27147 1028 27189 1037
rect 27147 988 27148 1028
rect 27188 988 27189 1028
rect 27147 979 27189 988
rect 27148 80 27188 979
rect 27340 80 27380 2500
rect 27436 1625 27476 3172
rect 27532 3163 27572 3172
rect 27628 2540 27668 3415
rect 27724 3305 27764 3424
rect 27723 3296 27765 3305
rect 27723 3256 27724 3296
rect 27764 3256 27765 3296
rect 27723 3247 27765 3256
rect 27820 2540 27860 3592
rect 28107 3464 28149 3473
rect 28107 3424 28108 3464
rect 28148 3424 28149 3464
rect 28107 3415 28149 3424
rect 28108 3330 28148 3415
rect 27915 3212 27957 3221
rect 27915 3172 27916 3212
rect 27956 3172 27957 3212
rect 27915 3163 27957 3172
rect 27916 3078 27956 3163
rect 28204 2540 28244 3928
rect 28492 3893 28532 4684
rect 28587 4556 28629 4565
rect 28587 4516 28588 4556
rect 28628 4516 28629 4556
rect 28587 4507 28629 4516
rect 28588 4145 28628 4507
rect 28587 4136 28629 4145
rect 28587 4096 28588 4136
rect 28628 4096 28629 4136
rect 28587 4087 28629 4096
rect 28588 3968 28628 3977
rect 28491 3884 28533 3893
rect 28491 3844 28492 3884
rect 28532 3844 28533 3884
rect 28491 3835 28533 3844
rect 28491 3716 28533 3725
rect 28491 3676 28492 3716
rect 28532 3676 28533 3716
rect 28491 3667 28533 3676
rect 28492 3464 28532 3667
rect 28492 3415 28532 3424
rect 28300 3212 28340 3221
rect 28340 3172 28436 3212
rect 28300 3163 28340 3172
rect 27628 2500 27764 2540
rect 27820 2500 27956 2540
rect 28204 2500 28340 2540
rect 27531 2456 27573 2465
rect 27531 2416 27532 2456
rect 27572 2416 27573 2456
rect 27531 2407 27573 2416
rect 27435 1616 27477 1625
rect 27435 1576 27436 1616
rect 27476 1576 27477 1616
rect 27435 1567 27477 1576
rect 27532 80 27572 2407
rect 27724 80 27764 2500
rect 27916 80 27956 2500
rect 28107 1784 28149 1793
rect 28107 1744 28108 1784
rect 28148 1744 28149 1784
rect 28107 1735 28149 1744
rect 28108 80 28148 1735
rect 28300 80 28340 2500
rect 28396 1037 28436 3172
rect 28491 2708 28533 2717
rect 28491 2668 28492 2708
rect 28532 2668 28533 2708
rect 28491 2659 28533 2668
rect 28395 1028 28437 1037
rect 28395 988 28396 1028
rect 28436 988 28437 1028
rect 28395 979 28437 988
rect 28492 80 28532 2659
rect 28588 1289 28628 3928
rect 28684 3809 28724 5104
rect 28780 4892 28820 5683
rect 28876 4901 28916 7792
rect 28972 7782 29012 7867
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 28971 5732 29013 5741
rect 28971 5692 28972 5732
rect 29012 5692 29013 5732
rect 28971 5683 29013 5692
rect 29164 5732 29204 6439
rect 29164 5683 29204 5692
rect 28972 5598 29012 5683
rect 29260 5564 29300 10639
rect 30316 10604 30356 11236
rect 30892 11192 30932 11236
rect 30892 11143 30932 11152
rect 30603 11108 30645 11117
rect 30603 11068 30604 11108
rect 30644 11068 30645 11108
rect 30603 11059 30645 11068
rect 31371 11108 31413 11117
rect 31371 11068 31372 11108
rect 31412 11068 31413 11108
rect 31371 11059 31413 11068
rect 30507 10940 30549 10949
rect 30507 10900 30508 10940
rect 30548 10900 30549 10940
rect 30507 10891 30549 10900
rect 30124 10564 30356 10604
rect 29643 9512 29685 9521
rect 29643 9472 29644 9512
rect 29684 9472 29685 9512
rect 29643 9463 29685 9472
rect 29355 8756 29397 8765
rect 29355 8716 29356 8756
rect 29396 8716 29397 8756
rect 29355 8707 29397 8716
rect 29547 8756 29589 8765
rect 29547 8716 29548 8756
rect 29588 8716 29589 8756
rect 29547 8707 29589 8716
rect 29356 8622 29396 8707
rect 29548 8622 29588 8707
rect 29547 7412 29589 7421
rect 29547 7372 29548 7412
rect 29588 7372 29589 7412
rect 29547 7363 29589 7372
rect 29548 5648 29588 7363
rect 29644 5648 29684 9463
rect 30028 9428 30068 9437
rect 30028 8765 30068 9388
rect 30124 9260 30164 10564
rect 30219 10436 30261 10445
rect 30411 10436 30453 10445
rect 30219 10396 30220 10436
rect 30260 10396 30356 10436
rect 30219 10387 30261 10396
rect 30316 10277 30356 10396
rect 30411 10396 30412 10436
rect 30452 10396 30453 10436
rect 30411 10387 30453 10396
rect 30220 10268 30260 10277
rect 30220 9428 30260 10228
rect 30315 10268 30357 10277
rect 30315 10228 30316 10268
rect 30356 10228 30357 10268
rect 30315 10219 30357 10228
rect 30412 10268 30452 10387
rect 30412 10109 30452 10228
rect 30316 10100 30356 10109
rect 30316 9941 30356 10060
rect 30411 10100 30453 10109
rect 30411 10060 30412 10100
rect 30452 10060 30453 10100
rect 30411 10051 30453 10060
rect 30315 9932 30357 9941
rect 30315 9892 30316 9932
rect 30356 9892 30357 9932
rect 30315 9883 30357 9892
rect 30508 9605 30548 10891
rect 30604 10865 30644 11059
rect 30987 11024 31029 11033
rect 30987 10984 30988 11024
rect 31028 10984 31029 11024
rect 30987 10975 31029 10984
rect 30795 10940 30837 10949
rect 30700 10900 30796 10940
rect 30836 10900 30837 10940
rect 30603 10856 30645 10865
rect 30603 10816 30604 10856
rect 30644 10816 30645 10856
rect 30603 10807 30645 10816
rect 30604 10268 30644 10277
rect 30700 10268 30740 10900
rect 30795 10891 30837 10900
rect 30988 10940 31028 10975
rect 30796 10806 30836 10891
rect 30988 10889 31028 10900
rect 31179 10940 31221 10949
rect 31179 10900 31180 10940
rect 31220 10900 31221 10940
rect 31179 10891 31221 10900
rect 31372 10940 31412 11059
rect 36171 11024 36213 11033
rect 36171 10984 36172 11024
rect 36212 10984 36213 11024
rect 36171 10975 36213 10984
rect 31083 10856 31125 10865
rect 31083 10816 31084 10856
rect 31124 10816 31125 10856
rect 31083 10807 31125 10816
rect 30795 10688 30837 10697
rect 30987 10688 31029 10697
rect 30795 10648 30796 10688
rect 30836 10648 30837 10688
rect 30795 10639 30837 10648
rect 30892 10648 30988 10688
rect 31028 10648 31029 10688
rect 30796 10277 30836 10639
rect 30644 10228 30740 10268
rect 30795 10268 30837 10277
rect 30795 10228 30796 10268
rect 30836 10228 30837 10268
rect 30604 10025 30644 10228
rect 30795 10219 30837 10228
rect 30796 10134 30836 10219
rect 30699 10100 30741 10109
rect 30699 10060 30700 10100
rect 30740 10060 30741 10100
rect 30699 10051 30741 10060
rect 30603 10016 30645 10025
rect 30603 9976 30604 10016
rect 30644 9976 30645 10016
rect 30603 9967 30645 9976
rect 30507 9596 30549 9605
rect 30507 9556 30508 9596
rect 30548 9556 30549 9596
rect 30507 9547 30549 9556
rect 30604 9428 30644 9967
rect 30700 9966 30740 10051
rect 30892 9773 30932 10648
rect 30987 10639 31029 10648
rect 30988 10268 31028 10277
rect 30988 10025 31028 10228
rect 31084 10184 31124 10807
rect 31180 10806 31220 10891
rect 31276 10856 31316 10865
rect 31180 10361 31220 10384
rect 31179 10352 31221 10361
rect 31179 10312 31180 10352
rect 31220 10312 31221 10352
rect 31179 10303 31221 10312
rect 31180 10289 31220 10303
rect 31180 10240 31220 10249
rect 31084 10144 31220 10184
rect 30987 10016 31029 10025
rect 30987 9976 30988 10016
rect 31028 9976 31029 10016
rect 30987 9967 31029 9976
rect 31084 10016 31124 10025
rect 30891 9764 30933 9773
rect 30891 9724 30892 9764
rect 30932 9724 30933 9764
rect 30891 9715 30933 9724
rect 31084 9605 31124 9976
rect 31083 9596 31125 9605
rect 31083 9556 31084 9596
rect 31124 9556 31125 9596
rect 31083 9547 31125 9556
rect 30891 9512 30933 9521
rect 30891 9472 30892 9512
rect 30932 9472 30933 9512
rect 30891 9463 30933 9472
rect 30260 9388 30604 9428
rect 30220 9379 30260 9388
rect 30604 9269 30644 9388
rect 30795 9428 30837 9437
rect 30795 9388 30796 9428
rect 30836 9388 30837 9428
rect 30795 9379 30837 9388
rect 30700 9344 30740 9353
rect 30603 9260 30645 9269
rect 30124 9220 30356 9260
rect 30027 8756 30069 8765
rect 30027 8716 30028 8756
rect 30068 8716 30069 8756
rect 30027 8707 30069 8716
rect 30219 8756 30261 8765
rect 30219 8716 30220 8756
rect 30260 8716 30261 8756
rect 30219 8707 30261 8716
rect 30220 8168 30260 8707
rect 30220 8119 30260 8128
rect 29932 7916 29972 7925
rect 29836 7876 29932 7916
rect 29740 7706 29780 7715
rect 29740 7076 29780 7666
rect 29836 7169 29876 7876
rect 29932 7867 29972 7876
rect 30028 7916 30068 7925
rect 30028 7505 30068 7876
rect 30027 7496 30069 7505
rect 30027 7456 30028 7496
rect 30068 7456 30069 7496
rect 30027 7447 30069 7456
rect 30027 7244 30069 7253
rect 30027 7204 30028 7244
rect 30068 7204 30069 7244
rect 30027 7195 30069 7204
rect 29835 7160 29877 7169
rect 29835 7120 29836 7160
rect 29876 7120 29877 7160
rect 29835 7111 29877 7120
rect 29740 6833 29780 7036
rect 29739 6824 29781 6833
rect 29739 6784 29740 6824
rect 29780 6784 29781 6824
rect 29739 6775 29781 6784
rect 29740 6404 29780 6775
rect 29836 6446 29876 7111
rect 30028 7110 30068 7195
rect 29932 6572 29972 6581
rect 29972 6532 30164 6572
rect 29932 6523 29972 6532
rect 29836 6406 29972 6446
rect 29740 6355 29780 6364
rect 29932 6404 29972 6406
rect 29932 6355 29972 6364
rect 30027 6404 30069 6413
rect 30027 6364 30028 6404
rect 30068 6364 30069 6404
rect 30027 6355 30069 6364
rect 29835 6320 29877 6329
rect 29835 6280 29836 6320
rect 29876 6280 29877 6320
rect 29835 6271 29877 6280
rect 29836 6152 29876 6271
rect 30028 6270 30068 6355
rect 29836 6112 30068 6152
rect 29932 5648 29972 5657
rect 29644 5608 29932 5648
rect 29548 5599 29588 5608
rect 29932 5599 29972 5608
rect 29164 5524 29300 5564
rect 28971 5228 29013 5237
rect 28971 5188 28972 5228
rect 29012 5188 29013 5228
rect 28971 5179 29013 5188
rect 28780 4817 28820 4852
rect 28875 4892 28917 4901
rect 28875 4852 28876 4892
rect 28916 4852 28917 4892
rect 28875 4843 28917 4852
rect 28972 4892 29012 5179
rect 29164 4976 29204 5524
rect 29356 5480 29396 5489
rect 29740 5480 29780 5489
rect 29164 4927 29204 4936
rect 29260 5440 29356 5480
rect 28972 4843 29012 4852
rect 28779 4808 28821 4817
rect 28779 4768 28780 4808
rect 28820 4768 28821 4808
rect 28779 4759 28821 4768
rect 28780 4728 28820 4759
rect 28876 4724 28916 4733
rect 28971 4724 29013 4733
rect 28916 4684 28972 4724
rect 29012 4684 29013 4724
rect 28876 4675 28916 4684
rect 28971 4675 29013 4684
rect 29163 4556 29205 4565
rect 29163 4516 29164 4556
rect 29204 4516 29205 4556
rect 29163 4507 29205 4516
rect 28875 4388 28917 4397
rect 28875 4348 28876 4388
rect 28916 4348 28917 4388
rect 28875 4339 28917 4348
rect 28779 4220 28821 4229
rect 28779 4180 28780 4220
rect 28820 4180 28821 4220
rect 28779 4171 28821 4180
rect 28780 4136 28820 4171
rect 28780 4085 28820 4096
rect 28683 3800 28725 3809
rect 28683 3760 28684 3800
rect 28724 3760 28725 3800
rect 28683 3751 28725 3760
rect 28876 3464 28916 4339
rect 29164 4304 29204 4507
rect 29260 4472 29300 5440
rect 29356 5431 29396 5440
rect 29644 5440 29740 5480
rect 29451 5312 29493 5321
rect 29451 5272 29452 5312
rect 29492 5272 29493 5312
rect 29451 5263 29493 5272
rect 29355 4724 29397 4733
rect 29355 4684 29356 4724
rect 29396 4684 29397 4724
rect 29355 4675 29397 4684
rect 29356 4590 29396 4675
rect 29260 4432 29396 4472
rect 29164 4264 29300 4304
rect 29260 4219 29300 4264
rect 29260 4170 29300 4179
rect 29260 4052 29300 4061
rect 29260 3977 29300 4012
rect 28876 3415 28916 3424
rect 28972 3968 29012 3977
rect 28684 3212 28724 3221
rect 28684 2717 28724 3172
rect 28683 2708 28725 2717
rect 28683 2668 28684 2708
rect 28724 2668 28725 2708
rect 28683 2659 28725 2668
rect 28683 1868 28725 1877
rect 28683 1828 28684 1868
rect 28724 1828 28725 1868
rect 28683 1819 28725 1828
rect 28587 1280 28629 1289
rect 28587 1240 28588 1280
rect 28628 1240 28629 1280
rect 28587 1231 28629 1240
rect 28684 80 28724 1819
rect 28875 1532 28917 1541
rect 28875 1492 28876 1532
rect 28916 1492 28917 1532
rect 28875 1483 28917 1492
rect 28876 80 28916 1483
rect 28972 1205 29012 3928
rect 29260 3968 29302 3977
rect 29260 3928 29261 3968
rect 29301 3928 29302 3968
rect 29260 3919 29302 3928
rect 29259 3800 29301 3809
rect 29259 3760 29260 3800
rect 29300 3760 29301 3800
rect 29259 3751 29301 3760
rect 29260 3464 29300 3751
rect 29260 3415 29300 3424
rect 29068 3212 29108 3221
rect 29068 2801 29108 3172
rect 29067 2792 29109 2801
rect 29067 2752 29068 2792
rect 29108 2752 29109 2792
rect 29067 2743 29109 2752
rect 29356 2540 29396 4432
rect 29452 4220 29492 5263
rect 29547 5144 29589 5153
rect 29547 5104 29548 5144
rect 29588 5104 29589 5144
rect 29547 5095 29589 5104
rect 29548 4976 29588 5095
rect 29548 4927 29588 4936
rect 29452 4061 29492 4180
rect 29451 4052 29493 4061
rect 29451 4012 29452 4052
rect 29492 4012 29493 4052
rect 29451 4003 29493 4012
rect 29644 3632 29684 5440
rect 29740 5431 29780 5440
rect 29932 4976 29972 4985
rect 30028 4976 30068 6112
rect 30124 5741 30164 6532
rect 30316 6161 30356 9220
rect 30603 9220 30604 9260
rect 30644 9220 30645 9260
rect 30603 9211 30645 9220
rect 30700 9101 30740 9304
rect 30796 9294 30836 9379
rect 30699 9092 30741 9101
rect 30699 9052 30700 9092
rect 30740 9052 30741 9092
rect 30699 9043 30741 9052
rect 30892 8420 30932 9463
rect 31084 9428 31124 9437
rect 30988 9415 31028 9424
rect 30988 9269 31028 9375
rect 30987 9260 31029 9269
rect 30987 9220 30988 9260
rect 31028 9220 31029 9260
rect 30987 9211 31029 9220
rect 31084 9017 31124 9388
rect 31180 9428 31220 10144
rect 31180 9379 31220 9388
rect 31083 9008 31125 9017
rect 31083 8968 31084 9008
rect 31124 8968 31125 9008
rect 31083 8959 31125 8968
rect 30700 8380 30932 8420
rect 30412 7160 30452 7169
rect 30315 6152 30357 6161
rect 30315 6112 30316 6152
rect 30356 6112 30357 6152
rect 30315 6103 30357 6112
rect 30315 5900 30357 5909
rect 30315 5860 30316 5900
rect 30356 5860 30357 5900
rect 30315 5851 30357 5860
rect 30123 5732 30165 5741
rect 30123 5692 30124 5732
rect 30164 5692 30165 5732
rect 30123 5683 30165 5692
rect 30316 5732 30356 5851
rect 30316 5683 30356 5692
rect 30124 5598 30164 5683
rect 30412 5657 30452 7120
rect 30603 5732 30645 5741
rect 30603 5692 30604 5732
rect 30644 5692 30645 5732
rect 30603 5683 30645 5692
rect 30411 5648 30453 5657
rect 30411 5608 30412 5648
rect 30452 5608 30453 5648
rect 30411 5599 30453 5608
rect 30604 5598 30644 5683
rect 30507 5564 30549 5573
rect 30507 5524 30508 5564
rect 30548 5524 30549 5564
rect 30507 5515 30549 5524
rect 30411 5480 30453 5489
rect 30411 5440 30412 5480
rect 30452 5440 30453 5480
rect 30411 5431 30453 5440
rect 29972 4936 30068 4976
rect 29932 4927 29972 4936
rect 30316 4892 30356 4901
rect 30316 4733 30356 4852
rect 29548 3592 29684 3632
rect 29740 4724 29780 4733
rect 29260 2500 29396 2540
rect 29452 3212 29492 3221
rect 29067 1364 29109 1373
rect 29067 1324 29068 1364
rect 29108 1324 29109 1364
rect 29067 1315 29109 1324
rect 28971 1196 29013 1205
rect 28971 1156 28972 1196
rect 29012 1156 29013 1196
rect 28971 1147 29013 1156
rect 29068 80 29108 1315
rect 29260 80 29300 2500
rect 29452 1793 29492 3172
rect 29548 2540 29588 3592
rect 29643 3464 29685 3473
rect 29643 3424 29644 3464
rect 29684 3424 29685 3464
rect 29643 3415 29685 3424
rect 29644 3330 29684 3415
rect 29548 2500 29684 2540
rect 29451 1784 29493 1793
rect 29451 1744 29452 1784
rect 29492 1744 29493 1784
rect 29451 1735 29493 1744
rect 29451 1616 29493 1625
rect 29451 1576 29452 1616
rect 29492 1576 29493 1616
rect 29451 1567 29493 1576
rect 29452 80 29492 1567
rect 29644 80 29684 2500
rect 29740 953 29780 4684
rect 29835 4724 29877 4733
rect 30124 4724 30164 4733
rect 29835 4684 29836 4724
rect 29876 4684 29877 4724
rect 29835 4675 29877 4684
rect 30028 4684 30124 4724
rect 29836 3632 29876 4675
rect 29931 4220 29973 4229
rect 29931 4180 29932 4220
rect 29972 4180 29973 4220
rect 29931 4171 29973 4180
rect 29932 4086 29972 4171
rect 30028 3632 30068 4684
rect 30124 4675 30164 4684
rect 30315 4724 30357 4733
rect 30315 4684 30316 4724
rect 30356 4684 30357 4724
rect 30315 4675 30357 4684
rect 30219 4640 30261 4649
rect 30219 4600 30220 4640
rect 30260 4600 30261 4640
rect 30219 4591 30261 4600
rect 30123 4220 30165 4229
rect 30123 4180 30124 4220
rect 30164 4180 30165 4220
rect 30123 4171 30165 4180
rect 30124 4086 30164 4171
rect 30124 3968 30164 3977
rect 30220 3968 30260 4591
rect 30315 4220 30357 4229
rect 30315 4180 30316 4220
rect 30356 4180 30357 4220
rect 30315 4171 30357 4180
rect 30316 4086 30356 4171
rect 30164 3928 30260 3968
rect 30316 3968 30356 3977
rect 30124 3919 30164 3928
rect 29836 3592 29972 3632
rect 30028 3592 30164 3632
rect 29836 3212 29876 3221
rect 29836 1700 29876 3172
rect 29932 2372 29972 3592
rect 30028 3464 30068 3475
rect 30028 3389 30068 3424
rect 30027 3380 30069 3389
rect 30027 3340 30028 3380
rect 30068 3340 30069 3380
rect 30027 3331 30069 3340
rect 29932 2332 30068 2372
rect 29836 1660 29972 1700
rect 29932 1373 29972 1660
rect 29931 1364 29973 1373
rect 29931 1324 29932 1364
rect 29972 1324 29973 1364
rect 29931 1315 29973 1324
rect 29835 1280 29877 1289
rect 29835 1240 29836 1280
rect 29876 1240 29877 1280
rect 29835 1231 29877 1240
rect 29739 944 29781 953
rect 29739 904 29740 944
rect 29780 904 29781 944
rect 29739 895 29781 904
rect 29836 80 29876 1231
rect 30028 80 30068 2332
rect 30124 1121 30164 3592
rect 30316 3473 30356 3928
rect 30315 3464 30357 3473
rect 30315 3424 30316 3464
rect 30356 3424 30357 3464
rect 30315 3415 30357 3424
rect 30412 3464 30452 5431
rect 30508 5144 30548 5515
rect 30603 5228 30645 5237
rect 30603 5188 30604 5228
rect 30644 5188 30645 5228
rect 30603 5179 30645 5188
rect 30508 5095 30548 5104
rect 30507 4892 30549 4901
rect 30507 4852 30508 4892
rect 30548 4852 30549 4892
rect 30507 4843 30549 4852
rect 30508 4758 30548 4843
rect 30508 4220 30548 4229
rect 30604 4220 30644 5179
rect 30700 5153 30740 8380
rect 30795 8252 30837 8261
rect 30795 8212 30796 8252
rect 30836 8212 30837 8252
rect 30795 8203 30837 8212
rect 30796 7925 30836 8203
rect 31276 8093 31316 10816
rect 31372 10697 31412 10900
rect 36075 10940 36117 10949
rect 36075 10900 36076 10940
rect 36116 10900 36117 10940
rect 36075 10891 36117 10900
rect 31371 10688 31413 10697
rect 31371 10648 31372 10688
rect 31412 10648 31413 10688
rect 31371 10639 31413 10648
rect 31563 10604 31605 10613
rect 31563 10564 31564 10604
rect 31604 10564 31605 10604
rect 31563 10555 31605 10564
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 31372 10268 31412 10277
rect 31372 10025 31412 10228
rect 31564 10268 31604 10555
rect 31947 10520 31989 10529
rect 31947 10480 31948 10520
rect 31988 10480 31989 10520
rect 31947 10471 31989 10480
rect 31564 10193 31604 10228
rect 31563 10184 31605 10193
rect 31563 10144 31564 10184
rect 31604 10144 31605 10184
rect 31563 10135 31605 10144
rect 31564 10104 31604 10135
rect 31371 10016 31413 10025
rect 31371 9976 31372 10016
rect 31412 9976 31413 10016
rect 31371 9967 31413 9976
rect 31468 10016 31508 10025
rect 31508 9976 31892 10016
rect 31468 9967 31508 9976
rect 31755 8672 31797 8681
rect 31755 8632 31756 8672
rect 31796 8632 31797 8672
rect 31755 8623 31797 8632
rect 31275 8084 31317 8093
rect 31275 8044 31276 8084
rect 31316 8044 31317 8084
rect 31275 8035 31317 8044
rect 30795 7916 30837 7925
rect 30795 7876 30796 7916
rect 30836 7876 30837 7916
rect 30795 7867 30837 7876
rect 30987 7916 31029 7925
rect 30987 7876 30988 7916
rect 31028 7876 31029 7916
rect 30987 7867 31029 7876
rect 31179 7916 31221 7925
rect 31179 7876 31180 7916
rect 31220 7876 31221 7916
rect 31179 7867 31221 7876
rect 31372 7916 31412 7925
rect 30796 7782 30836 7867
rect 30891 7832 30933 7841
rect 30891 7792 30892 7832
rect 30932 7792 30933 7832
rect 30891 7783 30933 7792
rect 30892 7698 30932 7783
rect 30988 7782 31028 7867
rect 31180 7782 31220 7867
rect 31275 7832 31317 7841
rect 31275 7792 31276 7832
rect 31316 7792 31317 7832
rect 31275 7783 31317 7792
rect 31276 7698 31316 7783
rect 31372 7757 31412 7876
rect 31563 7916 31605 7925
rect 31563 7876 31564 7916
rect 31604 7876 31605 7916
rect 31563 7867 31605 7876
rect 31756 7916 31796 8623
rect 31756 7867 31796 7876
rect 31564 7782 31604 7867
rect 31659 7832 31701 7841
rect 31659 7792 31660 7832
rect 31700 7792 31701 7832
rect 31659 7783 31701 7792
rect 31371 7748 31413 7757
rect 31371 7708 31372 7748
rect 31412 7708 31413 7748
rect 31371 7699 31413 7708
rect 31660 7698 31700 7783
rect 30987 7496 31029 7505
rect 30987 7456 30988 7496
rect 31028 7456 31029 7496
rect 30987 7447 31029 7456
rect 30988 7001 31028 7447
rect 31852 7412 31892 9976
rect 31948 8924 31988 10471
rect 35595 10436 35637 10445
rect 35595 10396 35596 10436
rect 35636 10396 35637 10436
rect 35595 10387 35637 10396
rect 32044 10268 32084 10277
rect 35596 10268 35636 10387
rect 36076 10352 36116 10891
rect 36172 10529 36212 10975
rect 36460 10940 36500 10949
rect 36364 10900 36460 10940
rect 36171 10520 36213 10529
rect 36171 10480 36172 10520
rect 36212 10480 36213 10520
rect 36171 10471 36213 10480
rect 36076 10303 36116 10312
rect 32084 10228 32180 10268
rect 32044 10219 32084 10228
rect 32043 10016 32085 10025
rect 32043 9976 32044 10016
rect 32084 9976 32085 10016
rect 32043 9967 32085 9976
rect 32044 9882 32084 9967
rect 31948 8875 31988 8884
rect 32140 8756 32180 10228
rect 35596 10219 35636 10228
rect 35787 10268 35829 10277
rect 35787 10228 35788 10268
rect 35828 10228 35829 10268
rect 35787 10219 35829 10228
rect 35979 10268 36021 10277
rect 35979 10228 35980 10268
rect 36020 10228 36021 10268
rect 35979 10219 36021 10228
rect 36172 10268 36212 10471
rect 36364 10277 36404 10900
rect 36460 10891 36500 10900
rect 36652 10940 36692 10949
rect 36844 10940 36884 10949
rect 36556 10856 36596 10865
rect 36459 10688 36501 10697
rect 36459 10648 36460 10688
rect 36500 10648 36501 10688
rect 36459 10639 36501 10648
rect 36460 10352 36500 10639
rect 36556 10436 36596 10816
rect 36652 10781 36692 10900
rect 36748 10900 36844 10940
rect 36651 10772 36693 10781
rect 36651 10732 36652 10772
rect 36692 10732 36693 10772
rect 36651 10723 36693 10732
rect 36652 10613 36692 10723
rect 36651 10604 36693 10613
rect 36651 10564 36652 10604
rect 36692 10564 36693 10604
rect 36651 10555 36693 10564
rect 36556 10396 36692 10436
rect 36460 10303 36500 10312
rect 36363 10268 36405 10277
rect 36172 10219 36212 10228
rect 36268 10228 36364 10268
rect 36404 10228 36405 10268
rect 32236 10184 32276 10193
rect 32236 9437 32276 10144
rect 35788 10134 35828 10219
rect 35980 10134 36020 10219
rect 35883 10100 35925 10109
rect 35883 10060 35884 10100
rect 35924 10060 35925 10100
rect 35883 10051 35925 10060
rect 35691 10016 35733 10025
rect 35691 9976 35692 10016
rect 35732 9976 35733 10016
rect 35691 9967 35733 9976
rect 34539 9932 34581 9941
rect 34539 9892 34540 9932
rect 34580 9892 34581 9932
rect 34539 9883 34581 9892
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 34540 9680 34580 9883
rect 35692 9882 35732 9967
rect 34540 9631 34580 9640
rect 35115 9680 35157 9689
rect 35115 9640 35116 9680
rect 35156 9640 35157 9680
rect 35115 9631 35157 9640
rect 32235 9428 32277 9437
rect 32235 9388 32236 9428
rect 32276 9388 32277 9428
rect 32235 9379 32277 9388
rect 34444 9428 34484 9437
rect 33387 9176 33429 9185
rect 33387 9136 33388 9176
rect 33428 9136 33429 9176
rect 33387 9127 33429 9136
rect 32619 8924 32661 8933
rect 32619 8884 32620 8924
rect 32660 8884 32661 8924
rect 32619 8875 32661 8884
rect 32332 8756 32372 8765
rect 32140 8716 32332 8756
rect 32139 8420 32181 8429
rect 32139 8380 32140 8420
rect 32180 8380 32181 8420
rect 32139 8371 32181 8380
rect 32140 8009 32180 8371
rect 32139 8000 32181 8009
rect 32139 7960 32140 8000
rect 32180 7960 32181 8000
rect 32139 7951 32181 7960
rect 31947 7916 31989 7925
rect 31947 7876 31948 7916
rect 31988 7876 31989 7916
rect 31947 7867 31989 7876
rect 32140 7916 32180 7951
rect 31948 7782 31988 7867
rect 32140 7865 32180 7876
rect 32043 7832 32085 7841
rect 32043 7792 32044 7832
rect 32084 7792 32085 7832
rect 32043 7783 32085 7792
rect 32044 7698 32084 7783
rect 32236 7580 32276 8716
rect 32332 8707 32372 8716
rect 32523 8588 32565 8597
rect 32523 8548 32524 8588
rect 32564 8548 32565 8588
rect 32523 8539 32565 8548
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 32332 7916 32372 7927
rect 32332 7841 32372 7876
rect 32428 7866 32468 7951
rect 32524 7916 32564 8539
rect 32524 7867 32564 7876
rect 32331 7832 32373 7841
rect 32331 7792 32332 7832
rect 32372 7792 32373 7832
rect 32331 7783 32373 7792
rect 32620 7748 32660 8875
rect 32907 8336 32949 8345
rect 32907 8296 32908 8336
rect 32948 8296 32949 8336
rect 32907 8287 32949 8296
rect 32908 8177 32948 8287
rect 32907 8168 32949 8177
rect 32907 8128 32908 8168
rect 32948 8128 32949 8168
rect 32907 8119 32949 8128
rect 32716 7916 32756 7927
rect 32716 7841 32756 7876
rect 32811 7916 32853 7925
rect 32811 7876 32812 7916
rect 32852 7876 32853 7916
rect 32811 7867 32853 7876
rect 32908 7916 32948 8119
rect 32908 7867 32948 7876
rect 33100 7916 33140 7927
rect 32715 7832 32757 7841
rect 32715 7792 32716 7832
rect 32756 7792 32757 7832
rect 32715 7783 32757 7792
rect 31756 7372 31892 7412
rect 32044 7540 32276 7580
rect 32524 7708 32660 7748
rect 31180 7244 31220 7253
rect 31180 7001 31220 7204
rect 31660 7244 31700 7255
rect 31660 7169 31700 7204
rect 31659 7160 31701 7169
rect 31659 7120 31660 7160
rect 31700 7120 31701 7160
rect 31659 7111 31701 7120
rect 30987 6992 31029 7001
rect 30987 6952 30988 6992
rect 31028 6952 31029 6992
rect 30987 6943 31029 6952
rect 31179 6992 31221 7001
rect 31179 6952 31180 6992
rect 31220 6952 31221 6992
rect 31179 6943 31221 6952
rect 30891 5900 30933 5909
rect 30891 5860 30892 5900
rect 30932 5860 30933 5900
rect 30891 5851 30933 5860
rect 31083 5900 31125 5909
rect 31083 5860 31084 5900
rect 31124 5860 31125 5900
rect 31083 5851 31125 5860
rect 30795 5732 30837 5741
rect 30795 5692 30796 5732
rect 30836 5692 30837 5732
rect 30795 5683 30837 5692
rect 30796 5598 30836 5683
rect 30699 5144 30741 5153
rect 30699 5104 30700 5144
rect 30740 5104 30741 5144
rect 30699 5095 30741 5104
rect 30700 4985 30740 5016
rect 30699 4976 30741 4985
rect 30699 4936 30700 4976
rect 30740 4936 30741 4976
rect 30699 4927 30741 4936
rect 30700 4892 30740 4927
rect 30892 4901 30932 5851
rect 31084 5732 31124 5851
rect 31084 5683 31124 5692
rect 31180 5564 31220 6943
rect 31659 6824 31701 6833
rect 31659 6784 31660 6824
rect 31700 6784 31701 6824
rect 31659 6775 31701 6784
rect 31563 6740 31605 6749
rect 31563 6700 31564 6740
rect 31604 6700 31605 6740
rect 31563 6691 31605 6700
rect 31564 6488 31604 6691
rect 31660 6665 31700 6775
rect 31659 6656 31701 6665
rect 31659 6616 31660 6656
rect 31700 6616 31701 6656
rect 31659 6607 31701 6616
rect 31468 6448 31604 6488
rect 31468 6404 31508 6448
rect 31468 6355 31508 6364
rect 31660 6404 31700 6413
rect 31660 6329 31700 6364
rect 31659 6320 31701 6329
rect 31659 6280 31660 6320
rect 31700 6280 31701 6320
rect 31659 6271 31701 6280
rect 31467 6236 31509 6245
rect 31467 6196 31468 6236
rect 31508 6196 31509 6236
rect 31467 6187 31509 6196
rect 31564 6236 31604 6245
rect 31275 5816 31317 5825
rect 31275 5776 31276 5816
rect 31316 5776 31317 5816
rect 31275 5767 31317 5776
rect 31276 5732 31316 5767
rect 31276 5681 31316 5692
rect 31468 5732 31508 6187
rect 31180 5524 31316 5564
rect 31083 5480 31125 5489
rect 31083 5440 31084 5480
rect 31124 5440 31125 5480
rect 31083 5431 31125 5440
rect 31084 5346 31124 5431
rect 31180 5060 31220 5069
rect 30988 5020 31180 5060
rect 30700 4397 30740 4852
rect 30891 4892 30933 4901
rect 30891 4852 30892 4892
rect 30932 4852 30933 4892
rect 30891 4843 30933 4852
rect 30795 4724 30837 4733
rect 30795 4684 30796 4724
rect 30836 4684 30837 4724
rect 30795 4675 30837 4684
rect 30796 4590 30836 4675
rect 30795 4472 30837 4481
rect 30795 4432 30796 4472
rect 30836 4432 30837 4472
rect 30795 4423 30837 4432
rect 30699 4388 30741 4397
rect 30699 4348 30700 4388
rect 30740 4348 30741 4388
rect 30699 4339 30741 4348
rect 30700 4220 30740 4229
rect 30604 4180 30700 4220
rect 30508 3893 30548 4180
rect 30700 4171 30740 4180
rect 30507 3884 30549 3893
rect 30507 3844 30508 3884
rect 30548 3844 30549 3884
rect 30507 3835 30549 3844
rect 30508 3725 30548 3835
rect 30507 3716 30549 3725
rect 30507 3676 30508 3716
rect 30548 3676 30549 3716
rect 30507 3667 30549 3676
rect 30412 3415 30452 3424
rect 30796 3464 30836 4423
rect 30892 4229 30932 4843
rect 30891 4220 30933 4229
rect 30891 4180 30892 4220
rect 30932 4180 30933 4220
rect 30891 4171 30933 4180
rect 30891 4052 30933 4061
rect 30891 4012 30892 4052
rect 30932 4012 30933 4052
rect 30891 4003 30933 4012
rect 30892 3918 30932 4003
rect 30988 3632 31028 5020
rect 31180 5011 31220 5020
rect 31180 4892 31220 4901
rect 31276 4892 31316 5524
rect 31468 4905 31508 5692
rect 31220 4852 31316 4892
rect 31372 4892 31508 4905
rect 31564 4901 31604 6196
rect 31660 5741 31700 6271
rect 31659 5732 31701 5741
rect 31659 5692 31660 5732
rect 31700 5692 31701 5732
rect 31659 5683 31701 5692
rect 31659 5480 31701 5489
rect 31659 5440 31660 5480
rect 31700 5440 31701 5480
rect 31659 5431 31701 5440
rect 31660 5346 31700 5431
rect 31660 5069 31700 5154
rect 31659 5060 31701 5069
rect 31756 5060 31796 7372
rect 31860 7244 31900 7252
rect 31947 7244 31989 7253
rect 31860 7243 31948 7244
rect 31900 7204 31948 7243
rect 31988 7204 31989 7244
rect 31860 7194 31900 7203
rect 31947 7195 31989 7204
rect 31852 7076 31892 7085
rect 32044 7076 32084 7540
rect 32332 7253 32372 7338
rect 32139 7244 32181 7253
rect 32331 7244 32373 7253
rect 32139 7204 32140 7244
rect 32180 7204 32276 7244
rect 32139 7195 32181 7204
rect 31892 7036 32084 7076
rect 32236 7076 32276 7204
rect 32331 7204 32332 7244
rect 32372 7204 32373 7244
rect 32331 7195 32373 7204
rect 32331 7076 32373 7085
rect 32236 7036 32332 7076
rect 32372 7036 32373 7076
rect 31852 7027 31892 7036
rect 32331 7027 32373 7036
rect 32139 6992 32181 7001
rect 32139 6952 32140 6992
rect 32180 6952 32181 6992
rect 32139 6943 32181 6952
rect 32043 6908 32085 6917
rect 32043 6868 32044 6908
rect 32084 6868 32085 6908
rect 32043 6859 32085 6868
rect 31851 6656 31893 6665
rect 31851 6616 31852 6656
rect 31892 6616 31893 6656
rect 32044 6656 32084 6859
rect 32140 6858 32180 6943
rect 32332 6942 32372 7027
rect 32235 6824 32277 6833
rect 32235 6784 32236 6824
rect 32276 6784 32277 6824
rect 32235 6775 32277 6784
rect 32044 6616 32180 6656
rect 31851 6607 31893 6616
rect 31852 6404 31892 6607
rect 32044 6413 32084 6498
rect 31852 6355 31892 6364
rect 32043 6404 32085 6413
rect 32043 6364 32044 6404
rect 32084 6364 32085 6404
rect 32043 6355 32085 6364
rect 32140 6320 32180 6616
rect 32236 6581 32276 6775
rect 32235 6572 32277 6581
rect 32235 6532 32236 6572
rect 32276 6532 32277 6572
rect 32235 6523 32277 6532
rect 32236 6417 32276 6523
rect 32236 6368 32276 6377
rect 32428 6404 32468 6413
rect 32331 6320 32373 6329
rect 32140 6280 32276 6320
rect 31948 6236 31988 6245
rect 31988 6196 32180 6236
rect 31948 6187 31988 6196
rect 31851 6068 31893 6077
rect 31851 6028 31852 6068
rect 31892 6028 31893 6068
rect 31851 6019 31893 6028
rect 31852 5825 31892 6019
rect 31851 5816 31893 5825
rect 31851 5776 31852 5816
rect 31892 5776 31893 5816
rect 31851 5767 31893 5776
rect 31852 5732 31892 5767
rect 32044 5741 32084 5826
rect 31852 5681 31892 5692
rect 32043 5732 32085 5741
rect 32043 5692 32044 5732
rect 32084 5692 32085 5732
rect 32043 5683 32085 5692
rect 31947 5480 31989 5489
rect 31947 5440 31948 5480
rect 31988 5440 31989 5480
rect 31947 5431 31989 5440
rect 32044 5480 32084 5489
rect 31851 5396 31893 5405
rect 31851 5356 31852 5396
rect 31892 5356 31893 5396
rect 31851 5347 31893 5356
rect 31659 5020 31660 5060
rect 31700 5020 31701 5060
rect 31659 5011 31701 5020
rect 31755 5020 31796 5060
rect 31755 4976 31795 5020
rect 31755 4936 31796 4976
rect 31412 4865 31508 4892
rect 31563 4892 31605 4901
rect 31180 4843 31220 4852
rect 31372 4843 31412 4852
rect 31563 4852 31564 4892
rect 31604 4852 31605 4892
rect 31563 4843 31605 4852
rect 31660 4881 31700 4890
rect 31563 4724 31605 4733
rect 31563 4684 31564 4724
rect 31604 4684 31605 4724
rect 31563 4675 31605 4684
rect 31083 4472 31125 4481
rect 31083 4432 31084 4472
rect 31124 4432 31125 4472
rect 31083 4423 31125 4432
rect 31084 4313 31124 4423
rect 31083 4304 31125 4313
rect 31083 4264 31084 4304
rect 31124 4264 31125 4304
rect 31083 4255 31125 4264
rect 31467 4304 31509 4313
rect 31467 4264 31468 4304
rect 31508 4264 31509 4304
rect 31467 4255 31509 4264
rect 31084 4220 31124 4255
rect 31084 4169 31124 4180
rect 31275 4220 31317 4229
rect 31275 4180 31276 4220
rect 31316 4180 31317 4220
rect 31275 4171 31317 4180
rect 30796 3415 30836 3424
rect 30892 3592 31028 3632
rect 31180 4136 31220 4145
rect 30219 3212 30261 3221
rect 30219 3172 30220 3212
rect 30260 3172 30261 3212
rect 30219 3163 30261 3172
rect 30604 3212 30644 3221
rect 30220 3078 30260 3163
rect 30315 3128 30357 3137
rect 30315 3088 30316 3128
rect 30356 3088 30357 3128
rect 30315 3079 30357 3088
rect 30219 1784 30261 1793
rect 30219 1744 30220 1784
rect 30260 1744 30261 1784
rect 30219 1735 30261 1744
rect 30220 1289 30260 1735
rect 30219 1280 30261 1289
rect 30219 1240 30220 1280
rect 30260 1240 30261 1280
rect 30219 1231 30261 1240
rect 30123 1112 30165 1121
rect 30316 1112 30356 3079
rect 30604 2885 30644 3172
rect 30603 2876 30645 2885
rect 30603 2836 30604 2876
rect 30644 2836 30645 2876
rect 30603 2827 30645 2836
rect 30892 2297 30932 3592
rect 31180 3464 31220 4096
rect 31276 4086 31316 4171
rect 31468 4136 31508 4255
rect 31468 4087 31508 4096
rect 31275 3968 31317 3977
rect 31275 3928 31276 3968
rect 31316 3928 31317 3968
rect 31275 3919 31317 3928
rect 31180 3415 31220 3424
rect 30988 3212 31028 3221
rect 30891 2288 30933 2297
rect 30891 2248 30892 2288
rect 30932 2248 30933 2288
rect 30891 2239 30933 2248
rect 30988 1625 31028 3172
rect 31276 3137 31316 3919
rect 31564 3464 31604 4675
rect 31660 4229 31700 4841
rect 31659 4220 31701 4229
rect 31659 4180 31660 4220
rect 31700 4180 31701 4220
rect 31659 4171 31701 4180
rect 31564 3415 31604 3424
rect 31660 3968 31700 3977
rect 31372 3212 31412 3221
rect 31275 3128 31317 3137
rect 31275 3088 31276 3128
rect 31316 3088 31317 3128
rect 31275 3079 31317 3088
rect 31275 2792 31317 2801
rect 31275 2752 31276 2792
rect 31316 2752 31317 2792
rect 31275 2743 31317 2752
rect 31179 2708 31221 2717
rect 31179 2668 31180 2708
rect 31220 2668 31221 2708
rect 31179 2659 31221 2668
rect 30987 1616 31029 1625
rect 30987 1576 30988 1616
rect 31028 1576 31029 1616
rect 30987 1567 31029 1576
rect 30411 1196 30453 1205
rect 30411 1156 30412 1196
rect 30452 1156 30453 1196
rect 30411 1147 30453 1156
rect 30123 1072 30124 1112
rect 30164 1072 30165 1112
rect 30123 1063 30165 1072
rect 30220 1072 30356 1112
rect 30220 80 30260 1072
rect 30412 80 30452 1147
rect 30987 1112 31029 1121
rect 30987 1072 30988 1112
rect 31028 1072 31029 1112
rect 30987 1063 31029 1072
rect 30795 1028 30837 1037
rect 30795 988 30796 1028
rect 30836 988 30837 1028
rect 30795 979 30837 988
rect 30603 944 30645 953
rect 30603 904 30604 944
rect 30644 904 30645 944
rect 30603 895 30645 904
rect 30604 80 30644 895
rect 30796 80 30836 979
rect 30988 80 31028 1063
rect 31180 80 31220 2659
rect 31276 1028 31316 2743
rect 31372 1205 31412 3172
rect 31563 3212 31605 3221
rect 31563 3172 31564 3212
rect 31604 3172 31605 3212
rect 31563 3163 31605 3172
rect 31564 1616 31604 3163
rect 31660 2045 31700 3928
rect 31756 3389 31796 4936
rect 31852 4892 31892 5347
rect 31852 4843 31892 4852
rect 31852 4136 31892 4147
rect 31852 4061 31892 4096
rect 31851 4052 31893 4061
rect 31851 4012 31852 4052
rect 31892 4012 31893 4052
rect 31851 4003 31893 4012
rect 31948 3641 31988 5431
rect 32044 4145 32084 5440
rect 32140 4808 32180 6196
rect 32236 5732 32276 6280
rect 32331 6280 32332 6320
rect 32372 6280 32373 6320
rect 32331 6271 32373 6280
rect 32332 6186 32372 6271
rect 32331 5984 32373 5993
rect 32331 5944 32332 5984
rect 32372 5944 32373 5984
rect 32331 5935 32373 5944
rect 32236 5683 32276 5692
rect 32332 5573 32372 5935
rect 32428 5741 32468 6364
rect 32524 5984 32564 7708
rect 32620 7244 32660 7253
rect 32716 7244 32756 7783
rect 32812 7782 32852 7867
rect 33100 7841 33140 7876
rect 33195 7916 33237 7925
rect 33195 7876 33196 7916
rect 33236 7876 33237 7916
rect 33195 7867 33237 7876
rect 33292 7916 33332 7925
rect 33099 7832 33141 7841
rect 33099 7792 33100 7832
rect 33140 7792 33141 7832
rect 33099 7783 33141 7792
rect 33196 7782 33236 7867
rect 33292 7673 33332 7876
rect 33291 7664 33333 7673
rect 33291 7624 33292 7664
rect 33332 7624 33333 7664
rect 33291 7615 33333 7624
rect 32811 7580 32853 7589
rect 32811 7540 32812 7580
rect 32852 7540 32853 7580
rect 32811 7531 32853 7540
rect 32660 7204 32756 7244
rect 32812 7244 32852 7531
rect 33291 7412 33333 7421
rect 33291 7372 33292 7412
rect 33332 7372 33333 7412
rect 33291 7363 33333 7372
rect 32620 7195 32660 7204
rect 32812 7195 32852 7204
rect 33195 7160 33237 7169
rect 33195 7120 33196 7160
rect 33236 7120 33237 7160
rect 33195 7111 33237 7120
rect 32716 6992 32756 7001
rect 32619 6404 32661 6413
rect 32619 6364 32620 6404
rect 32660 6364 32661 6404
rect 32619 6355 32661 6364
rect 32620 6270 32660 6355
rect 32716 6161 32756 6952
rect 32812 6572 32852 6581
rect 32852 6532 32948 6572
rect 32812 6523 32852 6532
rect 32812 6404 32852 6413
rect 32715 6152 32757 6161
rect 32715 6112 32716 6152
rect 32756 6112 32757 6152
rect 32715 6103 32757 6112
rect 32524 5944 32756 5984
rect 32427 5732 32469 5741
rect 32427 5692 32428 5732
rect 32468 5692 32469 5732
rect 32427 5683 32469 5692
rect 32620 5732 32660 5741
rect 32523 5648 32565 5657
rect 32523 5608 32524 5648
rect 32564 5608 32565 5648
rect 32523 5599 32565 5608
rect 32331 5564 32373 5573
rect 32331 5524 32332 5564
rect 32372 5524 32373 5564
rect 32331 5515 32373 5524
rect 32235 5480 32277 5489
rect 32235 5440 32236 5480
rect 32276 5440 32277 5480
rect 32235 5431 32277 5440
rect 32427 5480 32469 5489
rect 32427 5440 32428 5480
rect 32468 5440 32469 5480
rect 32427 5431 32469 5440
rect 32236 4976 32276 5431
rect 32428 5346 32468 5431
rect 32236 4927 32276 4936
rect 32524 4808 32564 5599
rect 32620 5573 32660 5692
rect 32619 5564 32661 5573
rect 32619 5524 32620 5564
rect 32660 5524 32661 5564
rect 32619 5515 32661 5524
rect 32620 4976 32660 4985
rect 32716 4976 32756 5944
rect 32812 5741 32852 6364
rect 32811 5732 32853 5741
rect 32811 5692 32812 5732
rect 32852 5692 32853 5732
rect 32811 5683 32853 5692
rect 32812 5480 32852 5489
rect 32812 5321 32852 5440
rect 32811 5312 32853 5321
rect 32811 5272 32812 5312
rect 32852 5272 32853 5312
rect 32811 5263 32853 5272
rect 32660 4936 32756 4976
rect 32620 4927 32660 4936
rect 32715 4808 32757 4817
rect 32140 4768 32372 4808
rect 32524 4768 32660 4808
rect 32235 4304 32277 4313
rect 32235 4264 32236 4304
rect 32276 4264 32277 4304
rect 32235 4255 32277 4264
rect 32043 4136 32085 4145
rect 32043 4096 32044 4136
rect 32084 4096 32085 4136
rect 32043 4087 32085 4096
rect 32236 4136 32276 4255
rect 32236 4087 32276 4096
rect 32044 3968 32084 3977
rect 32084 3928 32276 3968
rect 32044 3919 32084 3928
rect 31947 3632 31989 3641
rect 31947 3592 31948 3632
rect 31988 3592 31989 3632
rect 31947 3583 31989 3592
rect 31947 3464 31989 3473
rect 31947 3424 31948 3464
rect 31988 3424 31989 3464
rect 31947 3415 31989 3424
rect 31755 3380 31797 3389
rect 31755 3340 31756 3380
rect 31796 3340 31797 3380
rect 31755 3331 31797 3340
rect 31948 3330 31988 3415
rect 31756 3212 31796 3221
rect 31756 2801 31796 3172
rect 32140 3212 32180 3221
rect 32140 2969 32180 3172
rect 32139 2960 32181 2969
rect 32139 2920 32140 2960
rect 32180 2920 32181 2960
rect 32139 2911 32181 2920
rect 32043 2876 32085 2885
rect 32043 2836 32044 2876
rect 32084 2836 32085 2876
rect 32043 2827 32085 2836
rect 31755 2792 31797 2801
rect 31755 2752 31756 2792
rect 31796 2752 31797 2792
rect 31755 2743 31797 2752
rect 31659 2036 31701 2045
rect 31659 1996 31660 2036
rect 31700 1996 31701 2036
rect 31659 1987 31701 1996
rect 32044 1616 32084 2827
rect 31564 1576 31988 1616
rect 32044 1576 32180 1616
rect 31755 1364 31797 1373
rect 31755 1324 31756 1364
rect 31796 1324 31797 1364
rect 31755 1315 31797 1324
rect 31563 1280 31605 1289
rect 31563 1240 31564 1280
rect 31604 1240 31605 1280
rect 31563 1231 31605 1240
rect 31371 1196 31413 1205
rect 31371 1156 31372 1196
rect 31412 1156 31413 1196
rect 31371 1147 31413 1156
rect 31276 988 31412 1028
rect 31372 80 31412 988
rect 31564 80 31604 1231
rect 31756 80 31796 1315
rect 31948 80 31988 1576
rect 32140 80 32180 1576
rect 32236 785 32276 3928
rect 32332 3464 32372 4768
rect 32428 4724 32468 4733
rect 32468 4684 32564 4724
rect 32428 4675 32468 4684
rect 32332 3415 32372 3424
rect 32428 3968 32468 3977
rect 32331 2036 32373 2045
rect 32331 1996 32332 2036
rect 32372 1996 32373 2036
rect 32331 1987 32373 1996
rect 32235 776 32277 785
rect 32235 736 32236 776
rect 32276 736 32277 776
rect 32235 727 32277 736
rect 32332 80 32372 1987
rect 32428 1289 32468 3928
rect 32524 3632 32564 4684
rect 32620 4136 32660 4768
rect 32715 4768 32716 4808
rect 32756 4768 32757 4808
rect 32908 4808 32948 6532
rect 33196 6497 33236 7111
rect 33292 7085 33332 7363
rect 33291 7076 33333 7085
rect 33291 7036 33292 7076
rect 33332 7036 33333 7076
rect 33291 7027 33333 7036
rect 33003 6488 33045 6497
rect 33003 6448 33004 6488
rect 33044 6448 33045 6488
rect 33003 6439 33045 6448
rect 33195 6488 33237 6497
rect 33195 6448 33196 6488
rect 33236 6448 33237 6488
rect 33195 6439 33237 6448
rect 33004 6236 33044 6439
rect 33099 6404 33141 6413
rect 33099 6364 33100 6404
rect 33140 6364 33141 6404
rect 33099 6355 33141 6364
rect 33196 6404 33236 6439
rect 33004 6187 33044 6196
rect 33100 5909 33140 6355
rect 33196 6354 33236 6364
rect 33292 6404 33332 7027
rect 33292 6355 33332 6364
rect 33388 5993 33428 9127
rect 33483 9008 33525 9017
rect 33483 8968 33484 9008
rect 33524 8968 33525 9008
rect 33483 8959 33525 8968
rect 33387 5984 33429 5993
rect 33387 5944 33388 5984
rect 33428 5944 33429 5984
rect 33387 5935 33429 5944
rect 33099 5900 33141 5909
rect 33099 5860 33100 5900
rect 33140 5860 33141 5900
rect 33099 5851 33141 5860
rect 33291 5480 33333 5489
rect 33291 5440 33292 5480
rect 33332 5440 33333 5480
rect 33484 5480 33524 8959
rect 33964 8756 34004 8765
rect 33772 8716 33964 8756
rect 33675 8672 33717 8681
rect 33675 8632 33676 8672
rect 33716 8632 33717 8672
rect 33675 8623 33717 8632
rect 33579 7916 33621 7925
rect 33579 7876 33580 7916
rect 33620 7876 33621 7916
rect 33579 7867 33621 7876
rect 33580 7782 33620 7867
rect 33676 7589 33716 8623
rect 33772 8252 33812 8716
rect 33964 8707 34004 8716
rect 34155 8756 34197 8765
rect 34155 8716 34156 8756
rect 34196 8716 34197 8756
rect 34155 8707 34197 8716
rect 34347 8756 34389 8765
rect 34444 8756 34484 9388
rect 34636 9428 34676 9437
rect 34828 9428 34868 9437
rect 34347 8716 34348 8756
rect 34388 8716 34484 8756
rect 34540 8756 34580 8765
rect 34347 8707 34389 8716
rect 34060 8672 34100 8681
rect 34060 8513 34100 8632
rect 34156 8622 34196 8707
rect 34059 8504 34101 8513
rect 34059 8464 34060 8504
rect 34100 8464 34101 8504
rect 34059 8455 34101 8464
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 33772 8212 33883 8252
rect 33843 8168 33883 8212
rect 33843 8128 33908 8168
rect 33771 8084 33813 8093
rect 33771 8044 33772 8084
rect 33812 8044 33813 8084
rect 33771 8035 33813 8044
rect 33772 7916 33812 8035
rect 33772 7867 33812 7876
rect 33868 7841 33908 8128
rect 34348 7916 34388 8707
rect 34540 8597 34580 8716
rect 34539 8588 34581 8597
rect 34539 8548 34540 8588
rect 34580 8548 34581 8588
rect 34539 8539 34581 8548
rect 34444 8504 34484 8513
rect 34444 8345 34484 8464
rect 34443 8336 34485 8345
rect 34443 8296 34444 8336
rect 34484 8296 34485 8336
rect 34443 8287 34485 8296
rect 34636 8177 34676 9388
rect 34732 9388 34828 9428
rect 34732 8765 34772 9388
rect 34828 9379 34868 9388
rect 35020 9428 35060 9437
rect 34923 9344 34965 9353
rect 34923 9304 34924 9344
rect 34964 9304 34965 9344
rect 34923 9295 34965 9304
rect 34827 9260 34869 9269
rect 34827 9220 34828 9260
rect 34868 9220 34869 9260
rect 34827 9211 34869 9220
rect 34828 9092 34868 9211
rect 34924 9210 34964 9295
rect 34828 9052 34964 9092
rect 34827 8924 34869 8933
rect 34827 8884 34828 8924
rect 34868 8884 34869 8924
rect 34827 8875 34869 8884
rect 34828 8840 34868 8875
rect 34828 8789 34868 8800
rect 34731 8756 34773 8765
rect 34731 8716 34732 8756
rect 34772 8716 34773 8756
rect 34731 8707 34773 8716
rect 34924 8756 34964 9052
rect 34732 8622 34772 8707
rect 34827 8252 34869 8261
rect 34924 8252 34964 8716
rect 35020 8429 35060 9388
rect 35116 9269 35156 9631
rect 35115 9260 35157 9269
rect 35115 9220 35116 9260
rect 35156 9220 35157 9260
rect 35115 9211 35157 9220
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35691 8840 35733 8849
rect 35691 8800 35692 8840
rect 35732 8800 35733 8840
rect 35691 8791 35733 8800
rect 35115 8756 35157 8765
rect 35115 8716 35116 8756
rect 35156 8716 35157 8756
rect 35115 8707 35157 8716
rect 35308 8756 35348 8767
rect 35116 8622 35156 8707
rect 35308 8681 35348 8716
rect 35499 8756 35541 8765
rect 35499 8716 35500 8756
rect 35540 8716 35541 8756
rect 35499 8707 35541 8716
rect 35692 8756 35732 8791
rect 35307 8672 35349 8681
rect 35307 8632 35308 8672
rect 35348 8632 35349 8672
rect 35307 8623 35349 8632
rect 35500 8622 35540 8707
rect 35692 8681 35732 8716
rect 35691 8672 35733 8681
rect 35691 8632 35692 8672
rect 35732 8632 35733 8672
rect 35691 8623 35733 8632
rect 35692 8592 35732 8623
rect 35212 8504 35252 8513
rect 35595 8504 35637 8513
rect 35252 8464 35540 8504
rect 35212 8455 35252 8464
rect 35019 8420 35061 8429
rect 35019 8380 35020 8420
rect 35060 8380 35061 8420
rect 35019 8371 35061 8380
rect 35020 8261 35060 8371
rect 34827 8212 34828 8252
rect 34868 8212 34964 8252
rect 35019 8252 35061 8261
rect 35019 8212 35020 8252
rect 35060 8212 35061 8252
rect 34827 8203 34869 8212
rect 35019 8203 35061 8212
rect 34635 8168 34677 8177
rect 34635 8128 34636 8168
rect 34676 8128 34677 8168
rect 34635 8119 34677 8128
rect 35307 8168 35349 8177
rect 35307 8128 35308 8168
rect 35348 8128 35349 8168
rect 35307 8119 35349 8128
rect 34923 8000 34965 8009
rect 34923 7960 34924 8000
rect 34964 7960 34965 8000
rect 34923 7951 34965 7960
rect 35308 8000 35348 8119
rect 35308 7951 35348 7960
rect 34443 7916 34485 7925
rect 34348 7876 34444 7916
rect 34484 7876 34485 7916
rect 34443 7867 34485 7876
rect 34636 7916 34676 7925
rect 33867 7832 33909 7841
rect 33867 7792 33868 7832
rect 33908 7792 33909 7832
rect 33867 7783 33909 7792
rect 33675 7580 33717 7589
rect 33675 7540 33676 7580
rect 33716 7540 33717 7580
rect 33675 7531 33717 7540
rect 33868 7421 33908 7783
rect 34444 7782 34484 7867
rect 34540 7832 34580 7841
rect 33867 7412 33909 7421
rect 33867 7372 33868 7412
rect 33908 7372 33909 7412
rect 33867 7363 33909 7372
rect 33867 7244 33909 7253
rect 33867 7204 33868 7244
rect 33908 7204 33909 7244
rect 33867 7195 33909 7204
rect 34059 7244 34101 7253
rect 34059 7204 34060 7244
rect 34100 7204 34101 7244
rect 34059 7195 34101 7204
rect 34252 7244 34292 7255
rect 33868 7110 33908 7195
rect 33964 7160 34004 7169
rect 33964 7001 34004 7120
rect 34060 7110 34100 7195
rect 34252 7169 34292 7204
rect 34347 7244 34389 7253
rect 34444 7244 34484 7253
rect 34347 7204 34348 7244
rect 34388 7204 34444 7244
rect 34347 7195 34389 7204
rect 34444 7195 34484 7204
rect 34251 7160 34293 7169
rect 34251 7120 34252 7160
rect 34292 7120 34293 7160
rect 34251 7111 34293 7120
rect 33963 6992 34005 7001
rect 33963 6952 33964 6992
rect 34004 6952 34005 6992
rect 33963 6943 34005 6952
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 33675 6740 33717 6749
rect 33675 6700 33676 6740
rect 33716 6700 33717 6740
rect 33675 6691 33717 6700
rect 33676 6404 33716 6691
rect 34059 6656 34101 6665
rect 34059 6616 34060 6656
rect 34100 6616 34101 6656
rect 34059 6607 34101 6616
rect 33676 6355 33716 6364
rect 33867 6404 33909 6413
rect 33867 6364 33868 6404
rect 33908 6364 33909 6404
rect 33867 6355 33909 6364
rect 34060 6404 34100 6607
rect 34348 6413 34388 7195
rect 34540 7085 34580 7792
rect 34636 7757 34676 7876
rect 34827 7916 34869 7925
rect 34827 7876 34828 7916
rect 34868 7876 34869 7916
rect 34827 7867 34869 7876
rect 34828 7782 34868 7867
rect 34924 7866 34964 7951
rect 35020 7916 35060 7925
rect 35020 7841 35060 7876
rect 35019 7832 35061 7841
rect 35019 7792 35020 7832
rect 35060 7792 35061 7832
rect 35019 7783 35061 7792
rect 34635 7748 34677 7757
rect 34635 7708 34636 7748
rect 34676 7708 34677 7748
rect 34635 7699 34677 7708
rect 34636 7421 34676 7699
rect 35020 7673 35060 7783
rect 35500 7748 35540 8464
rect 35595 8464 35596 8504
rect 35636 8464 35637 8504
rect 35595 8455 35637 8464
rect 35596 8370 35636 8455
rect 35884 8252 35924 10051
rect 36268 9437 36308 10228
rect 36363 10219 36405 10228
rect 36556 10268 36596 10279
rect 36364 10134 36404 10219
rect 36556 10193 36596 10228
rect 36555 10184 36597 10193
rect 36555 10144 36556 10184
rect 36596 10144 36597 10184
rect 36555 10135 36597 10144
rect 36652 9857 36692 10396
rect 36748 10277 36788 10900
rect 36844 10891 36884 10900
rect 37036 10940 37076 10951
rect 39052 10940 39092 14920
rect 49899 11444 49941 11453
rect 49899 11404 49900 11444
rect 49940 11404 49941 11444
rect 49899 11395 49941 11404
rect 49048 11360 49416 11369
rect 49088 11320 49130 11360
rect 49170 11320 49212 11360
rect 49252 11320 49294 11360
rect 49334 11320 49376 11360
rect 49048 11311 49416 11320
rect 39148 10940 39188 10949
rect 39340 10940 39380 10949
rect 39052 10900 39148 10940
rect 37036 10865 37076 10900
rect 39148 10891 39188 10900
rect 39244 10900 39340 10940
rect 36940 10856 36980 10865
rect 36940 10688 36980 10816
rect 37035 10856 37077 10865
rect 37035 10816 37036 10856
rect 37076 10816 37077 10856
rect 37035 10807 37077 10816
rect 37419 10856 37461 10865
rect 37419 10816 37420 10856
rect 37460 10816 37461 10856
rect 37419 10807 37461 10816
rect 37995 10856 38037 10865
rect 37995 10816 37996 10856
rect 38036 10816 38037 10856
rect 37995 10807 38037 10816
rect 36940 10648 37268 10688
rect 36939 10352 36981 10361
rect 36939 10312 36940 10352
rect 36980 10312 36981 10352
rect 36939 10303 36981 10312
rect 36747 10268 36789 10277
rect 36747 10228 36748 10268
rect 36788 10228 36789 10268
rect 36747 10219 36789 10228
rect 36940 10268 36980 10303
rect 36748 10134 36788 10219
rect 36940 10193 36980 10228
rect 36939 10184 36981 10193
rect 36939 10144 36940 10184
rect 36980 10144 36981 10184
rect 36939 10135 36981 10144
rect 36940 10104 36980 10135
rect 36844 10016 36884 10025
rect 36884 9976 36980 10016
rect 36844 9967 36884 9976
rect 36651 9848 36693 9857
rect 36651 9808 36652 9848
rect 36692 9808 36693 9848
rect 36651 9799 36693 9808
rect 36843 9764 36885 9773
rect 36843 9724 36844 9764
rect 36884 9724 36885 9764
rect 36843 9715 36885 9724
rect 36363 9596 36405 9605
rect 36363 9556 36364 9596
rect 36404 9556 36405 9596
rect 36363 9547 36405 9556
rect 36364 9462 36404 9547
rect 36459 9512 36501 9521
rect 36459 9472 36460 9512
rect 36500 9472 36501 9512
rect 36459 9463 36501 9472
rect 36267 9428 36309 9437
rect 36267 9388 36268 9428
rect 36308 9388 36309 9428
rect 36267 9379 36309 9388
rect 36460 9428 36500 9463
rect 36268 9294 36308 9379
rect 36460 9377 36500 9388
rect 36651 9428 36693 9437
rect 36651 9388 36652 9428
rect 36692 9388 36693 9428
rect 36651 9379 36693 9388
rect 36844 9428 36884 9715
rect 36652 9294 36692 9379
rect 36844 9353 36884 9388
rect 36748 9344 36788 9353
rect 36748 8261 36788 9304
rect 36843 9344 36885 9353
rect 36843 9304 36844 9344
rect 36884 9304 36885 9344
rect 36843 9295 36885 9304
rect 36844 9264 36884 9295
rect 36940 9269 36980 9976
rect 37132 9428 37172 9437
rect 36939 9260 36981 9269
rect 36939 9220 36940 9260
rect 36980 9220 36981 9260
rect 36939 9211 36981 9220
rect 36843 9008 36885 9017
rect 36843 8968 36844 9008
rect 36884 8968 36885 9008
rect 36843 8959 36885 8968
rect 36844 8840 36884 8959
rect 36844 8800 36980 8840
rect 35692 8212 35924 8252
rect 36747 8252 36789 8261
rect 36747 8212 36748 8252
rect 36788 8212 36789 8252
rect 35500 7708 35636 7748
rect 35019 7664 35061 7673
rect 35019 7624 35020 7664
rect 35060 7624 35061 7664
rect 35019 7615 35061 7624
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 34635 7412 34677 7421
rect 34635 7372 34636 7412
rect 34676 7372 34677 7412
rect 34635 7363 34677 7372
rect 34635 7244 34677 7253
rect 34635 7204 34636 7244
rect 34676 7204 34677 7244
rect 34635 7195 34677 7204
rect 34539 7076 34581 7085
rect 34539 7036 34540 7076
rect 34580 7036 34581 7076
rect 34539 7027 34581 7036
rect 34444 6992 34484 7001
rect 34444 6833 34484 6952
rect 34443 6824 34485 6833
rect 34443 6784 34444 6824
rect 34484 6784 34485 6824
rect 34443 6775 34485 6784
rect 34636 6581 34676 7195
rect 34731 7160 34773 7169
rect 34731 7120 34732 7160
rect 34772 7120 34773 7160
rect 34731 7111 34773 7120
rect 34635 6572 34677 6581
rect 34444 6532 34636 6572
rect 34676 6532 34677 6572
rect 34060 6355 34100 6364
rect 34252 6404 34292 6413
rect 34347 6404 34389 6413
rect 34292 6364 34348 6404
rect 34388 6364 34389 6404
rect 34252 6355 34292 6364
rect 34347 6355 34389 6364
rect 34444 6404 34484 6532
rect 34635 6523 34677 6532
rect 34444 6355 34484 6364
rect 34636 6393 34676 6402
rect 33772 6245 33812 6330
rect 33868 6270 33908 6355
rect 34155 6320 34197 6329
rect 34155 6280 34156 6320
rect 34196 6280 34197 6320
rect 34155 6271 34197 6280
rect 33771 6236 33813 6245
rect 33771 6196 33772 6236
rect 33812 6196 33813 6236
rect 33771 6187 33813 6196
rect 34156 6186 34196 6271
rect 33771 5984 33813 5993
rect 33771 5944 33772 5984
rect 33812 5944 33813 5984
rect 33771 5935 33813 5944
rect 33772 5648 33812 5935
rect 34155 5900 34197 5909
rect 34155 5860 34156 5900
rect 34196 5860 34197 5900
rect 34155 5851 34197 5860
rect 34156 5732 34196 5851
rect 34348 5741 34388 6355
rect 34539 6236 34581 6245
rect 34539 6196 34540 6236
rect 34580 6196 34581 6236
rect 34539 6187 34581 6196
rect 34540 6102 34580 6187
rect 34539 5816 34581 5825
rect 34539 5776 34540 5816
rect 34580 5776 34581 5816
rect 34539 5767 34581 5776
rect 34156 5683 34196 5692
rect 34347 5732 34389 5741
rect 34347 5692 34348 5732
rect 34388 5692 34389 5732
rect 34347 5683 34389 5692
rect 34540 5732 34580 5767
rect 34636 5732 34676 6353
rect 34732 6077 34772 7111
rect 34827 6908 34869 6917
rect 34827 6868 34828 6908
rect 34868 6868 34869 6908
rect 34827 6859 34869 6868
rect 34828 6404 34868 6859
rect 35499 6572 35541 6581
rect 35499 6532 35500 6572
rect 35540 6532 35541 6572
rect 35499 6523 35541 6532
rect 35500 6438 35540 6523
rect 34828 6355 34868 6364
rect 35019 6404 35061 6413
rect 35019 6364 35020 6404
rect 35060 6364 35061 6404
rect 35019 6355 35061 6364
rect 35020 6270 35060 6355
rect 34924 6236 34964 6245
rect 34828 6196 34924 6236
rect 34731 6068 34773 6077
rect 34731 6028 34732 6068
rect 34772 6028 34773 6068
rect 34731 6019 34773 6028
rect 34732 5741 34772 5826
rect 34731 5732 34773 5741
rect 34636 5692 34732 5732
rect 34772 5692 34773 5732
rect 34540 5681 34580 5692
rect 34731 5683 34773 5692
rect 33772 5599 33812 5608
rect 33964 5489 34004 5574
rect 33963 5480 34005 5489
rect 33484 5440 33620 5480
rect 33291 5431 33333 5440
rect 33004 4985 33044 5070
rect 33003 4976 33045 4985
rect 33003 4936 33004 4976
rect 33044 4936 33045 4976
rect 33003 4927 33045 4936
rect 33292 4808 33332 5431
rect 33483 5312 33525 5321
rect 33483 5272 33484 5312
rect 33524 5272 33525 5312
rect 33483 5263 33525 5272
rect 33388 4985 33428 5070
rect 33387 4976 33429 4985
rect 33387 4936 33388 4976
rect 33428 4936 33429 4976
rect 33387 4927 33429 4936
rect 32908 4768 33044 4808
rect 33292 4768 33428 4808
rect 32715 4759 32757 4768
rect 32716 4313 32756 4759
rect 32812 4724 32852 4733
rect 32852 4684 32948 4724
rect 32812 4675 32852 4684
rect 32715 4304 32757 4313
rect 32715 4264 32716 4304
rect 32756 4264 32757 4304
rect 32715 4255 32757 4264
rect 32620 4087 32660 4096
rect 32715 4136 32757 4145
rect 32715 4096 32716 4136
rect 32756 4096 32757 4136
rect 32715 4087 32757 4096
rect 32524 3592 32660 3632
rect 32524 3212 32564 3221
rect 32524 2717 32564 3172
rect 32523 2708 32565 2717
rect 32523 2668 32524 2708
rect 32564 2668 32565 2708
rect 32523 2659 32565 2668
rect 32620 2372 32660 3592
rect 32716 3464 32756 4087
rect 32716 3415 32756 3424
rect 32812 3968 32852 3977
rect 32524 2332 32660 2372
rect 32427 1280 32469 1289
rect 32427 1240 32428 1280
rect 32468 1240 32469 1280
rect 32427 1231 32469 1240
rect 32524 80 32564 2332
rect 32812 1793 32852 3928
rect 32908 3632 32948 4684
rect 33004 4304 33044 4768
rect 33196 4724 33236 4733
rect 33236 4684 33332 4724
rect 33196 4675 33236 4684
rect 33004 4264 33140 4304
rect 33003 4136 33045 4145
rect 33003 4096 33004 4136
rect 33044 4096 33045 4136
rect 33003 4087 33045 4096
rect 33004 4002 33044 4087
rect 33100 3641 33140 4264
rect 33196 3968 33236 3977
rect 33099 3632 33141 3641
rect 32908 3592 33044 3632
rect 32908 3212 32948 3221
rect 32811 1784 32853 1793
rect 32811 1744 32812 1784
rect 32852 1744 32853 1784
rect 32811 1735 32853 1744
rect 32715 1616 32757 1625
rect 32715 1576 32716 1616
rect 32756 1576 32757 1616
rect 32715 1567 32757 1576
rect 32716 80 32756 1567
rect 32908 953 32948 3172
rect 33004 2372 33044 3592
rect 33099 3592 33100 3632
rect 33140 3592 33141 3632
rect 33099 3583 33141 3592
rect 33100 3464 33140 3475
rect 33100 3389 33140 3424
rect 33099 3380 33141 3389
rect 33099 3340 33100 3380
rect 33140 3340 33141 3380
rect 33099 3331 33141 3340
rect 33004 2332 33140 2372
rect 32907 944 32949 953
rect 32907 904 32908 944
rect 32948 904 32949 944
rect 32907 895 32949 904
rect 32907 776 32949 785
rect 32907 736 32908 776
rect 32948 736 32949 776
rect 32907 727 32949 736
rect 32908 80 32948 727
rect 33100 80 33140 2332
rect 33196 2045 33236 3928
rect 33292 3632 33332 4684
rect 33388 4136 33428 4768
rect 33388 4087 33428 4096
rect 33292 3592 33428 3632
rect 33292 3212 33332 3221
rect 33195 2036 33237 2045
rect 33195 1996 33196 2036
rect 33236 1996 33237 2036
rect 33195 1987 33237 1996
rect 33292 1364 33332 3172
rect 33388 2372 33428 3592
rect 33484 3464 33524 5263
rect 33580 4985 33620 5440
rect 33963 5440 33964 5480
rect 34004 5440 34005 5480
rect 33963 5431 34005 5440
rect 34347 5480 34389 5489
rect 34347 5440 34348 5480
rect 34388 5440 34389 5480
rect 34347 5431 34389 5440
rect 34732 5480 34772 5489
rect 34348 5346 34388 5431
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34155 5144 34197 5153
rect 34155 5104 34156 5144
rect 34196 5104 34197 5144
rect 34155 5095 34197 5104
rect 33772 4985 33812 5070
rect 33579 4976 33621 4985
rect 33579 4936 33580 4976
rect 33620 4936 33621 4976
rect 33579 4927 33621 4936
rect 33771 4976 33813 4985
rect 33771 4936 33772 4976
rect 33812 4936 33813 4976
rect 33771 4927 33813 4936
rect 34156 4976 34196 5095
rect 34732 4987 34772 5440
rect 34828 5153 34868 6196
rect 34924 6187 34964 6196
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35596 5909 35636 7708
rect 35692 6488 35732 8212
rect 36747 8203 36789 8212
rect 36748 7925 36788 8010
rect 36171 7916 36213 7925
rect 36747 7916 36789 7925
rect 36171 7876 36172 7916
rect 36212 7876 36213 7916
rect 36171 7867 36213 7876
rect 36652 7876 36748 7916
rect 36788 7876 36789 7916
rect 36172 7782 36212 7867
rect 36652 7832 36692 7876
rect 36747 7867 36789 7876
rect 36844 7874 36884 7883
rect 36556 7792 36692 7832
rect 36459 7160 36501 7169
rect 36459 7120 36460 7160
rect 36500 7120 36501 7160
rect 36459 7111 36501 7120
rect 36460 7026 36500 7111
rect 36171 6992 36213 7001
rect 36171 6952 36172 6992
rect 36212 6952 36213 6992
rect 36171 6943 36213 6952
rect 35980 6572 36020 6581
rect 35692 6439 35732 6448
rect 35788 6532 35980 6572
rect 35595 5900 35637 5909
rect 35595 5860 35596 5900
rect 35636 5860 35637 5900
rect 35595 5851 35637 5860
rect 34924 5732 34964 5743
rect 35116 5732 35156 5741
rect 34924 5657 34964 5692
rect 35020 5692 35116 5732
rect 34923 5648 34965 5657
rect 34923 5608 34924 5648
rect 34964 5608 34965 5648
rect 34923 5599 34965 5608
rect 34923 5312 34965 5321
rect 34923 5272 34924 5312
rect 34964 5272 34965 5312
rect 34923 5263 34965 5272
rect 34827 5144 34869 5153
rect 34827 5104 34828 5144
rect 34868 5104 34869 5144
rect 34827 5095 34869 5104
rect 34156 4927 34196 4936
rect 34540 4901 34580 4986
rect 34732 4947 34868 4987
rect 34251 4892 34293 4901
rect 34251 4852 34252 4892
rect 34292 4852 34293 4892
rect 34251 4843 34293 4852
rect 34539 4892 34581 4901
rect 34539 4852 34540 4892
rect 34580 4852 34581 4892
rect 34539 4843 34581 4852
rect 34731 4892 34773 4901
rect 34731 4852 34732 4892
rect 34772 4852 34773 4892
rect 34731 4843 34773 4852
rect 33579 4724 33621 4733
rect 33579 4684 33580 4724
rect 33620 4684 33621 4724
rect 33579 4675 33621 4684
rect 33771 4724 33813 4733
rect 33771 4684 33772 4724
rect 33812 4684 33813 4724
rect 33771 4675 33813 4684
rect 33964 4724 34004 4733
rect 33580 4590 33620 4675
rect 33579 3968 33621 3977
rect 33579 3928 33580 3968
rect 33620 3928 33621 3968
rect 33579 3919 33621 3928
rect 33580 3834 33620 3919
rect 33772 3632 33812 4675
rect 33867 4556 33909 4565
rect 33867 4516 33868 4556
rect 33908 4516 33909 4556
rect 33867 4507 33909 4516
rect 33868 4229 33908 4507
rect 33867 4220 33909 4229
rect 33867 4180 33868 4220
rect 33908 4180 33909 4220
rect 33867 4171 33909 4180
rect 33868 4086 33908 4171
rect 33964 3968 34004 4684
rect 34059 4640 34101 4649
rect 34059 4600 34060 4640
rect 34100 4600 34101 4640
rect 34059 4591 34101 4600
rect 34060 4388 34100 4591
rect 34252 4397 34292 4843
rect 34732 4758 34772 4843
rect 34348 4724 34388 4733
rect 34636 4724 34676 4733
rect 34388 4684 34580 4724
rect 34348 4675 34388 4684
rect 34347 4556 34389 4565
rect 34347 4516 34348 4556
rect 34388 4516 34389 4556
rect 34347 4507 34389 4516
rect 34060 4339 34100 4348
rect 34251 4388 34293 4397
rect 34251 4348 34252 4388
rect 34292 4348 34293 4388
rect 34251 4339 34293 4348
rect 34060 4220 34100 4231
rect 34060 4145 34100 4180
rect 34252 4145 34292 4339
rect 34059 4136 34101 4145
rect 34059 4096 34060 4136
rect 34100 4096 34101 4136
rect 34059 4087 34101 4096
rect 34251 4136 34293 4145
rect 34251 4096 34252 4136
rect 34292 4096 34293 4136
rect 34251 4087 34293 4096
rect 34348 4052 34388 4507
rect 34444 4229 34484 4314
rect 34443 4220 34485 4229
rect 34443 4180 34444 4220
rect 34484 4180 34485 4220
rect 34443 4171 34485 4180
rect 34444 4052 34484 4061
rect 34348 4012 34444 4052
rect 34444 4003 34484 4012
rect 33964 3928 34388 3968
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34251 3632 34293 3641
rect 33772 3592 34004 3632
rect 33484 3415 33524 3424
rect 33579 3464 33621 3473
rect 33868 3464 33908 3473
rect 33579 3424 33580 3464
rect 33620 3424 33868 3464
rect 33579 3415 33621 3424
rect 33868 3415 33908 3424
rect 33676 3212 33716 3221
rect 33676 2540 33716 3172
rect 33867 2876 33909 2885
rect 33867 2836 33868 2876
rect 33908 2836 33909 2876
rect 33867 2827 33909 2836
rect 33676 2500 33812 2540
rect 33388 2332 33716 2372
rect 33292 1324 33428 1364
rect 33291 1196 33333 1205
rect 33291 1156 33292 1196
rect 33332 1156 33333 1196
rect 33291 1147 33333 1156
rect 33292 80 33332 1147
rect 33388 953 33428 1324
rect 33483 1280 33525 1289
rect 33483 1240 33484 1280
rect 33524 1240 33525 1280
rect 33483 1231 33525 1240
rect 33387 944 33429 953
rect 33387 904 33388 944
rect 33428 904 33429 944
rect 33387 895 33429 904
rect 33484 80 33524 1231
rect 33676 80 33716 2332
rect 33772 1037 33812 2500
rect 33771 1028 33813 1037
rect 33771 988 33772 1028
rect 33812 988 33813 1028
rect 33771 979 33813 988
rect 33868 80 33908 2827
rect 33964 2381 34004 3592
rect 34251 3592 34252 3632
rect 34292 3592 34293 3632
rect 34251 3583 34293 3592
rect 34252 3464 34292 3583
rect 34252 3415 34292 3424
rect 34060 3212 34100 3221
rect 34100 3172 34196 3212
rect 34060 3163 34100 3172
rect 34059 2792 34101 2801
rect 34059 2752 34060 2792
rect 34100 2752 34101 2792
rect 34059 2743 34101 2752
rect 33963 2372 34005 2381
rect 33963 2332 33964 2372
rect 34004 2332 34005 2372
rect 33963 2323 34005 2332
rect 34060 80 34100 2743
rect 34156 1121 34196 3172
rect 34348 2297 34388 3928
rect 34444 3212 34484 3221
rect 34540 3212 34580 4684
rect 34636 4481 34676 4684
rect 34635 4472 34677 4481
rect 34635 4432 34636 4472
rect 34676 4432 34677 4472
rect 34635 4423 34677 4432
rect 34636 4220 34676 4229
rect 34636 4061 34676 4180
rect 34731 4220 34773 4229
rect 34731 4180 34732 4220
rect 34772 4180 34773 4220
rect 34731 4171 34773 4180
rect 34635 4052 34677 4061
rect 34635 4012 34636 4052
rect 34676 4012 34677 4052
rect 34635 4003 34677 4012
rect 34732 3380 34772 4171
rect 34828 3968 34868 4947
rect 34924 4892 34964 5263
rect 35020 4892 35060 5692
rect 35116 5683 35156 5692
rect 35403 5732 35445 5741
rect 35403 5692 35404 5732
rect 35444 5692 35445 5732
rect 35403 5683 35445 5692
rect 35596 5732 35636 5741
rect 35788 5732 35828 6532
rect 35980 6523 36020 6532
rect 35877 6404 35924 6413
rect 35877 6364 35878 6404
rect 35877 6355 35924 6364
rect 35979 6404 36021 6413
rect 35979 6364 35980 6404
rect 36020 6364 36021 6404
rect 35979 6355 36021 6364
rect 36172 6404 36212 6943
rect 36556 6656 36596 7792
rect 36748 7748 36788 7757
rect 36748 7589 36788 7708
rect 36844 7673 36884 7834
rect 36843 7664 36885 7673
rect 36843 7624 36844 7664
rect 36884 7624 36885 7664
rect 36843 7615 36885 7624
rect 36747 7580 36789 7589
rect 36747 7540 36748 7580
rect 36788 7540 36789 7580
rect 36747 7531 36789 7540
rect 36652 7412 36692 7421
rect 36748 7412 36788 7531
rect 36692 7372 36788 7412
rect 36652 7363 36692 7372
rect 36651 6992 36693 7001
rect 36651 6952 36652 6992
rect 36692 6952 36693 6992
rect 36651 6943 36693 6952
rect 36652 6858 36692 6943
rect 36843 6824 36885 6833
rect 36843 6784 36844 6824
rect 36884 6784 36885 6824
rect 36843 6775 36885 6784
rect 36652 6656 36692 6665
rect 36556 6616 36652 6656
rect 36652 6607 36692 6616
rect 36844 6413 36884 6775
rect 36172 6355 36212 6364
rect 36363 6404 36405 6413
rect 36363 6364 36364 6404
rect 36404 6364 36405 6404
rect 36363 6355 36405 6364
rect 36843 6404 36885 6413
rect 36843 6364 36844 6404
rect 36884 6364 36885 6404
rect 36843 6355 36885 6364
rect 35878 6275 35918 6355
rect 35980 6270 36020 6355
rect 36364 6270 36404 6355
rect 36268 5741 36308 5826
rect 36076 5732 36116 5741
rect 36267 5732 36309 5741
rect 35636 5692 36020 5732
rect 35596 5683 35636 5692
rect 35404 5598 35444 5683
rect 35116 5480 35156 5489
rect 35116 5153 35156 5440
rect 35307 5396 35349 5405
rect 35307 5356 35308 5396
rect 35348 5356 35349 5396
rect 35307 5347 35349 5356
rect 35115 5144 35157 5153
rect 35115 5104 35116 5144
rect 35156 5104 35157 5144
rect 35115 5095 35157 5104
rect 35308 4976 35348 5347
rect 35403 5228 35445 5237
rect 35403 5188 35404 5228
rect 35444 5188 35445 5228
rect 35403 5179 35445 5188
rect 35404 5060 35444 5179
rect 35404 5020 35636 5060
rect 35308 4936 35444 4976
rect 35115 4892 35157 4901
rect 35020 4852 35116 4892
rect 35156 4852 35157 4892
rect 34924 4843 34964 4852
rect 35115 4843 35157 4852
rect 35308 4881 35348 4890
rect 35116 4758 35156 4843
rect 35308 4817 35348 4841
rect 35307 4808 35349 4817
rect 35307 4768 35308 4808
rect 35348 4768 35349 4808
rect 35307 4759 35349 4768
rect 35404 4808 35444 4936
rect 35596 4892 35636 5020
rect 35884 4901 35924 4986
rect 35692 4892 35732 4901
rect 35404 4759 35444 4768
rect 35500 4881 35540 4890
rect 35308 4746 35348 4759
rect 35500 4733 35540 4841
rect 35596 4852 35692 4892
rect 35019 4724 35061 4733
rect 35019 4684 35020 4724
rect 35060 4684 35061 4724
rect 35019 4675 35061 4684
rect 35499 4724 35541 4733
rect 35499 4684 35500 4724
rect 35540 4684 35541 4724
rect 35499 4675 35541 4684
rect 35020 4590 35060 4675
rect 35596 4565 35636 4852
rect 35692 4843 35732 4852
rect 35883 4892 35925 4901
rect 35883 4852 35884 4892
rect 35924 4852 35925 4892
rect 35980 4892 36020 5692
rect 36116 5692 36212 5732
rect 36076 5683 36116 5692
rect 36076 4892 36116 4901
rect 35980 4852 36076 4892
rect 35883 4843 35925 4852
rect 36076 4843 36116 4852
rect 36172 4733 36212 5692
rect 36267 5692 36268 5732
rect 36308 5692 36309 5732
rect 36267 5683 36309 5692
rect 36460 5732 36500 5743
rect 36460 5657 36500 5692
rect 36555 5732 36597 5741
rect 36652 5732 36692 5741
rect 36555 5692 36556 5732
rect 36596 5692 36652 5732
rect 36555 5683 36597 5692
rect 36652 5683 36692 5692
rect 36844 5732 36884 6355
rect 36844 5683 36884 5692
rect 36459 5648 36501 5657
rect 36459 5608 36460 5648
rect 36500 5608 36501 5648
rect 36459 5599 36501 5608
rect 36268 5480 36308 5489
rect 36308 5440 36404 5480
rect 36268 5431 36308 5440
rect 36267 4892 36309 4901
rect 36267 4852 36268 4892
rect 36308 4852 36309 4892
rect 36267 4843 36309 4852
rect 36268 4758 36308 4843
rect 35691 4724 35733 4733
rect 35691 4684 35692 4724
rect 35732 4684 35733 4724
rect 35691 4675 35733 4684
rect 35788 4724 35828 4733
rect 36171 4724 36213 4733
rect 35828 4684 35924 4724
rect 35788 4675 35828 4684
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35595 4556 35637 4565
rect 35595 4516 35596 4556
rect 35636 4516 35637 4556
rect 35595 4507 35637 4516
rect 35020 4430 35060 4483
rect 35596 4430 35636 4507
rect 35019 4390 35020 4397
rect 35060 4390 35061 4397
rect 35019 4388 35061 4390
rect 35404 4390 35636 4430
rect 35404 4388 35444 4390
rect 35019 4348 35020 4388
rect 35060 4348 35061 4388
rect 35019 4339 35061 4348
rect 35212 4348 35444 4388
rect 35019 4220 35061 4229
rect 35019 4180 35020 4220
rect 35060 4180 35061 4220
rect 35019 4171 35061 4180
rect 35212 4220 35252 4348
rect 35212 4171 35252 4180
rect 35499 4220 35541 4229
rect 35588 4220 35628 4228
rect 35499 4180 35500 4220
rect 35540 4219 35628 4220
rect 35540 4180 35588 4219
rect 35499 4171 35541 4180
rect 35692 4220 35732 4675
rect 35788 4397 35828 4482
rect 35787 4388 35829 4397
rect 35787 4348 35788 4388
rect 35828 4348 35829 4388
rect 35787 4339 35829 4348
rect 35788 4220 35828 4229
rect 35692 4180 35788 4220
rect 35020 4086 35060 4171
rect 35588 4170 35628 4179
rect 35115 4136 35157 4145
rect 35115 4096 35116 4136
rect 35156 4096 35157 4136
rect 35115 4087 35157 4096
rect 34828 3928 34964 3968
rect 34924 3557 34964 3928
rect 35019 3716 35061 3725
rect 35019 3676 35020 3716
rect 35060 3676 35061 3716
rect 35019 3667 35061 3676
rect 34923 3548 34965 3557
rect 34923 3508 34924 3548
rect 34964 3508 34965 3548
rect 34923 3499 34965 3508
rect 34732 3331 34772 3340
rect 34924 3380 34964 3389
rect 35020 3380 35060 3667
rect 35116 3641 35156 4087
rect 35595 3884 35637 3893
rect 35595 3844 35596 3884
rect 35636 3844 35637 3884
rect 35595 3835 35637 3844
rect 35307 3800 35349 3809
rect 35307 3760 35308 3800
rect 35348 3760 35349 3800
rect 35307 3751 35349 3760
rect 35115 3632 35157 3641
rect 35115 3592 35116 3632
rect 35156 3592 35157 3632
rect 35115 3583 35157 3592
rect 35308 3464 35348 3751
rect 35308 3415 35348 3424
rect 34964 3340 35060 3380
rect 34924 3331 34964 3340
rect 35500 3221 35540 3306
rect 34924 3212 34964 3221
rect 34540 3172 34772 3212
rect 34444 2540 34484 3172
rect 34635 2960 34677 2969
rect 34635 2920 34636 2960
rect 34676 2920 34677 2960
rect 34635 2911 34677 2920
rect 34444 2500 34580 2540
rect 34443 2372 34485 2381
rect 34443 2332 34444 2372
rect 34484 2332 34485 2372
rect 34443 2323 34485 2332
rect 34347 2288 34389 2297
rect 34347 2248 34348 2288
rect 34388 2248 34389 2288
rect 34347 2239 34389 2248
rect 34251 1784 34293 1793
rect 34251 1744 34252 1784
rect 34292 1744 34293 1784
rect 34251 1735 34293 1744
rect 34155 1112 34197 1121
rect 34155 1072 34156 1112
rect 34196 1072 34197 1112
rect 34155 1063 34197 1072
rect 34252 80 34292 1735
rect 34444 80 34484 2323
rect 34540 1625 34580 2500
rect 34539 1616 34581 1625
rect 34539 1576 34540 1616
rect 34580 1576 34581 1616
rect 34539 1567 34581 1576
rect 34636 80 34676 2911
rect 34732 1289 34772 3172
rect 34827 2036 34869 2045
rect 34827 1996 34828 2036
rect 34868 1996 34869 2036
rect 34827 1987 34869 1996
rect 34731 1280 34773 1289
rect 34731 1240 34732 1280
rect 34772 1240 34773 1280
rect 34731 1231 34773 1240
rect 34828 80 34868 1987
rect 34924 1373 34964 3172
rect 35499 3212 35541 3221
rect 35499 3172 35500 3212
rect 35540 3172 35541 3212
rect 35499 3163 35541 3172
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35211 2708 35253 2717
rect 35211 2668 35212 2708
rect 35252 2668 35253 2708
rect 35211 2659 35253 2668
rect 35019 2288 35061 2297
rect 35019 2248 35020 2288
rect 35060 2248 35061 2288
rect 35019 2239 35061 2248
rect 34923 1364 34965 1373
rect 34923 1324 34924 1364
rect 34964 1324 34965 1364
rect 34923 1315 34965 1324
rect 35020 80 35060 2239
rect 35212 80 35252 2659
rect 35403 1196 35445 1205
rect 35403 1156 35404 1196
rect 35444 1156 35445 1196
rect 35403 1147 35445 1156
rect 35404 80 35444 1147
rect 35596 80 35636 3835
rect 35691 3464 35733 3473
rect 35691 3424 35692 3464
rect 35732 3424 35733 3464
rect 35691 3415 35733 3424
rect 35692 3330 35732 3415
rect 35788 3305 35828 4180
rect 35884 3809 35924 4684
rect 36171 4684 36172 4724
rect 36212 4684 36213 4724
rect 36171 4675 36213 4684
rect 36075 4304 36117 4313
rect 36075 4264 36076 4304
rect 36116 4264 36117 4304
rect 36075 4255 36117 4264
rect 36076 4136 36116 4255
rect 36076 4087 36116 4096
rect 36172 4061 36212 4675
rect 36171 4052 36213 4061
rect 36171 4012 36172 4052
rect 36212 4012 36213 4052
rect 36364 4052 36404 5440
rect 36459 4976 36501 4985
rect 36459 4936 36460 4976
rect 36500 4936 36501 4976
rect 36459 4927 36501 4936
rect 36460 4149 36500 4927
rect 36556 4901 36596 5683
rect 36940 5648 36980 8800
rect 37035 8756 37077 8765
rect 37035 8716 37036 8756
rect 37076 8716 37077 8756
rect 37035 8707 37077 8716
rect 37132 8756 37172 9388
rect 37228 8924 37268 10648
rect 37323 10520 37365 10529
rect 37323 10480 37324 10520
rect 37364 10480 37365 10520
rect 37323 10471 37365 10480
rect 37324 10277 37364 10471
rect 37323 10268 37365 10277
rect 37323 10228 37324 10268
rect 37364 10228 37365 10268
rect 37323 10219 37365 10228
rect 37420 10268 37460 10807
rect 37996 10361 38036 10807
rect 38091 10604 38133 10613
rect 38091 10564 38092 10604
rect 38132 10564 38133 10604
rect 38091 10555 38133 10564
rect 37995 10352 38037 10361
rect 37995 10312 37996 10352
rect 38036 10312 38037 10352
rect 37995 10303 38037 10312
rect 37420 10219 37460 10228
rect 37611 10268 37653 10277
rect 37611 10228 37612 10268
rect 37652 10228 37653 10268
rect 37611 10219 37653 10228
rect 37803 10268 37845 10277
rect 37803 10228 37804 10268
rect 37844 10228 37845 10268
rect 37803 10219 37845 10228
rect 37996 10268 38036 10303
rect 37612 10134 37652 10219
rect 37804 10134 37844 10219
rect 37996 10218 38036 10228
rect 38092 10109 38132 10555
rect 38763 10520 38805 10529
rect 38763 10480 38764 10520
rect 38804 10480 38805 10520
rect 38763 10471 38805 10480
rect 38379 10436 38421 10445
rect 38379 10396 38380 10436
rect 38420 10396 38421 10436
rect 38379 10387 38421 10396
rect 38187 10268 38229 10277
rect 38187 10228 38188 10268
rect 38228 10228 38229 10268
rect 38187 10219 38229 10228
rect 38380 10268 38420 10387
rect 38764 10361 38804 10471
rect 38763 10352 38805 10361
rect 38763 10312 38764 10352
rect 38804 10312 38805 10352
rect 38763 10303 38805 10312
rect 38380 10219 38420 10228
rect 38571 10268 38613 10277
rect 38571 10228 38572 10268
rect 38612 10228 38613 10268
rect 38571 10219 38613 10228
rect 38764 10268 38804 10303
rect 37899 10100 37941 10109
rect 37899 10060 37900 10100
rect 37940 10060 37941 10100
rect 37899 10051 37941 10060
rect 38091 10100 38133 10109
rect 38091 10060 38092 10100
rect 38132 10060 38133 10100
rect 38091 10051 38133 10060
rect 37516 10016 37556 10025
rect 37516 9521 37556 9976
rect 37900 9966 37940 10051
rect 38188 9848 38228 10219
rect 38572 10134 38612 10219
rect 38764 10218 38804 10228
rect 38955 10268 38997 10277
rect 38955 10228 38956 10268
rect 38996 10228 38997 10268
rect 38955 10219 38997 10228
rect 39148 10268 39188 10279
rect 38956 10134 38996 10219
rect 39148 10193 39188 10228
rect 39147 10184 39189 10193
rect 39147 10144 39148 10184
rect 39188 10144 39189 10184
rect 39147 10135 39189 10144
rect 38379 10100 38421 10109
rect 38379 10060 38380 10100
rect 38420 10060 38421 10100
rect 38379 10051 38421 10060
rect 37996 9808 38228 9848
rect 38284 10016 38324 10025
rect 37899 9680 37941 9689
rect 37899 9640 37900 9680
rect 37940 9640 37941 9680
rect 37899 9631 37941 9640
rect 37515 9512 37557 9521
rect 37515 9472 37516 9512
rect 37556 9472 37557 9512
rect 37515 9463 37557 9472
rect 37900 9437 37940 9631
rect 37323 9428 37365 9437
rect 37323 9388 37324 9428
rect 37364 9388 37365 9428
rect 37323 9379 37365 9388
rect 37899 9428 37941 9437
rect 37899 9388 37900 9428
rect 37940 9388 37941 9428
rect 37899 9379 37941 9388
rect 37996 9428 38036 9808
rect 37324 9294 37364 9379
rect 37996 9269 38036 9388
rect 38187 9428 38229 9437
rect 38187 9388 38188 9428
rect 38228 9388 38229 9428
rect 38187 9379 38229 9388
rect 38092 9344 38132 9353
rect 37803 9260 37845 9269
rect 37803 9220 37804 9260
rect 37844 9220 37845 9260
rect 37803 9211 37845 9220
rect 37995 9260 38037 9269
rect 37995 9220 37996 9260
rect 38036 9220 38037 9260
rect 37995 9211 38037 9220
rect 37228 8884 37364 8924
rect 37228 8756 37268 8784
rect 37324 8765 37364 8884
rect 37132 8716 37228 8756
rect 37036 8622 37076 8707
rect 37036 8168 37076 8177
rect 37132 8168 37172 8716
rect 37228 8707 37268 8716
rect 37323 8756 37365 8765
rect 37323 8716 37324 8756
rect 37364 8716 37365 8756
rect 37323 8707 37365 8716
rect 37323 8504 37365 8513
rect 37323 8464 37324 8504
rect 37364 8464 37365 8504
rect 37323 8455 37365 8464
rect 37076 8128 37172 8168
rect 37036 8119 37076 8128
rect 37227 7496 37269 7505
rect 37227 7456 37228 7496
rect 37268 7456 37269 7496
rect 37227 7447 37269 7456
rect 37228 6161 37268 7447
rect 37324 7412 37364 8455
rect 37707 8084 37749 8093
rect 37707 8044 37708 8084
rect 37748 8044 37749 8084
rect 37707 8035 37749 8044
rect 37420 7925 37460 8010
rect 37708 7950 37748 8035
rect 37419 7916 37461 7925
rect 37419 7876 37420 7916
rect 37460 7876 37461 7916
rect 37419 7867 37461 7876
rect 37516 7916 37556 7925
rect 37420 7748 37460 7757
rect 37420 7589 37460 7708
rect 37419 7580 37461 7589
rect 37419 7540 37420 7580
rect 37460 7540 37461 7580
rect 37419 7531 37461 7540
rect 37516 7505 37556 7876
rect 37611 7580 37653 7589
rect 37611 7540 37612 7580
rect 37652 7540 37653 7580
rect 37611 7531 37653 7540
rect 37515 7496 37557 7505
rect 37515 7456 37516 7496
rect 37556 7456 37557 7496
rect 37515 7447 37557 7456
rect 37324 7372 37460 7412
rect 37323 7244 37365 7253
rect 37323 7204 37324 7244
rect 37364 7204 37365 7244
rect 37323 7195 37365 7204
rect 37324 7110 37364 7195
rect 37324 6497 37364 6528
rect 37323 6488 37365 6497
rect 37323 6448 37324 6488
rect 37364 6448 37365 6488
rect 37323 6439 37365 6448
rect 37324 6404 37364 6439
rect 37324 6245 37364 6364
rect 37323 6236 37365 6245
rect 37323 6196 37324 6236
rect 37364 6196 37365 6236
rect 37323 6187 37365 6196
rect 37227 6152 37269 6161
rect 37227 6112 37228 6152
rect 37268 6112 37269 6152
rect 37227 6103 37269 6112
rect 37228 5984 37268 6103
rect 37228 5944 37273 5984
rect 37036 5825 37076 5838
rect 37035 5816 37077 5825
rect 37035 5776 37036 5816
rect 37076 5776 37077 5816
rect 37035 5767 37077 5776
rect 37036 5743 37076 5767
rect 37233 5741 37273 5944
rect 37036 5694 37076 5703
rect 37228 5732 37273 5741
rect 37268 5692 37273 5732
rect 37228 5683 37268 5692
rect 36940 5608 37172 5648
rect 36652 5480 36692 5489
rect 37036 5480 37076 5489
rect 36692 5440 36884 5480
rect 36652 5431 36692 5440
rect 36651 4976 36693 4985
rect 36651 4936 36652 4976
rect 36692 4936 36693 4976
rect 36651 4927 36693 4936
rect 36555 4892 36597 4901
rect 36555 4852 36556 4892
rect 36596 4852 36597 4892
rect 36555 4843 36597 4852
rect 36556 4758 36596 4843
rect 36652 4842 36692 4927
rect 36748 4892 36788 4901
rect 36748 4565 36788 4852
rect 36747 4556 36789 4565
rect 36747 4516 36748 4556
rect 36788 4516 36789 4556
rect 36747 4507 36789 4516
rect 36460 4100 36500 4109
rect 36844 4136 36884 5440
rect 36844 4087 36884 4096
rect 36940 5440 37036 5480
rect 36364 4012 36500 4052
rect 36171 4003 36213 4012
rect 36268 3968 36308 3977
rect 36308 3928 36404 3968
rect 36268 3919 36308 3928
rect 35883 3800 35925 3809
rect 35883 3760 35884 3800
rect 35924 3760 35925 3800
rect 35883 3751 35925 3760
rect 36075 3464 36117 3473
rect 36075 3424 36076 3464
rect 36116 3424 36117 3464
rect 36075 3415 36117 3424
rect 36076 3330 36116 3415
rect 35787 3296 35829 3305
rect 35787 3256 35788 3296
rect 35828 3256 35829 3296
rect 35787 3247 35829 3256
rect 35788 2969 35828 3247
rect 35884 3212 35924 3221
rect 35787 2960 35829 2969
rect 35787 2920 35788 2960
rect 35828 2920 35829 2960
rect 35787 2911 35829 2920
rect 35884 1709 35924 3172
rect 36268 3212 36308 3221
rect 35883 1700 35925 1709
rect 35883 1660 35884 1700
rect 35924 1660 35925 1700
rect 35883 1651 35925 1660
rect 35787 1280 35829 1289
rect 35787 1240 35788 1280
rect 35828 1240 35829 1280
rect 35787 1231 35829 1240
rect 35788 80 35828 1231
rect 36171 944 36213 953
rect 36171 904 36172 944
rect 36212 904 36213 944
rect 36171 895 36213 904
rect 35979 860 36021 869
rect 35979 820 35980 860
rect 36020 820 36021 860
rect 35979 811 36021 820
rect 35980 80 36020 811
rect 36172 80 36212 895
rect 36268 197 36308 3172
rect 36364 1289 36404 3928
rect 36460 3464 36500 4012
rect 36652 3968 36692 3977
rect 36692 3928 36788 3968
rect 36652 3919 36692 3928
rect 36460 3415 36500 3424
rect 36652 3212 36692 3221
rect 36652 1457 36692 3172
rect 36748 2045 36788 3928
rect 36843 3800 36885 3809
rect 36843 3760 36844 3800
rect 36884 3760 36885 3800
rect 36843 3751 36885 3760
rect 36844 3464 36884 3751
rect 36844 3415 36884 3424
rect 36940 3305 36980 5440
rect 37036 5431 37076 5440
rect 37132 4976 37172 5608
rect 37323 5480 37365 5489
rect 37323 5440 37324 5480
rect 37364 5440 37365 5480
rect 37323 5431 37365 5440
rect 37324 5346 37364 5431
rect 37132 4927 37172 4936
rect 37035 4892 37077 4901
rect 37035 4852 37036 4892
rect 37076 4852 37077 4892
rect 37035 4843 37077 4852
rect 37227 4892 37269 4901
rect 37227 4852 37228 4892
rect 37268 4852 37269 4892
rect 37227 4843 37269 4852
rect 37036 4136 37076 4843
rect 37228 4149 37268 4843
rect 37036 4096 37172 4136
rect 37228 4100 37268 4109
rect 37324 4724 37364 4733
rect 37132 4052 37172 4096
rect 37132 4012 37268 4052
rect 37036 3968 37076 3977
rect 37076 3928 37172 3968
rect 37036 3919 37076 3928
rect 36939 3296 36981 3305
rect 36939 3256 36940 3296
rect 36980 3256 36981 3296
rect 36939 3247 36981 3256
rect 37036 3212 37076 3221
rect 36939 3128 36981 3137
rect 36939 3088 36940 3128
rect 36980 3088 36981 3128
rect 36939 3079 36981 3088
rect 36747 2036 36789 2045
rect 36747 1996 36748 2036
rect 36788 1996 36789 2036
rect 36747 1987 36789 1996
rect 36747 1616 36789 1625
rect 36747 1576 36748 1616
rect 36788 1576 36789 1616
rect 36747 1567 36789 1576
rect 36651 1448 36693 1457
rect 36651 1408 36652 1448
rect 36692 1408 36693 1448
rect 36651 1399 36693 1408
rect 36363 1280 36405 1289
rect 36363 1240 36364 1280
rect 36404 1240 36405 1280
rect 36363 1231 36405 1240
rect 36555 1112 36597 1121
rect 36555 1072 36556 1112
rect 36596 1072 36597 1112
rect 36555 1063 36597 1072
rect 36363 1028 36405 1037
rect 36363 988 36364 1028
rect 36404 988 36405 1028
rect 36363 979 36405 988
rect 36267 188 36309 197
rect 36267 148 36268 188
rect 36308 148 36309 188
rect 36267 139 36309 148
rect 36364 80 36404 979
rect 36556 80 36596 1063
rect 36748 80 36788 1567
rect 36940 80 36980 3079
rect 37036 1205 37076 3172
rect 37132 2129 37172 3928
rect 37228 3464 37268 4012
rect 37228 3415 37268 3424
rect 37227 3296 37269 3305
rect 37227 3256 37228 3296
rect 37268 3256 37269 3296
rect 37227 3247 37269 3256
rect 37228 2465 37268 3247
rect 37227 2456 37269 2465
rect 37227 2416 37228 2456
rect 37268 2416 37269 2456
rect 37227 2407 37269 2416
rect 37131 2120 37173 2129
rect 37131 2080 37132 2120
rect 37172 2080 37173 2120
rect 37131 2071 37173 2080
rect 37131 1280 37173 1289
rect 37131 1240 37132 1280
rect 37172 1240 37173 1280
rect 37131 1231 37173 1240
rect 37035 1196 37077 1205
rect 37035 1156 37036 1196
rect 37076 1156 37077 1196
rect 37035 1147 37077 1156
rect 37132 80 37172 1231
rect 37324 80 37364 4684
rect 37420 4136 37460 7372
rect 37516 7253 37556 7338
rect 37515 7244 37557 7253
rect 37515 7204 37516 7244
rect 37556 7204 37557 7244
rect 37515 7195 37557 7204
rect 37515 6992 37557 7001
rect 37515 6952 37516 6992
rect 37556 6952 37557 6992
rect 37515 6943 37557 6952
rect 37516 6858 37556 6943
rect 37612 6404 37652 7531
rect 37707 7328 37749 7337
rect 37707 7288 37708 7328
rect 37748 7288 37749 7328
rect 37707 7279 37749 7288
rect 37708 7244 37748 7279
rect 37708 7169 37748 7204
rect 37707 7160 37749 7169
rect 37707 7120 37708 7160
rect 37748 7120 37749 7160
rect 37707 7111 37749 7120
rect 37708 7080 37748 7111
rect 37804 6656 37844 9211
rect 38092 9185 38132 9304
rect 38188 9294 38228 9379
rect 38091 9176 38133 9185
rect 38091 9136 38092 9176
rect 38132 9136 38133 9176
rect 38091 9127 38133 9136
rect 37995 8924 38037 8933
rect 38284 8924 38324 9976
rect 38380 9932 38420 10051
rect 38668 10016 38708 10025
rect 38380 9892 38612 9932
rect 38380 9428 38420 9437
rect 38380 9269 38420 9388
rect 38572 9428 38612 9892
rect 38572 9379 38612 9388
rect 38475 9344 38517 9353
rect 38475 9304 38476 9344
rect 38516 9304 38517 9344
rect 38475 9295 38517 9304
rect 38379 9260 38421 9269
rect 38379 9220 38380 9260
rect 38420 9220 38421 9260
rect 38379 9211 38421 9220
rect 38380 9017 38420 9211
rect 38476 9210 38516 9295
rect 38571 9092 38613 9101
rect 38571 9052 38572 9092
rect 38612 9052 38613 9092
rect 38571 9043 38613 9052
rect 38379 9008 38421 9017
rect 38379 8968 38380 9008
rect 38420 8968 38421 9008
rect 38379 8959 38421 8968
rect 37995 8884 37996 8924
rect 38036 8884 38037 8924
rect 37995 8875 38037 8884
rect 38188 8884 38324 8924
rect 37900 7253 37940 7338
rect 37899 7244 37941 7253
rect 37899 7204 37900 7244
rect 37940 7204 37941 7244
rect 37899 7195 37941 7204
rect 37612 6355 37652 6364
rect 37708 6616 37844 6656
rect 37900 6992 37940 7001
rect 37708 6320 37748 6616
rect 37900 6581 37940 6952
rect 37899 6572 37941 6581
rect 37804 6497 37844 6541
rect 37899 6532 37900 6572
rect 37940 6532 37941 6572
rect 37899 6523 37941 6532
rect 37803 6488 37845 6497
rect 37803 6448 37804 6488
rect 37844 6448 37845 6488
rect 37803 6446 37845 6448
rect 37803 6439 37804 6446
rect 37844 6439 37845 6446
rect 37804 6397 37844 6406
rect 37900 6404 37940 6415
rect 37900 6329 37940 6364
rect 37899 6320 37941 6329
rect 37708 6280 37844 6320
rect 37612 6236 37652 6245
rect 37652 6196 37748 6236
rect 37612 6187 37652 6196
rect 37516 5825 37556 5856
rect 37515 5816 37557 5825
rect 37515 5776 37516 5816
rect 37556 5776 37557 5816
rect 37515 5767 37557 5776
rect 37516 5732 37556 5767
rect 37708 5741 37748 6196
rect 37516 5573 37556 5692
rect 37707 5732 37749 5741
rect 37707 5692 37708 5732
rect 37748 5692 37749 5732
rect 37707 5683 37749 5692
rect 37515 5564 37557 5573
rect 37515 5524 37516 5564
rect 37556 5524 37557 5564
rect 37515 5515 37557 5524
rect 37707 5480 37749 5489
rect 37707 5440 37708 5480
rect 37748 5440 37749 5480
rect 37707 5431 37749 5440
rect 37708 5346 37748 5431
rect 37515 4976 37557 4985
rect 37515 4936 37516 4976
rect 37556 4936 37557 4976
rect 37515 4927 37557 4936
rect 37516 4842 37556 4927
rect 37611 4808 37653 4817
rect 37611 4768 37612 4808
rect 37652 4768 37653 4808
rect 37611 4759 37653 4768
rect 37612 4313 37652 4759
rect 37708 4724 37748 4733
rect 37611 4304 37653 4313
rect 37611 4264 37612 4304
rect 37652 4264 37653 4304
rect 37611 4255 37653 4264
rect 37612 4220 37652 4255
rect 37612 4169 37652 4180
rect 37420 4096 37556 4136
rect 37420 3968 37460 3977
rect 37420 3389 37460 3928
rect 37516 3464 37556 4096
rect 37612 3464 37652 3473
rect 37516 3424 37612 3464
rect 37612 3415 37652 3424
rect 37419 3380 37461 3389
rect 37419 3340 37420 3380
rect 37460 3340 37461 3380
rect 37419 3331 37461 3340
rect 37420 3212 37460 3221
rect 37420 1625 37460 3172
rect 37515 3212 37557 3221
rect 37515 3172 37516 3212
rect 37556 3172 37557 3212
rect 37515 3163 37557 3172
rect 37516 3053 37556 3163
rect 37515 3044 37557 3053
rect 37515 3004 37516 3044
rect 37556 3004 37557 3044
rect 37515 2995 37557 3004
rect 37708 2540 37748 4684
rect 37804 4397 37844 6280
rect 37899 6280 37900 6320
rect 37940 6280 37941 6320
rect 37899 6271 37941 6280
rect 37899 6068 37941 6077
rect 37899 6028 37900 6068
rect 37940 6028 37941 6068
rect 37899 6019 37941 6028
rect 37900 5732 37940 6019
rect 37900 5489 37940 5692
rect 37899 5480 37941 5489
rect 37899 5440 37900 5480
rect 37940 5440 37941 5480
rect 37899 5431 37941 5440
rect 37900 4976 37940 4985
rect 37996 4976 38036 8875
rect 38188 8261 38228 8884
rect 38284 8756 38324 8765
rect 38380 8756 38420 8959
rect 38476 8756 38516 8765
rect 38380 8716 38476 8756
rect 38187 8252 38229 8261
rect 38187 8212 38188 8252
rect 38228 8212 38229 8252
rect 38187 8203 38229 8212
rect 38284 8093 38324 8716
rect 38476 8707 38516 8716
rect 38283 8084 38325 8093
rect 38283 8044 38284 8084
rect 38324 8044 38325 8084
rect 38283 8035 38325 8044
rect 38283 7244 38325 7253
rect 38283 7204 38284 7244
rect 38324 7204 38325 7244
rect 38283 7195 38325 7204
rect 38091 6740 38133 6749
rect 38091 6700 38092 6740
rect 38132 6700 38133 6740
rect 38091 6691 38133 6700
rect 38092 6413 38132 6691
rect 38091 6404 38133 6413
rect 38091 6364 38092 6404
rect 38132 6364 38133 6404
rect 38091 6355 38133 6364
rect 38284 6404 38324 7195
rect 38284 6329 38324 6364
rect 38283 6320 38325 6329
rect 38572 6320 38612 9043
rect 38668 8345 38708 9976
rect 39052 10016 39092 10025
rect 38764 9428 38804 9437
rect 38764 9017 38804 9388
rect 38955 9428 38997 9437
rect 38955 9388 38956 9428
rect 38996 9388 38997 9428
rect 38955 9379 38997 9388
rect 38860 9344 38900 9353
rect 38860 9101 38900 9304
rect 38956 9294 38996 9379
rect 38859 9092 38901 9101
rect 38859 9052 38860 9092
rect 38900 9052 38901 9092
rect 38859 9043 38901 9052
rect 38763 9008 38805 9017
rect 38763 8968 38764 9008
rect 38804 8968 38805 9008
rect 38763 8959 38805 8968
rect 38667 8336 38709 8345
rect 38667 8296 38668 8336
rect 38708 8296 38709 8336
rect 38667 8287 38709 8296
rect 39052 8177 39092 9976
rect 39051 8168 39093 8177
rect 39051 8128 39052 8168
rect 39092 8128 39093 8168
rect 39051 8119 39093 8128
rect 39244 7505 39284 10900
rect 39340 10891 39380 10900
rect 40779 10940 40821 10949
rect 40779 10900 40780 10940
rect 40820 10900 40821 10940
rect 40779 10891 40821 10900
rect 40587 10772 40629 10781
rect 40587 10732 40588 10772
rect 40628 10732 40629 10772
rect 40587 10723 40629 10732
rect 40588 10268 40628 10723
rect 40588 10219 40628 10228
rect 40683 10184 40725 10193
rect 40683 10144 40684 10184
rect 40724 10144 40725 10184
rect 40683 10135 40725 10144
rect 40203 9932 40245 9941
rect 40203 9892 40204 9932
rect 40244 9892 40245 9932
rect 40203 9883 40245 9892
rect 40011 9848 40053 9857
rect 40011 9808 40012 9848
rect 40052 9808 40053 9848
rect 40011 9799 40053 9808
rect 39339 9428 39381 9437
rect 39339 9388 39340 9428
rect 39380 9388 39381 9428
rect 39339 9379 39381 9388
rect 39340 9294 39380 9379
rect 39915 8588 39957 8597
rect 39915 8548 39916 8588
rect 39956 8548 39957 8588
rect 39915 8539 39957 8548
rect 39627 8420 39669 8429
rect 39627 8380 39628 8420
rect 39668 8380 39669 8420
rect 39627 8371 39669 8380
rect 39436 7916 39476 7925
rect 39243 7496 39285 7505
rect 39243 7456 39244 7496
rect 39284 7456 39285 7496
rect 39243 7447 39285 7456
rect 39148 7244 39188 7253
rect 38667 6824 38709 6833
rect 38667 6784 38668 6824
rect 38708 6784 38709 6824
rect 38667 6775 38709 6784
rect 38668 6665 38708 6775
rect 38667 6656 38709 6665
rect 38667 6616 38668 6656
rect 38708 6616 38709 6656
rect 38667 6607 38709 6616
rect 38668 6404 38708 6607
rect 38763 6488 38805 6497
rect 38763 6448 38764 6488
rect 38804 6448 38805 6488
rect 38763 6439 38805 6448
rect 38668 6355 38708 6364
rect 38764 6354 38804 6439
rect 39148 6413 39188 7204
rect 39339 7076 39381 7085
rect 39339 7036 39340 7076
rect 39380 7036 39381 7076
rect 39339 7027 39381 7036
rect 38860 6404 38900 6413
rect 38860 6329 38900 6364
rect 39147 6404 39189 6413
rect 39147 6364 39148 6404
rect 39188 6364 39189 6404
rect 39147 6355 39189 6364
rect 39340 6404 39380 7027
rect 39436 6917 39476 7876
rect 39532 7916 39572 7925
rect 39532 7337 39572 7876
rect 39531 7328 39573 7337
rect 39531 7288 39532 7328
rect 39572 7288 39573 7328
rect 39531 7279 39573 7288
rect 39435 6908 39477 6917
rect 39435 6868 39436 6908
rect 39476 6868 39477 6908
rect 39435 6859 39477 6868
rect 39340 6355 39380 6364
rect 38283 6280 38284 6320
rect 38324 6280 38325 6320
rect 38283 6271 38325 6280
rect 38476 6280 38612 6320
rect 38859 6320 38901 6329
rect 38859 6280 38860 6320
rect 38900 6280 38901 6320
rect 38188 6236 38228 6245
rect 38188 6077 38228 6196
rect 38187 6068 38229 6077
rect 38187 6028 38188 6068
rect 38228 6028 38229 6068
rect 38187 6019 38229 6028
rect 38092 5732 38132 5743
rect 38092 5657 38132 5692
rect 38091 5648 38133 5657
rect 38091 5608 38092 5648
rect 38132 5608 38133 5648
rect 38091 5599 38133 5608
rect 38092 5480 38132 5489
rect 38092 5321 38132 5440
rect 38091 5312 38133 5321
rect 38091 5272 38092 5312
rect 38132 5272 38133 5312
rect 38091 5263 38133 5272
rect 38476 5060 38516 6280
rect 38859 6271 38901 6280
rect 38860 6152 38900 6271
rect 38764 6112 38900 6152
rect 38764 5741 38804 6112
rect 38955 6068 38997 6077
rect 38955 6028 38956 6068
rect 38996 6028 38997 6068
rect 38955 6019 38997 6028
rect 38571 5732 38613 5741
rect 38571 5692 38572 5732
rect 38612 5692 38613 5732
rect 38571 5683 38613 5692
rect 38763 5732 38805 5741
rect 38763 5692 38764 5732
rect 38804 5692 38805 5732
rect 38763 5683 38805 5692
rect 38572 5598 38612 5683
rect 38571 5480 38613 5489
rect 38571 5440 38572 5480
rect 38612 5440 38613 5480
rect 38571 5431 38613 5440
rect 37940 4936 38036 4976
rect 38188 5020 38516 5060
rect 37900 4927 37940 4936
rect 38188 4892 38228 5020
rect 37996 4852 38228 4892
rect 38284 4892 38324 4901
rect 37996 4808 38036 4852
rect 37900 4768 38036 4808
rect 37803 4388 37845 4397
rect 37803 4348 37804 4388
rect 37844 4348 37845 4388
rect 37803 4339 37845 4348
rect 37803 4220 37845 4229
rect 37803 4180 37804 4220
rect 37844 4180 37845 4220
rect 37803 4171 37845 4180
rect 37804 4086 37844 4171
rect 37803 3968 37845 3977
rect 37803 3928 37804 3968
rect 37844 3928 37845 3968
rect 37803 3919 37845 3928
rect 37804 3834 37844 3919
rect 37900 3464 37940 4768
rect 38092 4724 38132 4733
rect 37995 4556 38037 4565
rect 37995 4516 37996 4556
rect 38036 4516 38037 4556
rect 37995 4507 38037 4516
rect 37996 4220 38036 4507
rect 37996 3725 38036 4180
rect 37995 3716 38037 3725
rect 37995 3676 37996 3716
rect 38036 3676 38037 3716
rect 37995 3667 38037 3676
rect 37996 3464 38036 3473
rect 37900 3424 37996 3464
rect 37996 3415 38036 3424
rect 37804 3212 37844 3221
rect 37844 3172 38036 3212
rect 37804 3163 37844 3172
rect 37708 2500 37940 2540
rect 37707 2036 37749 2045
rect 37707 1996 37708 2036
rect 37748 1996 37749 2036
rect 37707 1987 37749 1996
rect 37515 1700 37557 1709
rect 37515 1660 37516 1700
rect 37556 1660 37557 1700
rect 37515 1651 37557 1660
rect 37419 1616 37461 1625
rect 37419 1576 37420 1616
rect 37460 1576 37461 1616
rect 37419 1567 37461 1576
rect 37516 80 37556 1651
rect 37708 80 37748 1987
rect 37900 80 37940 2500
rect 37996 1709 38036 3172
rect 38092 2381 38132 4684
rect 38187 4220 38229 4229
rect 38187 4180 38188 4220
rect 38228 4180 38229 4220
rect 38187 4171 38229 4180
rect 38188 4086 38228 4171
rect 38187 3968 38229 3977
rect 38187 3928 38188 3968
rect 38228 3928 38229 3968
rect 38187 3919 38229 3928
rect 38188 3834 38228 3919
rect 38188 3212 38228 3221
rect 38091 2372 38133 2381
rect 38091 2332 38092 2372
rect 38132 2332 38133 2372
rect 38091 2323 38133 2332
rect 38188 1793 38228 3172
rect 38284 3053 38324 4852
rect 38476 4892 38516 4901
rect 38379 4724 38421 4733
rect 38379 4684 38380 4724
rect 38420 4684 38421 4724
rect 38379 4675 38421 4684
rect 38380 4590 38420 4675
rect 38380 4220 38420 4229
rect 38476 4220 38516 4852
rect 38572 4472 38612 5431
rect 38668 4892 38708 4903
rect 38668 4817 38708 4852
rect 38860 4892 38900 4901
rect 38667 4808 38709 4817
rect 38667 4768 38668 4808
rect 38708 4768 38709 4808
rect 38667 4759 38709 4768
rect 38764 4724 38804 4733
rect 38572 4432 38708 4472
rect 38572 4229 38612 4314
rect 38571 4220 38613 4229
rect 38420 4180 38423 4220
rect 38476 4180 38572 4220
rect 38612 4180 38613 4220
rect 38380 4171 38423 4180
rect 38571 4171 38613 4180
rect 38383 4136 38423 4171
rect 38383 4096 38516 4136
rect 38476 3800 38516 4096
rect 38571 4052 38613 4061
rect 38571 4012 38572 4052
rect 38612 4012 38613 4052
rect 38571 4003 38613 4012
rect 38572 3918 38612 4003
rect 38668 3977 38708 4432
rect 38764 4397 38804 4684
rect 38763 4388 38805 4397
rect 38763 4348 38764 4388
rect 38804 4348 38805 4388
rect 38763 4339 38805 4348
rect 38764 4220 38804 4231
rect 38860 4220 38900 4852
rect 38956 4565 38996 6019
rect 39147 5900 39189 5909
rect 39147 5860 39148 5900
rect 39188 5860 39189 5900
rect 39147 5851 39189 5860
rect 39148 5741 39188 5851
rect 39147 5732 39189 5741
rect 39147 5692 39148 5732
rect 39188 5692 39189 5732
rect 39147 5683 39189 5692
rect 39340 5732 39380 5743
rect 39051 5648 39093 5657
rect 39051 5608 39052 5648
rect 39092 5608 39093 5648
rect 39051 5599 39093 5608
rect 39052 4892 39092 5599
rect 39148 5598 39188 5683
rect 39340 5657 39380 5692
rect 39244 5648 39284 5657
rect 39244 5060 39284 5608
rect 39339 5648 39381 5657
rect 39339 5608 39340 5648
rect 39380 5608 39381 5648
rect 39339 5599 39381 5608
rect 39532 5480 39572 5489
rect 39052 4843 39092 4852
rect 39148 5020 39284 5060
rect 39436 5440 39532 5480
rect 38955 4556 38997 4565
rect 38955 4516 38956 4556
rect 38996 4516 38997 4556
rect 38955 4507 38997 4516
rect 39148 4388 39188 5020
rect 39244 4892 39284 4901
rect 39339 4892 39381 4901
rect 39284 4852 39340 4892
rect 39380 4852 39381 4892
rect 39244 4843 39284 4852
rect 39339 4843 39381 4852
rect 39148 4348 39284 4388
rect 38955 4220 38997 4229
rect 39148 4220 39188 4229
rect 38860 4180 38956 4220
rect 38996 4180 38997 4220
rect 38764 4145 38804 4180
rect 38955 4171 38997 4180
rect 39052 4180 39148 4220
rect 38763 4136 38805 4145
rect 38763 4096 38764 4136
rect 38804 4096 38805 4136
rect 38763 4087 38805 4096
rect 38956 4086 38996 4171
rect 38667 3968 38709 3977
rect 38667 3928 38668 3968
rect 38708 3928 38709 3968
rect 38667 3919 38709 3928
rect 38956 3968 38996 3977
rect 38475 3760 38516 3800
rect 38763 3800 38805 3809
rect 38763 3760 38764 3800
rect 38804 3760 38805 3800
rect 38475 3716 38515 3760
rect 38763 3751 38805 3760
rect 38475 3676 38516 3716
rect 38379 3464 38421 3473
rect 38379 3424 38380 3464
rect 38420 3424 38421 3464
rect 38379 3415 38421 3424
rect 38380 3330 38420 3415
rect 38283 3044 38325 3053
rect 38283 3004 38284 3044
rect 38324 3004 38325 3044
rect 38283 2995 38325 3004
rect 38476 2969 38516 3676
rect 38764 3464 38804 3751
rect 38956 3473 38996 3928
rect 39052 3641 39092 4180
rect 39148 4171 39188 4180
rect 39051 3632 39093 3641
rect 39051 3592 39052 3632
rect 39092 3592 39093 3632
rect 39051 3583 39093 3592
rect 38764 3415 38804 3424
rect 38955 3464 38997 3473
rect 38955 3424 38956 3464
rect 38996 3424 38997 3464
rect 38955 3415 38997 3424
rect 38859 3380 38901 3389
rect 38859 3340 38860 3380
rect 38900 3340 38901 3380
rect 38859 3331 38901 3340
rect 38572 3212 38612 3221
rect 38475 2960 38517 2969
rect 38475 2920 38476 2960
rect 38516 2920 38517 2960
rect 38475 2911 38517 2920
rect 38475 2372 38517 2381
rect 38475 2332 38476 2372
rect 38516 2332 38517 2372
rect 38475 2323 38517 2332
rect 38283 2120 38325 2129
rect 38283 2080 38284 2120
rect 38324 2080 38325 2120
rect 38283 2071 38325 2080
rect 38187 1784 38229 1793
rect 38187 1744 38188 1784
rect 38228 1744 38229 1784
rect 38187 1735 38229 1744
rect 37995 1700 38037 1709
rect 37995 1660 37996 1700
rect 38036 1660 38037 1700
rect 37995 1651 38037 1660
rect 38091 104 38133 113
rect 38091 80 38092 104
rect 824 0 904 80
rect 1016 0 1096 80
rect 1208 0 1288 80
rect 1400 0 1480 80
rect 1592 0 1672 80
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 0 33544 80
rect 33656 0 33736 80
rect 33848 0 33928 80
rect 34040 0 34120 80
rect 34232 0 34312 80
rect 34424 0 34504 80
rect 34616 0 34696 80
rect 34808 0 34888 80
rect 35000 0 35080 80
rect 35192 0 35272 80
rect 35384 0 35464 80
rect 35576 0 35656 80
rect 35768 0 35848 80
rect 35960 0 36040 80
rect 36152 0 36232 80
rect 36344 0 36424 80
rect 36536 0 36616 80
rect 36728 0 36808 80
rect 36920 0 37000 80
rect 37112 0 37192 80
rect 37304 0 37384 80
rect 37496 0 37576 80
rect 37688 0 37768 80
rect 37880 0 37960 80
rect 38072 64 38092 80
rect 38132 80 38133 104
rect 38284 80 38324 2071
rect 38476 80 38516 2323
rect 38572 1541 38612 3172
rect 38571 1532 38613 1541
rect 38571 1492 38572 1532
rect 38612 1492 38613 1532
rect 38571 1483 38613 1492
rect 38667 1448 38709 1457
rect 38667 1408 38668 1448
rect 38708 1408 38709 1448
rect 38667 1399 38709 1408
rect 38668 80 38708 1399
rect 38860 80 38900 3331
rect 38956 3212 38996 3221
rect 38956 1121 38996 3172
rect 39052 2885 39092 3583
rect 39148 3464 39188 3473
rect 39148 3137 39188 3424
rect 39147 3128 39189 3137
rect 39147 3088 39148 3128
rect 39188 3088 39189 3128
rect 39147 3079 39189 3088
rect 39051 2876 39093 2885
rect 39051 2836 39052 2876
rect 39092 2836 39093 2876
rect 39051 2827 39093 2836
rect 39244 2801 39284 4348
rect 39340 4229 39380 4843
rect 39339 4220 39381 4229
rect 39339 4180 39340 4220
rect 39380 4180 39381 4220
rect 39339 4171 39381 4180
rect 39340 4086 39380 4171
rect 39339 3968 39381 3977
rect 39339 3928 39340 3968
rect 39380 3928 39381 3968
rect 39339 3919 39381 3928
rect 39340 3834 39380 3919
rect 39340 3212 39380 3221
rect 39243 2792 39285 2801
rect 39243 2752 39244 2792
rect 39284 2752 39285 2792
rect 39243 2743 39285 2752
rect 39243 1616 39285 1625
rect 39243 1576 39244 1616
rect 39284 1576 39285 1616
rect 39243 1567 39285 1576
rect 39051 1196 39093 1205
rect 39051 1156 39052 1196
rect 39092 1156 39093 1196
rect 39051 1147 39093 1156
rect 38955 1112 38997 1121
rect 38955 1072 38956 1112
rect 38996 1072 38997 1112
rect 38955 1063 38997 1072
rect 39052 80 39092 1147
rect 39244 80 39284 1567
rect 39340 617 39380 3172
rect 39339 608 39381 617
rect 39339 568 39340 608
rect 39380 568 39381 608
rect 39339 559 39381 568
rect 39436 80 39476 5440
rect 39532 5431 39572 5440
rect 39628 5228 39668 8371
rect 39723 8084 39765 8093
rect 39723 8044 39724 8084
rect 39764 8044 39765 8084
rect 39723 8035 39765 8044
rect 39724 7916 39764 8035
rect 39724 7867 39764 7876
rect 39916 7916 39956 8539
rect 39916 7867 39956 7876
rect 39723 7748 39765 7757
rect 39723 7708 39724 7748
rect 39764 7708 39765 7748
rect 39723 7699 39765 7708
rect 39724 7614 39764 7699
rect 39724 5648 39764 5657
rect 39724 5405 39764 5608
rect 39916 5480 39956 5489
rect 39723 5396 39765 5405
rect 39723 5356 39724 5396
rect 39764 5356 39765 5396
rect 39723 5347 39765 5356
rect 39532 5188 39668 5228
rect 39819 5228 39861 5237
rect 39819 5188 39820 5228
rect 39860 5188 39861 5228
rect 39532 4149 39572 5188
rect 39819 5179 39861 5188
rect 39627 4892 39669 4901
rect 39627 4852 39628 4892
rect 39668 4852 39669 4892
rect 39627 4843 39669 4852
rect 39820 4892 39860 5179
rect 39628 4758 39668 4843
rect 39724 4724 39764 4733
rect 39724 4136 39764 4684
rect 39820 4481 39860 4852
rect 39819 4472 39861 4481
rect 39819 4432 39820 4472
rect 39860 4432 39861 4472
rect 39819 4423 39861 4432
rect 39916 4304 39956 5440
rect 39532 4100 39572 4109
rect 39628 4096 39764 4136
rect 39820 4264 39956 4304
rect 39628 4052 39668 4096
rect 39532 4012 39668 4052
rect 39532 3641 39572 4012
rect 39724 3968 39764 3977
rect 39628 3928 39724 3968
rect 39531 3632 39573 3641
rect 39531 3592 39532 3632
rect 39572 3592 39573 3632
rect 39531 3583 39573 3592
rect 39532 3464 39572 3473
rect 39532 3305 39572 3424
rect 39531 3296 39573 3305
rect 39531 3256 39532 3296
rect 39572 3256 39573 3296
rect 39531 3247 39573 3256
rect 39531 1700 39573 1709
rect 39531 1660 39532 1700
rect 39572 1660 39573 1700
rect 39531 1651 39573 1660
rect 39532 1112 39572 1651
rect 39628 1289 39668 3928
rect 39724 3919 39764 3928
rect 39724 3212 39764 3221
rect 39724 1625 39764 3172
rect 39723 1616 39765 1625
rect 39723 1576 39724 1616
rect 39764 1576 39765 1616
rect 39723 1567 39765 1576
rect 39627 1280 39669 1289
rect 39627 1240 39628 1280
rect 39668 1240 39669 1280
rect 39627 1231 39669 1240
rect 39532 1072 39668 1112
rect 39628 80 39668 1072
rect 39820 80 39860 4264
rect 39916 4136 39956 4145
rect 40012 4136 40052 9799
rect 40204 7832 40244 9883
rect 40684 9512 40724 10135
rect 40684 9463 40724 9472
rect 40300 9428 40340 9439
rect 40300 9353 40340 9388
rect 40299 9344 40341 9353
rect 40299 9304 40300 9344
rect 40340 9304 40341 9344
rect 40299 9295 40341 9304
rect 40587 8756 40629 8765
rect 40587 8716 40588 8756
rect 40628 8716 40629 8756
rect 40587 8707 40629 8716
rect 40395 8000 40437 8009
rect 40395 7960 40396 8000
rect 40436 7960 40437 8000
rect 40395 7951 40437 7960
rect 40204 7792 40340 7832
rect 40107 7244 40149 7253
rect 40107 7204 40108 7244
rect 40148 7204 40149 7244
rect 40107 7195 40149 7204
rect 40108 7110 40148 7195
rect 40203 6656 40245 6665
rect 40203 6616 40204 6656
rect 40244 6616 40245 6656
rect 40203 6607 40245 6616
rect 40204 6404 40244 6607
rect 40204 6355 40244 6364
rect 40108 5648 40148 5657
rect 40108 4649 40148 5608
rect 40204 4976 40244 4985
rect 40300 4976 40340 7792
rect 40396 7244 40436 7951
rect 40396 7195 40436 7204
rect 40244 4936 40340 4976
rect 40588 4976 40628 8707
rect 40780 8168 40820 10891
rect 41259 10688 41301 10697
rect 41259 10648 41260 10688
rect 41300 10648 41301 10688
rect 41259 10639 41301 10648
rect 48651 10688 48693 10697
rect 48651 10648 48652 10688
rect 48692 10648 48693 10688
rect 48651 10639 48693 10648
rect 40875 8504 40917 8513
rect 40875 8464 40876 8504
rect 40916 8464 40917 8504
rect 40875 8455 40917 8464
rect 40204 4927 40244 4936
rect 40588 4927 40628 4936
rect 40684 8128 40820 8168
rect 40396 4724 40436 4733
rect 40107 4640 40149 4649
rect 40107 4600 40108 4640
rect 40148 4600 40149 4640
rect 40107 4591 40149 4600
rect 39956 4096 40052 4136
rect 40299 4136 40341 4145
rect 40299 4096 40300 4136
rect 40340 4096 40341 4136
rect 39916 4087 39956 4096
rect 40299 4087 40341 4096
rect 40300 4002 40340 4087
rect 40108 3968 40148 3977
rect 40148 3928 40244 3968
rect 40108 3919 40148 3928
rect 39916 3464 39956 3473
rect 39916 3221 39956 3424
rect 39915 3212 39957 3221
rect 39915 3172 39916 3212
rect 39956 3172 39957 3212
rect 39915 3163 39957 3172
rect 40108 3212 40148 3221
rect 40011 1784 40053 1793
rect 40011 1744 40012 1784
rect 40052 1744 40053 1784
rect 40011 1735 40053 1744
rect 40012 80 40052 1735
rect 40108 1709 40148 3172
rect 40204 1952 40244 3928
rect 40299 3800 40341 3809
rect 40299 3760 40300 3800
rect 40340 3760 40341 3800
rect 40299 3751 40341 3760
rect 40300 3464 40340 3751
rect 40300 3415 40340 3424
rect 40204 1912 40340 1952
rect 40107 1700 40149 1709
rect 40107 1660 40108 1700
rect 40148 1660 40149 1700
rect 40107 1651 40149 1660
rect 40203 1532 40245 1541
rect 40203 1492 40204 1532
rect 40244 1492 40245 1532
rect 40203 1483 40245 1492
rect 40204 80 40244 1483
rect 40300 1205 40340 1912
rect 40299 1196 40341 1205
rect 40299 1156 40300 1196
rect 40340 1156 40341 1196
rect 40299 1147 40341 1156
rect 40396 80 40436 4684
rect 40587 4136 40629 4145
rect 40587 4096 40588 4136
rect 40628 4096 40629 4136
rect 40587 4087 40629 4096
rect 40684 4136 40724 8128
rect 40876 7916 40916 8455
rect 40876 7867 40916 7876
rect 41163 7916 41205 7925
rect 41163 7876 41164 7916
rect 41204 7876 41205 7916
rect 41163 7867 41205 7876
rect 41164 7782 41204 7867
rect 40780 6320 40820 6329
rect 41260 6320 41300 10639
rect 41547 10436 41589 10445
rect 41547 10396 41548 10436
rect 41588 10396 41589 10436
rect 41547 10387 41589 10396
rect 41548 10268 41588 10387
rect 48652 10277 48692 10639
rect 49803 10436 49845 10445
rect 49803 10396 49804 10436
rect 49844 10396 49845 10436
rect 49803 10387 49845 10396
rect 49419 10352 49461 10361
rect 49419 10312 49420 10352
rect 49460 10312 49461 10352
rect 49419 10303 49461 10312
rect 41548 10219 41588 10228
rect 41836 10268 41876 10277
rect 41836 10109 41876 10228
rect 42795 10268 42837 10277
rect 42795 10228 42796 10268
rect 42836 10228 42837 10268
rect 42795 10219 42837 10228
rect 48651 10268 48693 10277
rect 48651 10228 48652 10268
rect 48692 10228 48693 10268
rect 48651 10219 48693 10228
rect 42796 10134 42836 10219
rect 41835 10100 41877 10109
rect 41835 10060 41836 10100
rect 41876 10060 41877 10100
rect 41835 10051 41877 10060
rect 42315 9764 42357 9773
rect 42315 9724 42316 9764
rect 42356 9724 42357 9764
rect 42315 9715 42357 9724
rect 46251 9764 46293 9773
rect 46251 9724 46252 9764
rect 46292 9724 46293 9764
rect 46251 9715 46293 9724
rect 41548 9428 41588 9437
rect 41548 9017 41588 9388
rect 42316 9428 42356 9715
rect 43659 9680 43701 9689
rect 43659 9640 43660 9680
rect 43700 9640 43701 9680
rect 43659 9631 43701 9640
rect 43083 9596 43125 9605
rect 43083 9556 43084 9596
rect 43124 9556 43125 9596
rect 43083 9547 43125 9556
rect 42316 9379 42356 9388
rect 42699 9176 42741 9185
rect 42699 9136 42700 9176
rect 42740 9136 42741 9176
rect 42699 9127 42741 9136
rect 41547 9008 41589 9017
rect 41547 8968 41548 9008
rect 41588 8968 41589 9008
rect 41547 8959 41589 8968
rect 42507 8672 42549 8681
rect 42507 8632 42508 8672
rect 42548 8632 42549 8672
rect 42507 8623 42549 8632
rect 42508 8538 42548 8623
rect 42411 8420 42453 8429
rect 42411 8380 42412 8420
rect 42452 8380 42453 8420
rect 42411 8371 42453 8380
rect 42028 7916 42068 7925
rect 41355 7748 41397 7757
rect 41355 7708 41356 7748
rect 41396 7708 41397 7748
rect 41355 7699 41397 7708
rect 41356 7244 41396 7699
rect 42028 7673 42068 7876
rect 42123 7916 42165 7925
rect 42123 7876 42124 7916
rect 42164 7876 42165 7916
rect 42123 7867 42165 7876
rect 42412 7916 42452 8371
rect 42412 7867 42452 7876
rect 42027 7664 42069 7673
rect 42027 7624 42028 7664
rect 42068 7624 42069 7664
rect 42027 7615 42069 7624
rect 41356 7195 41396 7204
rect 41931 7160 41973 7169
rect 41931 7120 41932 7160
rect 41972 7120 41973 7160
rect 41931 7111 41973 7120
rect 41739 6824 41781 6833
rect 41739 6784 41740 6824
rect 41780 6784 41781 6824
rect 41739 6775 41781 6784
rect 41644 6413 41684 6498
rect 41643 6404 41685 6413
rect 41643 6364 41644 6404
rect 41684 6364 41685 6404
rect 41643 6355 41685 6364
rect 41260 6280 41396 6320
rect 40780 5741 40820 6280
rect 41259 5984 41301 5993
rect 41259 5944 41260 5984
rect 41300 5944 41301 5984
rect 41259 5935 41301 5944
rect 40779 5732 40821 5741
rect 40779 5692 40780 5732
rect 40820 5692 40821 5732
rect 40779 5683 40821 5692
rect 41260 5648 41300 5935
rect 41260 5599 41300 5608
rect 41068 5480 41108 5489
rect 40875 5228 40917 5237
rect 40875 5188 40876 5228
rect 40916 5188 40917 5228
rect 40875 5179 40917 5188
rect 40684 4087 40724 4096
rect 40780 4724 40820 4733
rect 40492 3968 40532 3977
rect 40492 3389 40532 3928
rect 40588 3557 40628 4087
rect 40587 3548 40629 3557
rect 40587 3508 40588 3548
rect 40628 3508 40629 3548
rect 40587 3499 40629 3508
rect 40684 3464 40724 3473
rect 40491 3380 40533 3389
rect 40491 3340 40492 3380
rect 40532 3340 40533 3380
rect 40491 3331 40533 3340
rect 40684 3305 40724 3424
rect 40683 3296 40725 3305
rect 40683 3256 40684 3296
rect 40724 3256 40725 3296
rect 40683 3247 40725 3256
rect 40492 3212 40532 3221
rect 40492 785 40532 3172
rect 40780 2381 40820 4684
rect 40876 4145 40916 5179
rect 40971 5060 41013 5069
rect 40971 5020 40972 5060
rect 41012 5020 41013 5060
rect 40971 5011 41013 5020
rect 40972 4976 41012 5011
rect 40972 4925 41012 4936
rect 41068 4304 41108 5440
rect 41356 4976 41396 6280
rect 41740 5816 41780 6775
rect 41932 6404 41972 7111
rect 41932 6355 41972 6364
rect 41740 5767 41780 5776
rect 41739 5480 41781 5489
rect 41739 5440 41740 5480
rect 41780 5440 41781 5480
rect 41739 5431 41781 5440
rect 41547 5060 41589 5069
rect 41547 5020 41548 5060
rect 41588 5020 41589 5060
rect 41547 5011 41589 5020
rect 41356 4927 41396 4936
rect 41548 4926 41588 5011
rect 41740 4976 41780 5431
rect 41740 4927 41780 4936
rect 40972 4264 41108 4304
rect 41164 4724 41204 4733
rect 40875 4136 40917 4145
rect 40875 4096 40876 4136
rect 40916 4096 40917 4136
rect 40875 4087 40917 4096
rect 40876 3968 40916 3977
rect 40876 3557 40916 3928
rect 40875 3548 40917 3557
rect 40875 3508 40876 3548
rect 40916 3508 40917 3548
rect 40875 3499 40917 3508
rect 40876 3212 40916 3221
rect 40779 2372 40821 2381
rect 40779 2332 40780 2372
rect 40820 2332 40821 2372
rect 40779 2323 40821 2332
rect 40876 1457 40916 3172
rect 40875 1448 40917 1457
rect 40875 1408 40876 1448
rect 40916 1408 40917 1448
rect 40875 1399 40917 1408
rect 40779 1280 40821 1289
rect 40779 1240 40780 1280
rect 40820 1240 40821 1280
rect 40779 1231 40821 1240
rect 40587 1112 40629 1121
rect 40587 1072 40588 1112
rect 40628 1072 40629 1112
rect 40587 1063 40629 1072
rect 40491 776 40533 785
rect 40491 736 40492 776
rect 40532 736 40533 776
rect 40491 727 40533 736
rect 40588 80 40628 1063
rect 40780 80 40820 1231
rect 40972 80 41012 4264
rect 41067 4136 41109 4145
rect 41067 4096 41068 4136
rect 41108 4096 41109 4136
rect 41067 4087 41109 4096
rect 41068 4002 41108 4087
rect 41067 3800 41109 3809
rect 41067 3760 41068 3800
rect 41108 3760 41109 3800
rect 41067 3751 41109 3760
rect 41068 3464 41108 3751
rect 41068 3415 41108 3424
rect 41164 2549 41204 4684
rect 41835 4724 41877 4733
rect 41835 4684 41836 4724
rect 41876 4684 41877 4724
rect 41835 4675 41877 4684
rect 41932 4724 41972 4733
rect 41355 4388 41397 4397
rect 41355 4348 41356 4388
rect 41396 4348 41397 4388
rect 41355 4339 41397 4348
rect 41260 3968 41300 3977
rect 41260 3809 41300 3928
rect 41356 3884 41396 4339
rect 41451 4136 41493 4145
rect 41451 4096 41452 4136
rect 41492 4096 41493 4136
rect 41451 4087 41493 4096
rect 41836 4136 41876 4675
rect 41836 4087 41876 4096
rect 41452 4002 41492 4087
rect 41644 3968 41684 3977
rect 41684 3928 41780 3968
rect 41644 3919 41684 3928
rect 41356 3844 41492 3884
rect 41259 3800 41301 3809
rect 41259 3760 41260 3800
rect 41300 3760 41301 3800
rect 41259 3751 41301 3760
rect 41355 3548 41397 3557
rect 41355 3508 41356 3548
rect 41396 3508 41397 3548
rect 41355 3499 41397 3508
rect 41260 3212 41300 3221
rect 41163 2540 41205 2549
rect 41163 2500 41164 2540
rect 41204 2500 41205 2540
rect 41163 2491 41205 2500
rect 41163 2372 41205 2381
rect 41163 2332 41164 2372
rect 41204 2332 41205 2372
rect 41163 2323 41205 2332
rect 41164 80 41204 2323
rect 41260 365 41300 3172
rect 41356 2045 41396 3499
rect 41452 3464 41492 3844
rect 41452 3415 41492 3424
rect 41644 3212 41684 3221
rect 41547 3128 41589 3137
rect 41547 3088 41548 3128
rect 41588 3088 41589 3128
rect 41547 3079 41589 3088
rect 41548 2717 41588 3079
rect 41547 2708 41589 2717
rect 41547 2668 41548 2708
rect 41588 2668 41589 2708
rect 41547 2659 41589 2668
rect 41355 2036 41397 2045
rect 41355 1996 41356 2036
rect 41396 1996 41397 2036
rect 41355 1987 41397 1996
rect 41547 1196 41589 1205
rect 41547 1156 41548 1196
rect 41588 1156 41589 1196
rect 41547 1147 41589 1156
rect 41355 608 41397 617
rect 41355 568 41356 608
rect 41396 568 41397 608
rect 41355 559 41397 568
rect 41259 356 41301 365
rect 41259 316 41260 356
rect 41300 316 41301 356
rect 41259 307 41301 316
rect 41356 80 41396 559
rect 41548 80 41588 1147
rect 41644 953 41684 3172
rect 41740 2717 41780 3928
rect 41835 3464 41877 3473
rect 41835 3424 41836 3464
rect 41876 3424 41877 3464
rect 41835 3415 41877 3424
rect 41836 3330 41876 3415
rect 41739 2708 41781 2717
rect 41739 2668 41740 2708
rect 41780 2668 41781 2708
rect 41739 2659 41781 2668
rect 41932 2549 41972 4684
rect 42124 4136 42164 7867
rect 42604 5732 42644 5741
rect 42604 5405 42644 5692
rect 42603 5396 42645 5405
rect 42603 5356 42604 5396
rect 42644 5356 42645 5396
rect 42603 5347 42645 5356
rect 42700 5153 42740 9127
rect 42987 7412 43029 7421
rect 42987 7372 42988 7412
rect 43028 7372 43029 7412
rect 42987 7363 43029 7372
rect 42988 7278 43028 7363
rect 42891 7076 42933 7085
rect 42891 7036 42892 7076
rect 42932 7036 42933 7076
rect 42891 7027 42933 7036
rect 42796 6404 42836 6413
rect 42892 6404 42932 7027
rect 42836 6364 42932 6404
rect 42796 6355 42836 6364
rect 43084 6320 43124 9547
rect 43276 9428 43316 9439
rect 43276 9353 43316 9388
rect 43275 9344 43317 9353
rect 43275 9304 43276 9344
rect 43316 9304 43317 9344
rect 43275 9295 43317 9304
rect 43371 8756 43413 8765
rect 43371 8716 43372 8756
rect 43412 8716 43413 8756
rect 43371 8707 43413 8716
rect 43660 8756 43700 9631
rect 43755 9092 43797 9101
rect 43755 9052 43756 9092
rect 43796 9052 43797 9092
rect 43755 9043 43797 9052
rect 43660 8707 43700 8716
rect 43372 8622 43412 8707
rect 43371 7916 43413 7925
rect 43371 7876 43372 7916
rect 43412 7876 43413 7916
rect 43371 7867 43413 7876
rect 43372 7782 43412 7867
rect 43467 7244 43509 7253
rect 43467 7204 43468 7244
rect 43508 7204 43509 7244
rect 43467 7195 43509 7204
rect 43468 7110 43508 7195
rect 43467 6572 43509 6581
rect 43467 6532 43468 6572
rect 43508 6532 43509 6572
rect 43467 6523 43509 6532
rect 43468 6404 43508 6523
rect 43468 6355 43508 6364
rect 42892 6280 43124 6320
rect 42892 5648 42932 6280
rect 42892 5599 42932 5608
rect 43275 5648 43317 5657
rect 43275 5608 43276 5648
rect 43316 5608 43317 5648
rect 43275 5599 43317 5608
rect 43659 5648 43701 5657
rect 43659 5608 43660 5648
rect 43700 5608 43701 5648
rect 43659 5599 43701 5608
rect 43276 5514 43316 5599
rect 43660 5514 43700 5599
rect 43084 5480 43124 5489
rect 42699 5144 42741 5153
rect 42699 5104 42700 5144
rect 42740 5104 42741 5144
rect 42699 5095 42741 5104
rect 42507 5060 42549 5069
rect 42507 5020 42508 5060
rect 42548 5020 42549 5060
rect 42507 5011 42549 5020
rect 42987 5060 43029 5069
rect 42987 5020 42988 5060
rect 43028 5020 43029 5060
rect 42987 5011 43029 5020
rect 42219 4808 42261 4817
rect 42219 4768 42220 4808
rect 42260 4768 42261 4808
rect 42219 4759 42261 4768
rect 42220 4674 42260 4759
rect 42220 4136 42260 4145
rect 42124 4096 42220 4136
rect 42220 4087 42260 4096
rect 42028 3968 42068 3977
rect 42412 3968 42452 3977
rect 42028 3557 42068 3928
rect 42316 3928 42412 3968
rect 42219 3884 42261 3893
rect 42219 3844 42220 3884
rect 42260 3844 42261 3884
rect 42219 3835 42261 3844
rect 42027 3548 42069 3557
rect 42027 3508 42028 3548
rect 42068 3508 42069 3548
rect 42027 3499 42069 3508
rect 42220 3464 42260 3835
rect 42220 3415 42260 3424
rect 42123 3380 42165 3389
rect 42123 3340 42124 3380
rect 42164 3340 42165 3380
rect 42123 3331 42165 3340
rect 42028 3212 42068 3221
rect 41739 2540 41781 2549
rect 41739 2500 41740 2540
rect 41780 2500 41781 2540
rect 41739 2491 41781 2500
rect 41931 2540 41973 2549
rect 41931 2500 41932 2540
rect 41972 2500 41973 2540
rect 41931 2491 41973 2500
rect 41643 944 41685 953
rect 41643 904 41644 944
rect 41684 904 41685 944
rect 41643 895 41685 904
rect 41740 80 41780 2491
rect 41931 1616 41973 1625
rect 41931 1576 41932 1616
rect 41972 1576 41973 1616
rect 41931 1567 41973 1576
rect 41932 80 41972 1567
rect 42028 1037 42068 3172
rect 42027 1028 42069 1037
rect 42027 988 42028 1028
rect 42068 988 42069 1028
rect 42027 979 42069 988
rect 42124 80 42164 3331
rect 42219 2708 42261 2717
rect 42219 2668 42220 2708
rect 42260 2668 42261 2708
rect 42219 2659 42261 2668
rect 42220 188 42260 2659
rect 42316 281 42356 3928
rect 42412 3919 42452 3928
rect 42412 3212 42452 3221
rect 42412 1625 42452 3172
rect 42508 2717 42548 5011
rect 42988 4892 43028 5011
rect 42988 4843 43028 4852
rect 42603 4136 42645 4145
rect 42603 4096 42604 4136
rect 42644 4096 42645 4136
rect 42603 4087 42645 4096
rect 42987 4136 43029 4145
rect 42987 4096 42988 4136
rect 43028 4096 43029 4136
rect 42987 4087 43029 4096
rect 42604 4002 42644 4087
rect 42795 4052 42837 4061
rect 42795 4012 42796 4052
rect 42836 4012 42837 4052
rect 42795 4003 42837 4012
rect 42796 3918 42836 4003
rect 42988 4002 43028 4087
rect 42987 3884 43029 3893
rect 42987 3844 42988 3884
rect 43028 3844 43029 3884
rect 42987 3835 43029 3844
rect 42603 3632 42645 3641
rect 42603 3592 42604 3632
rect 42644 3592 42645 3632
rect 42603 3583 42645 3592
rect 42891 3632 42933 3641
rect 42891 3592 42892 3632
rect 42932 3592 42933 3632
rect 42891 3583 42933 3592
rect 42604 3464 42644 3583
rect 42604 3415 42644 3424
rect 42796 3212 42836 3221
rect 42507 2708 42549 2717
rect 42507 2668 42508 2708
rect 42548 2668 42549 2708
rect 42507 2659 42549 2668
rect 42699 2036 42741 2045
rect 42699 1996 42700 2036
rect 42740 1996 42741 2036
rect 42699 1987 42741 1996
rect 42507 1700 42549 1709
rect 42507 1660 42508 1700
rect 42548 1660 42549 1700
rect 42507 1651 42549 1660
rect 42411 1616 42453 1625
rect 42411 1576 42412 1616
rect 42452 1576 42453 1616
rect 42411 1567 42453 1576
rect 42315 272 42357 281
rect 42315 232 42316 272
rect 42356 232 42357 272
rect 42315 223 42357 232
rect 42220 148 42271 188
rect 42231 104 42271 148
rect 42231 80 42356 104
rect 42508 80 42548 1651
rect 42700 80 42740 1987
rect 42796 1289 42836 3172
rect 42892 2969 42932 3583
rect 42988 3464 43028 3835
rect 42988 3415 43028 3424
rect 43084 2969 43124 5440
rect 43468 5480 43508 5489
rect 43508 5440 43604 5480
rect 43468 5431 43508 5440
rect 43468 4808 43508 4817
rect 43371 4136 43413 4145
rect 43371 4096 43372 4136
rect 43412 4096 43413 4136
rect 43371 4087 43413 4096
rect 43372 4002 43412 4087
rect 43179 3968 43221 3977
rect 43179 3928 43180 3968
rect 43220 3928 43221 3968
rect 43179 3919 43221 3928
rect 43180 3834 43220 3919
rect 43275 3800 43317 3809
rect 43275 3760 43276 3800
rect 43316 3760 43317 3800
rect 43275 3751 43317 3760
rect 43180 3212 43220 3221
rect 43180 3053 43220 3172
rect 43179 3044 43221 3053
rect 43179 3004 43180 3044
rect 43220 3004 43221 3044
rect 43179 2995 43221 3004
rect 42891 2960 42933 2969
rect 42891 2920 42892 2960
rect 42932 2920 42933 2960
rect 42891 2911 42933 2920
rect 43083 2960 43125 2969
rect 43083 2920 43084 2960
rect 43124 2920 43125 2960
rect 43083 2911 43125 2920
rect 42891 2540 42933 2549
rect 42891 2500 42892 2540
rect 42932 2500 42933 2540
rect 42891 2491 42933 2500
rect 42795 1280 42837 1289
rect 42795 1240 42796 1280
rect 42836 1240 42837 1280
rect 42795 1231 42837 1240
rect 42892 80 42932 2491
rect 43083 776 43125 785
rect 43083 736 43084 776
rect 43124 736 43125 776
rect 43083 727 43125 736
rect 43084 80 43124 727
rect 43276 80 43316 3751
rect 43468 3725 43508 4768
rect 43564 4136 43604 5440
rect 43564 4096 43700 4136
rect 43564 3968 43604 3977
rect 43564 3809 43604 3928
rect 43563 3800 43605 3809
rect 43563 3760 43564 3800
rect 43604 3760 43605 3800
rect 43563 3751 43605 3760
rect 43467 3716 43509 3725
rect 43467 3676 43468 3716
rect 43508 3676 43509 3716
rect 43467 3667 43509 3676
rect 43371 3464 43413 3473
rect 43371 3424 43372 3464
rect 43412 3424 43413 3464
rect 43371 3415 43413 3424
rect 43372 3330 43412 3415
rect 43564 3212 43604 3221
rect 43467 2960 43509 2969
rect 43467 2920 43468 2960
rect 43508 2920 43509 2960
rect 43467 2911 43509 2920
rect 43468 80 43508 2911
rect 43564 2885 43604 3172
rect 43563 2876 43605 2885
rect 43563 2836 43564 2876
rect 43604 2836 43605 2876
rect 43563 2827 43605 2836
rect 43660 2792 43700 4096
rect 43756 3464 43796 9043
rect 44716 8968 45044 9008
rect 44139 8840 44181 8849
rect 44139 8800 44140 8840
rect 44180 8800 44181 8840
rect 44139 8791 44181 8800
rect 44140 8420 44180 8791
rect 44620 8756 44660 8765
rect 44620 8429 44660 8716
rect 43948 8380 44180 8420
rect 44619 8420 44661 8429
rect 44619 8380 44620 8420
rect 44660 8380 44661 8420
rect 43948 7253 43988 8380
rect 44619 8371 44661 8380
rect 44139 8252 44181 8261
rect 44139 8212 44140 8252
rect 44180 8212 44181 8252
rect 44139 8203 44181 8212
rect 44619 8252 44661 8261
rect 44619 8212 44620 8252
rect 44660 8212 44661 8252
rect 44619 8203 44661 8212
rect 44043 7916 44085 7925
rect 44043 7876 44044 7916
rect 44084 7876 44085 7916
rect 44043 7867 44085 7876
rect 44044 7782 44084 7867
rect 43947 7244 43989 7253
rect 43947 7204 43948 7244
rect 43988 7204 43989 7244
rect 43947 7195 43989 7204
rect 44140 5909 44180 8203
rect 44236 7916 44276 7927
rect 44236 7841 44276 7876
rect 44332 7916 44372 7925
rect 44372 7876 44468 7916
rect 44332 7867 44372 7876
rect 44235 7832 44277 7841
rect 44235 7792 44236 7832
rect 44276 7792 44277 7832
rect 44235 7783 44277 7792
rect 44331 7664 44373 7673
rect 44331 7624 44332 7664
rect 44372 7624 44373 7664
rect 44331 7615 44373 7624
rect 44332 7244 44372 7615
rect 44428 7253 44468 7876
rect 44524 7706 44564 7715
rect 44524 7412 44564 7666
rect 44620 7589 44660 8203
rect 44716 7706 44756 8968
rect 45004 8924 45044 8968
rect 45196 8924 45236 8933
rect 45004 8884 45196 8924
rect 45196 8875 45236 8884
rect 44907 8840 44949 8849
rect 44907 8800 44908 8840
rect 44948 8800 44949 8840
rect 44907 8791 44949 8800
rect 44908 8756 44948 8791
rect 46252 8765 46292 9715
rect 48459 9596 48501 9605
rect 48459 9556 48460 9596
rect 48500 9556 48501 9596
rect 48459 9547 48501 9556
rect 48652 9596 48692 10219
rect 49420 10218 49460 10303
rect 49048 9848 49416 9857
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49048 9799 49416 9808
rect 48652 9547 48692 9556
rect 48939 9596 48981 9605
rect 48939 9556 48940 9596
rect 48980 9556 48981 9596
rect 48939 9547 48981 9556
rect 47595 9512 47637 9521
rect 47595 9472 47596 9512
rect 47636 9472 47637 9512
rect 47595 9463 47637 9472
rect 48268 9512 48308 9521
rect 47019 9260 47061 9269
rect 47019 9220 47020 9260
rect 47060 9220 47061 9260
rect 47019 9211 47061 9220
rect 44908 8705 44948 8716
rect 45100 8756 45140 8765
rect 44907 8588 44949 8597
rect 44907 8548 44908 8588
rect 44948 8548 44949 8588
rect 44907 8539 44949 8548
rect 44619 7580 44661 7589
rect 44619 7540 44620 7580
rect 44660 7540 44661 7580
rect 44619 7531 44661 7540
rect 44620 7412 44660 7421
rect 44716 7412 44756 7666
rect 44524 7372 44620 7412
rect 44660 7372 44756 7412
rect 44620 7363 44660 7372
rect 44332 7195 44372 7204
rect 44427 7244 44469 7253
rect 44524 7245 44564 7254
rect 44427 7204 44428 7244
rect 44468 7205 44524 7244
rect 44468 7204 44564 7205
rect 44427 7195 44469 7204
rect 44524 7196 44564 7204
rect 44620 7244 44660 7253
rect 44523 6992 44565 7001
rect 44620 6992 44660 7204
rect 44236 6952 44524 6992
rect 44564 6952 44660 6992
rect 44139 5900 44181 5909
rect 44139 5860 44140 5900
rect 44180 5860 44181 5900
rect 44139 5851 44181 5860
rect 44044 5732 44084 5741
rect 44044 5489 44084 5692
rect 44236 5732 44276 6952
rect 44523 6943 44565 6952
rect 44524 6858 44564 6943
rect 44716 6824 44756 7372
rect 44908 7916 44948 8539
rect 44908 7253 44948 7876
rect 45003 7916 45045 7925
rect 45003 7876 45004 7916
rect 45044 7876 45045 7916
rect 45003 7867 45045 7876
rect 45004 7782 45044 7867
rect 44907 7244 44949 7253
rect 44907 7204 44908 7244
rect 44948 7204 44949 7244
rect 44907 7195 44949 7204
rect 44620 6784 44756 6824
rect 44427 6488 44469 6497
rect 44427 6448 44428 6488
rect 44468 6448 44469 6488
rect 44427 6439 44469 6448
rect 44332 6404 44372 6413
rect 44332 6077 44372 6364
rect 44331 6068 44373 6077
rect 44331 6028 44332 6068
rect 44372 6028 44373 6068
rect 44331 6019 44373 6028
rect 44331 5816 44373 5825
rect 44331 5776 44332 5816
rect 44372 5776 44373 5816
rect 44331 5767 44373 5776
rect 44236 5683 44276 5692
rect 44332 5732 44372 5767
rect 44332 5681 44372 5692
rect 43852 5480 43892 5489
rect 44043 5480 44085 5489
rect 43892 5440 43988 5480
rect 43852 5431 43892 5440
rect 43756 3415 43796 3424
rect 43948 3389 43988 5440
rect 44043 5440 44044 5480
rect 44084 5440 44085 5480
rect 44043 5431 44085 5440
rect 44236 5480 44276 5489
rect 44139 5228 44181 5237
rect 44139 5188 44140 5228
rect 44180 5188 44181 5228
rect 44139 5179 44181 5188
rect 44140 3464 44180 5179
rect 44236 5069 44276 5440
rect 44235 5060 44277 5069
rect 44235 5020 44236 5060
rect 44276 5020 44277 5060
rect 44235 5011 44277 5020
rect 44332 4892 44372 4901
rect 44332 4649 44372 4852
rect 44331 4640 44373 4649
rect 44331 4600 44332 4640
rect 44372 4600 44373 4640
rect 44331 4591 44373 4600
rect 44140 3415 44180 3424
rect 44236 3968 44276 3977
rect 43947 3380 43989 3389
rect 43947 3340 43948 3380
rect 43988 3340 43989 3380
rect 43947 3331 43989 3340
rect 43948 3212 43988 3221
rect 43948 2969 43988 3172
rect 44236 3137 44276 3928
rect 44331 3548 44373 3557
rect 44331 3508 44332 3548
rect 44372 3508 44373 3548
rect 44331 3499 44373 3508
rect 44332 3380 44372 3499
rect 44428 3464 44468 6439
rect 44524 5732 44564 5760
rect 44620 5732 44660 6784
rect 44716 6413 44756 6498
rect 45100 6497 45140 8716
rect 45196 8756 45236 8765
rect 46156 8756 46196 8765
rect 45196 8597 45236 8716
rect 45868 8716 46156 8756
rect 45195 8588 45237 8597
rect 45195 8548 45196 8588
rect 45236 8548 45237 8588
rect 45195 8539 45237 8548
rect 45387 8000 45429 8009
rect 45196 7960 45388 8000
rect 45428 7960 45429 8000
rect 45196 7916 45236 7960
rect 45387 7951 45429 7960
rect 45579 8000 45621 8009
rect 45579 7960 45580 8000
rect 45620 7960 45621 8000
rect 45579 7951 45621 7960
rect 45196 7867 45236 7876
rect 45580 7757 45620 7951
rect 45868 7925 45908 8716
rect 46156 8707 46196 8716
rect 46251 8756 46293 8765
rect 46251 8716 46252 8756
rect 46292 8716 46293 8756
rect 46251 8707 46293 8716
rect 46252 8084 46292 8707
rect 46539 8588 46581 8597
rect 46539 8548 46540 8588
rect 46580 8548 46581 8588
rect 46539 8539 46581 8548
rect 46252 8035 46292 8044
rect 46540 7925 46580 8539
rect 46923 8504 46965 8513
rect 46923 8464 46924 8504
rect 46964 8464 46965 8504
rect 46923 8455 46965 8464
rect 46924 7925 46964 8455
rect 45772 7916 45812 7925
rect 45579 7748 45621 7757
rect 45579 7708 45580 7748
rect 45620 7708 45621 7748
rect 45579 7699 45621 7708
rect 45772 7589 45812 7876
rect 45867 7916 45909 7925
rect 45867 7876 45868 7916
rect 45908 7876 45909 7916
rect 45867 7867 45909 7876
rect 46155 7916 46197 7925
rect 46155 7876 46156 7916
rect 46196 7876 46197 7916
rect 46155 7867 46197 7876
rect 46444 7916 46484 7925
rect 45867 7748 45909 7757
rect 45867 7708 45868 7748
rect 45908 7708 45909 7748
rect 45867 7699 45909 7708
rect 45291 7580 45333 7589
rect 45291 7540 45292 7580
rect 45332 7540 45333 7580
rect 45291 7531 45333 7540
rect 45771 7580 45813 7589
rect 45771 7540 45772 7580
rect 45812 7540 45813 7580
rect 45771 7531 45813 7540
rect 45195 7244 45237 7253
rect 45195 7204 45196 7244
rect 45236 7204 45237 7244
rect 45195 7195 45237 7204
rect 44811 6488 44853 6497
rect 44811 6448 44812 6488
rect 44852 6448 44853 6488
rect 44811 6439 44853 6448
rect 45099 6488 45141 6497
rect 45099 6448 45100 6488
rect 45140 6448 45141 6488
rect 45099 6439 45141 6448
rect 44715 6404 44757 6413
rect 44715 6364 44716 6404
rect 44756 6364 44757 6404
rect 44715 6355 44757 6364
rect 44715 5816 44757 5825
rect 44715 5776 44716 5816
rect 44756 5776 44757 5816
rect 44715 5767 44757 5776
rect 44564 5692 44660 5732
rect 44524 5683 44564 5692
rect 44620 5489 44660 5692
rect 44716 5732 44756 5767
rect 44716 5681 44756 5692
rect 44812 5732 44852 6439
rect 45099 6152 45141 6161
rect 45099 6112 45100 6152
rect 45140 6112 45141 6152
rect 45099 6103 45141 6112
rect 44812 5683 44852 5692
rect 45100 5732 45140 6103
rect 45196 5825 45236 7195
rect 45195 5816 45237 5825
rect 45195 5776 45196 5816
rect 45236 5776 45237 5816
rect 45195 5767 45237 5776
rect 44524 5480 44564 5489
rect 44524 4649 44564 5440
rect 44619 5480 44661 5489
rect 44619 5440 44620 5480
rect 44660 5440 44661 5480
rect 44619 5431 44661 5440
rect 44716 4808 44756 4817
rect 44523 4640 44565 4649
rect 44523 4600 44524 4640
rect 44564 4600 44565 4640
rect 44523 4591 44565 4600
rect 44619 4220 44661 4229
rect 44619 4180 44620 4220
rect 44660 4180 44661 4220
rect 44619 4171 44661 4180
rect 44620 4086 44660 4171
rect 44716 3473 44756 4768
rect 44524 3464 44564 3473
rect 44428 3424 44524 3464
rect 44524 3415 44564 3424
rect 44715 3464 44757 3473
rect 44715 3424 44716 3464
rect 44756 3424 44757 3464
rect 44715 3415 44757 3424
rect 44908 3464 44948 3473
rect 44619 3380 44661 3389
rect 44332 3340 44468 3380
rect 44332 3212 44372 3221
rect 44235 3128 44277 3137
rect 44235 3088 44236 3128
rect 44276 3088 44277 3128
rect 44235 3079 44277 3088
rect 43947 2960 43989 2969
rect 43947 2920 43948 2960
rect 43988 2920 43989 2960
rect 43947 2911 43989 2920
rect 44332 2801 44372 3172
rect 44331 2792 44373 2801
rect 43660 2752 44084 2792
rect 43851 2624 43893 2633
rect 43851 2584 43852 2624
rect 43892 2584 43893 2624
rect 43851 2575 43893 2584
rect 43659 1448 43701 1457
rect 43659 1408 43660 1448
rect 43700 1408 43701 1448
rect 43659 1399 43701 1408
rect 43660 80 43700 1399
rect 43852 80 43892 2575
rect 44044 80 44084 2752
rect 44331 2752 44332 2792
rect 44372 2752 44373 2792
rect 44331 2743 44373 2752
rect 44235 356 44277 365
rect 44235 316 44236 356
rect 44276 316 44277 356
rect 44235 307 44277 316
rect 44236 80 44276 307
rect 44428 80 44468 3340
rect 44619 3340 44620 3380
rect 44660 3340 44661 3380
rect 44619 3331 44661 3340
rect 44620 80 44660 3331
rect 44716 3212 44756 3221
rect 44716 2633 44756 3172
rect 44715 2624 44757 2633
rect 44715 2584 44716 2624
rect 44756 2584 44757 2624
rect 44715 2575 44757 2584
rect 44908 2465 44948 3424
rect 45100 3389 45140 5692
rect 45196 5732 45236 5767
rect 45196 5681 45236 5692
rect 45292 5657 45332 7531
rect 45772 7244 45812 7253
rect 45676 6413 45716 6498
rect 45675 6404 45717 6413
rect 45675 6364 45676 6404
rect 45716 6364 45717 6404
rect 45675 6355 45717 6364
rect 45772 6320 45812 7204
rect 45868 6404 45908 7699
rect 46156 7664 46196 7867
rect 46156 7624 46292 7664
rect 45963 7412 46005 7421
rect 45963 7372 45964 7412
rect 46004 7372 46005 7412
rect 45963 7363 46005 7372
rect 45964 7244 46004 7363
rect 45964 7195 46004 7204
rect 46156 6404 46196 6413
rect 45868 6364 46004 6404
rect 45772 6280 45908 6320
rect 45675 5984 45717 5993
rect 45675 5944 45676 5984
rect 45716 5944 45717 5984
rect 45675 5935 45717 5944
rect 45388 5900 45428 5909
rect 45428 5860 45620 5900
rect 45388 5851 45428 5860
rect 45388 5732 45428 5741
rect 45291 5648 45333 5657
rect 45291 5608 45292 5648
rect 45332 5608 45333 5648
rect 45291 5599 45333 5608
rect 45388 5489 45428 5692
rect 45387 5480 45429 5489
rect 45387 5440 45388 5480
rect 45428 5440 45429 5480
rect 45387 5431 45429 5440
rect 45580 5153 45620 5860
rect 45676 5732 45716 5935
rect 45676 5683 45716 5692
rect 45868 5489 45908 6280
rect 45964 5993 46004 6364
rect 46156 6320 46196 6364
rect 46060 6280 46196 6320
rect 45963 5984 46005 5993
rect 45963 5944 45964 5984
rect 46004 5944 46005 5984
rect 45963 5935 46005 5944
rect 46060 5825 46100 6280
rect 46059 5816 46101 5825
rect 46059 5776 46060 5816
rect 46100 5776 46101 5816
rect 46059 5767 46101 5776
rect 45867 5480 45909 5489
rect 45867 5440 45868 5480
rect 45908 5440 45909 5480
rect 45867 5431 45909 5440
rect 45675 5312 45717 5321
rect 45675 5272 45676 5312
rect 45716 5272 45717 5312
rect 45675 5263 45717 5272
rect 45579 5144 45621 5153
rect 45579 5104 45580 5144
rect 45620 5104 45621 5144
rect 45579 5095 45621 5104
rect 45580 4892 45620 5095
rect 45580 4843 45620 4852
rect 45579 4724 45621 4733
rect 45579 4684 45580 4724
rect 45620 4684 45621 4724
rect 45579 4675 45621 4684
rect 45483 4388 45525 4397
rect 45483 4348 45484 4388
rect 45524 4348 45525 4388
rect 45483 4339 45525 4348
rect 45484 4254 45524 4339
rect 45580 4229 45620 4675
rect 45579 4220 45621 4229
rect 45579 4180 45580 4220
rect 45620 4180 45621 4220
rect 45579 4171 45621 4180
rect 45387 4052 45429 4061
rect 45387 4012 45388 4052
rect 45428 4012 45429 4052
rect 45387 4003 45429 4012
rect 45292 3464 45332 3473
rect 45099 3380 45141 3389
rect 45099 3340 45100 3380
rect 45140 3340 45141 3380
rect 45099 3331 45141 3340
rect 45100 3212 45140 3221
rect 44907 2456 44949 2465
rect 44907 2416 44908 2456
rect 44948 2416 44949 2456
rect 44907 2407 44949 2416
rect 45100 1205 45140 3172
rect 45292 2717 45332 3424
rect 45291 2708 45333 2717
rect 45291 2668 45292 2708
rect 45332 2668 45333 2708
rect 45291 2659 45333 2668
rect 45099 1196 45141 1205
rect 45099 1156 45100 1196
rect 45140 1156 45141 1196
rect 45099 1147 45141 1156
rect 45195 1028 45237 1037
rect 45195 988 45196 1028
rect 45236 988 45237 1028
rect 45195 979 45237 988
rect 44811 944 44853 953
rect 44811 904 44812 944
rect 44852 904 44853 944
rect 44811 895 44853 904
rect 44812 80 44852 895
rect 45003 272 45045 281
rect 45003 232 45004 272
rect 45044 232 45045 272
rect 45003 223 45045 232
rect 45004 80 45044 223
rect 45196 80 45236 979
rect 45388 80 45428 4003
rect 45484 3212 45524 3221
rect 45484 2549 45524 3172
rect 45483 2540 45525 2549
rect 45483 2500 45484 2540
rect 45524 2500 45525 2540
rect 45483 2491 45525 2500
rect 45580 2465 45620 4171
rect 45676 3464 45716 5263
rect 45868 4892 45908 5431
rect 45868 4843 45908 4852
rect 46060 4892 46100 5767
rect 46252 5732 46292 7624
rect 46444 7589 46484 7876
rect 46539 7916 46581 7925
rect 46539 7876 46540 7916
rect 46580 7876 46581 7916
rect 46539 7867 46581 7876
rect 46923 7916 46965 7925
rect 46923 7876 46924 7916
rect 46964 7876 46965 7916
rect 46923 7867 46965 7876
rect 46924 7782 46964 7867
rect 46539 7748 46581 7757
rect 46539 7708 46540 7748
rect 46580 7708 46581 7748
rect 46539 7699 46581 7708
rect 46540 7614 46580 7699
rect 46443 7580 46485 7589
rect 46443 7540 46444 7580
rect 46484 7540 46485 7580
rect 46443 7531 46485 7540
rect 46444 7244 46484 7531
rect 46636 7421 46676 7506
rect 46635 7412 46677 7421
rect 46635 7372 46636 7412
rect 46676 7372 46772 7412
rect 46635 7363 46677 7372
rect 46540 7244 46580 7253
rect 46444 7204 46540 7244
rect 46540 7195 46580 7204
rect 46636 7244 46676 7255
rect 46636 7169 46676 7204
rect 46347 7160 46389 7169
rect 46347 7120 46348 7160
rect 46388 7120 46389 7160
rect 46347 7111 46389 7120
rect 46635 7160 46677 7169
rect 46635 7120 46636 7160
rect 46676 7120 46677 7160
rect 46635 7111 46677 7120
rect 46348 7026 46388 7111
rect 46636 7001 46676 7111
rect 46635 6992 46677 7001
rect 46635 6952 46636 6992
rect 46676 6952 46677 6992
rect 46635 6943 46677 6952
rect 46732 6833 46772 7372
rect 47020 7076 47060 9211
rect 47116 8756 47156 8767
rect 47116 8681 47156 8716
rect 47115 8672 47157 8681
rect 47115 8632 47116 8672
rect 47156 8632 47157 8672
rect 47115 8623 47157 8632
rect 47499 8168 47541 8177
rect 47212 8128 47444 8168
rect 47116 7916 47156 7925
rect 47116 7589 47156 7876
rect 47212 7916 47252 8128
rect 47307 8000 47349 8009
rect 47307 7960 47308 8000
rect 47348 7960 47349 8000
rect 47307 7951 47349 7960
rect 47212 7867 47252 7876
rect 47211 7748 47253 7757
rect 47211 7708 47212 7748
rect 47252 7708 47253 7748
rect 47211 7699 47253 7708
rect 47212 7614 47252 7699
rect 47115 7580 47157 7589
rect 47115 7540 47116 7580
rect 47156 7540 47157 7580
rect 47115 7531 47157 7540
rect 47116 7244 47156 7531
rect 47308 7244 47348 7951
rect 47156 7204 47252 7244
rect 47116 7195 47156 7204
rect 47212 7076 47252 7204
rect 47308 7195 47348 7204
rect 47020 7036 47156 7076
rect 47212 7036 47348 7076
rect 46731 6824 46773 6833
rect 46731 6784 46732 6824
rect 46772 6784 46773 6824
rect 46731 6775 46773 6784
rect 46636 6488 46676 6497
rect 46348 6404 46388 6413
rect 46348 6161 46388 6364
rect 46347 6152 46389 6161
rect 46347 6112 46348 6152
rect 46388 6112 46389 6152
rect 46347 6103 46389 6112
rect 46636 5900 46676 6448
rect 46828 6236 46868 6245
rect 47020 6236 47060 6245
rect 46868 6196 46964 6236
rect 46828 6187 46868 6196
rect 46827 5984 46869 5993
rect 46827 5944 46828 5984
rect 46868 5944 46869 5984
rect 46827 5935 46869 5944
rect 46156 5692 46292 5732
rect 46444 5860 46676 5900
rect 46156 4985 46196 5692
rect 46155 4976 46197 4985
rect 46155 4936 46156 4976
rect 46196 4936 46197 4976
rect 46155 4927 46197 4936
rect 46060 4843 46100 4852
rect 46156 4892 46196 4927
rect 46156 4841 46196 4852
rect 45867 4724 45909 4733
rect 45867 4684 45868 4724
rect 45908 4684 45909 4724
rect 45867 4675 45909 4684
rect 45868 4590 45908 4675
rect 45963 4388 46005 4397
rect 45963 4348 45964 4388
rect 46004 4348 46005 4388
rect 45963 4339 46005 4348
rect 45964 4220 46004 4339
rect 45771 3968 45813 3977
rect 45771 3928 45772 3968
rect 45812 3928 45813 3968
rect 45771 3919 45813 3928
rect 45676 3415 45716 3424
rect 45579 2456 45621 2465
rect 45579 2416 45580 2456
rect 45620 2416 45621 2456
rect 45579 2407 45621 2416
rect 45579 1616 45621 1625
rect 45579 1576 45580 1616
rect 45620 1576 45621 1616
rect 45579 1567 45621 1576
rect 45580 80 45620 1567
rect 45772 80 45812 3919
rect 45868 3212 45908 3221
rect 45964 3212 46004 4180
rect 46444 4145 46484 5860
rect 46636 5732 46676 5741
rect 46636 5237 46676 5692
rect 46635 5228 46677 5237
rect 46635 5188 46636 5228
rect 46676 5188 46677 5228
rect 46635 5179 46677 5188
rect 46636 4985 46676 5016
rect 46828 4985 46868 5935
rect 46635 4976 46677 4985
rect 46635 4936 46636 4976
rect 46676 4936 46677 4976
rect 46635 4927 46677 4936
rect 46827 4976 46869 4985
rect 46827 4936 46828 4976
rect 46868 4936 46869 4976
rect 46827 4934 46869 4936
rect 46827 4927 46828 4934
rect 46540 4892 46580 4901
rect 46540 4817 46580 4852
rect 46636 4892 46676 4927
rect 46868 4927 46869 4934
rect 46828 4885 46868 4894
rect 46539 4808 46581 4817
rect 46539 4768 46540 4808
rect 46580 4768 46581 4808
rect 46539 4759 46581 4768
rect 46443 4136 46485 4145
rect 46443 4096 46444 4136
rect 46484 4096 46485 4136
rect 46443 4087 46485 4096
rect 46059 4052 46101 4061
rect 46059 4012 46060 4052
rect 46100 4012 46101 4052
rect 46059 4003 46101 4012
rect 46060 3380 46100 4003
rect 46155 3800 46197 3809
rect 46155 3760 46156 3800
rect 46196 3760 46197 3800
rect 46155 3751 46197 3760
rect 46060 3331 46100 3340
rect 46060 3212 46100 3221
rect 45964 3172 46060 3212
rect 45868 2717 45908 3172
rect 46060 3163 46100 3172
rect 45867 2708 45909 2717
rect 45867 2668 45868 2708
rect 45908 2668 45909 2708
rect 45867 2659 45909 2668
rect 45963 1280 46005 1289
rect 45963 1240 45964 1280
rect 46004 1240 46005 1280
rect 45963 1231 46005 1240
rect 45964 80 46004 1231
rect 46156 80 46196 3751
rect 46251 3380 46293 3389
rect 46251 3340 46252 3380
rect 46292 3340 46293 3380
rect 46251 3331 46293 3340
rect 46348 3380 46388 3389
rect 46540 3380 46580 4759
rect 46636 4481 46676 4852
rect 46828 4724 46868 4733
rect 46635 4472 46677 4481
rect 46635 4432 46636 4472
rect 46676 4432 46677 4472
rect 46635 4423 46677 4432
rect 46732 3968 46772 3977
rect 46732 3641 46772 3928
rect 46828 3809 46868 4684
rect 46827 3800 46869 3809
rect 46827 3760 46828 3800
rect 46868 3760 46869 3800
rect 46827 3751 46869 3760
rect 46731 3632 46773 3641
rect 46731 3592 46732 3632
rect 46772 3592 46773 3632
rect 46731 3583 46773 3592
rect 46924 3464 46964 6196
rect 47020 5993 47060 6196
rect 47019 5984 47061 5993
rect 47019 5944 47020 5984
rect 47060 5944 47061 5984
rect 47019 5935 47061 5944
rect 47116 5648 47156 7036
rect 47211 6824 47253 6833
rect 47211 6784 47212 6824
rect 47252 6784 47253 6824
rect 47211 6775 47253 6784
rect 47212 6488 47252 6775
rect 47212 6439 47252 6448
rect 47308 6320 47348 7036
rect 47404 6497 47444 8128
rect 47499 8128 47500 8168
rect 47540 8128 47541 8168
rect 47499 8119 47541 8128
rect 47403 6488 47445 6497
rect 47403 6448 47404 6488
rect 47444 6448 47445 6488
rect 47403 6439 47445 6448
rect 47116 5599 47156 5608
rect 47212 6280 47348 6320
rect 47212 5480 47252 6280
rect 47404 6236 47444 6245
rect 47020 5440 47252 5480
rect 47308 5480 47348 5489
rect 47020 4892 47060 5440
rect 47308 5144 47348 5440
rect 47212 5104 47348 5144
rect 47020 4817 47060 4852
rect 47116 4892 47156 4901
rect 47019 4808 47061 4817
rect 47019 4768 47020 4808
rect 47060 4768 47061 4808
rect 47019 4759 47061 4768
rect 47116 4733 47156 4852
rect 47115 4724 47157 4733
rect 47115 4684 47116 4724
rect 47156 4684 47157 4724
rect 47115 4675 47157 4684
rect 47115 4220 47157 4229
rect 47115 4180 47116 4220
rect 47156 4180 47157 4220
rect 47115 4171 47157 4180
rect 47116 4086 47156 4171
rect 46388 3340 46580 3380
rect 46732 3424 46964 3464
rect 46348 3331 46388 3340
rect 46252 3246 46292 3331
rect 46635 3296 46677 3305
rect 46635 3256 46636 3296
rect 46676 3256 46677 3296
rect 46635 3247 46677 3256
rect 46636 3162 46676 3247
rect 46347 3044 46389 3053
rect 46347 3004 46348 3044
rect 46388 3004 46389 3044
rect 46347 2995 46389 3004
rect 46635 3044 46677 3053
rect 46635 3004 46636 3044
rect 46676 3004 46677 3044
rect 46635 2995 46677 3004
rect 46348 80 46388 2995
rect 46539 2876 46581 2885
rect 46539 2836 46540 2876
rect 46580 2836 46581 2876
rect 46539 2827 46581 2836
rect 46540 80 46580 2827
rect 46636 2633 46676 2995
rect 46635 2624 46677 2633
rect 46635 2584 46636 2624
rect 46676 2584 46677 2624
rect 46635 2575 46677 2584
rect 46732 80 46772 3424
rect 46923 2960 46965 2969
rect 46923 2920 46924 2960
rect 46964 2920 46965 2960
rect 46923 2911 46965 2920
rect 46924 80 46964 2911
rect 47115 2792 47157 2801
rect 47115 2752 47116 2792
rect 47156 2752 47157 2792
rect 47115 2743 47157 2752
rect 47116 80 47156 2743
rect 47212 1121 47252 5104
rect 47308 4985 47348 4987
rect 47307 4976 47349 4985
rect 47307 4936 47308 4976
rect 47348 4936 47349 4976
rect 47307 4927 47349 4936
rect 47308 4892 47348 4927
rect 47308 4843 47348 4852
rect 47308 4724 47348 4733
rect 47308 4229 47348 4684
rect 47307 4220 47349 4229
rect 47307 4180 47308 4220
rect 47348 4180 47349 4220
rect 47307 4171 47349 4180
rect 47404 3716 47444 6196
rect 47500 5648 47540 8119
rect 47596 6488 47636 9463
rect 48171 9176 48213 9185
rect 48171 9136 48172 9176
rect 48212 9136 48213 9176
rect 48171 9127 48213 9136
rect 48075 8588 48117 8597
rect 48075 8548 48076 8588
rect 48116 8548 48117 8588
rect 48075 8539 48117 8548
rect 48076 8454 48116 8539
rect 48172 8084 48212 9127
rect 48268 8681 48308 9472
rect 48460 9462 48500 9547
rect 48844 9428 48884 9437
rect 48844 9344 48884 9388
rect 48940 9428 48980 9547
rect 49804 9521 49844 10387
rect 49803 9512 49845 9521
rect 49803 9472 49804 9512
rect 49844 9472 49845 9512
rect 49803 9463 49845 9472
rect 49516 9428 49556 9437
rect 48940 9379 48980 9388
rect 49132 9388 49516 9428
rect 48460 9304 48884 9344
rect 48460 8849 48500 9304
rect 48940 9260 48980 9269
rect 48844 9220 48940 9260
rect 48844 9017 48884 9220
rect 48940 9211 48980 9220
rect 48843 9008 48885 9017
rect 48843 8968 48844 9008
rect 48884 8968 48885 9008
rect 48843 8959 48885 8968
rect 48459 8840 48501 8849
rect 48459 8800 48460 8840
rect 48500 8800 48501 8840
rect 48459 8791 48501 8800
rect 48363 8756 48405 8765
rect 48363 8716 48364 8756
rect 48404 8716 48405 8756
rect 48363 8707 48405 8716
rect 48267 8672 48309 8681
rect 48267 8632 48268 8672
rect 48308 8632 48309 8672
rect 48267 8623 48309 8632
rect 48268 8177 48308 8623
rect 48364 8622 48404 8707
rect 48460 8504 48500 8791
rect 48748 8765 48788 8796
rect 48747 8756 48789 8765
rect 48747 8716 48748 8756
rect 48788 8716 48789 8756
rect 48747 8707 48789 8716
rect 48364 8464 48500 8504
rect 48748 8672 48788 8707
rect 48267 8168 48309 8177
rect 48267 8128 48268 8168
rect 48308 8128 48309 8168
rect 48267 8119 48309 8128
rect 48172 8035 48212 8044
rect 48364 7916 48404 8464
rect 48364 7253 48404 7876
rect 48460 7916 48500 7925
rect 48500 7876 48692 7916
rect 48460 7867 48500 7876
rect 48460 7748 48500 7757
rect 48171 7244 48213 7253
rect 48171 7204 48172 7244
rect 48212 7204 48213 7244
rect 48171 7195 48213 7204
rect 48363 7244 48405 7253
rect 48363 7204 48364 7244
rect 48404 7204 48405 7244
rect 48363 7195 48405 7204
rect 47979 6908 48021 6917
rect 47979 6868 47980 6908
rect 48020 6868 48021 6908
rect 47979 6859 48021 6868
rect 47884 6581 47924 6666
rect 47883 6572 47925 6581
rect 47883 6532 47884 6572
rect 47924 6532 47925 6572
rect 47883 6523 47925 6532
rect 47596 6439 47636 6448
rect 47691 6488 47733 6497
rect 47691 6448 47692 6488
rect 47732 6448 47733 6488
rect 47691 6439 47733 6448
rect 47692 6320 47732 6439
rect 47884 6404 47924 6413
rect 47980 6404 48020 6859
rect 47924 6364 48020 6404
rect 48075 6404 48117 6413
rect 48075 6364 48076 6404
rect 48116 6364 48117 6404
rect 47884 6355 47924 6364
rect 48075 6355 48117 6364
rect 48172 6404 48212 7195
rect 48460 6833 48500 7708
rect 48556 7244 48596 7253
rect 48556 6917 48596 7204
rect 48652 7169 48692 7876
rect 48748 7841 48788 8632
rect 48747 7832 48789 7841
rect 48747 7792 48748 7832
rect 48788 7792 48789 7832
rect 48747 7783 48789 7792
rect 48748 7244 48788 7253
rect 48844 7244 48884 8959
rect 49132 8840 49172 9388
rect 49516 9379 49556 9388
rect 49612 9428 49652 9437
rect 49652 9388 49748 9428
rect 49612 9379 49652 9388
rect 49516 9260 49556 9269
rect 49323 9008 49365 9017
rect 49516 9008 49556 9220
rect 49611 9260 49653 9269
rect 49611 9220 49612 9260
rect 49652 9220 49653 9260
rect 49611 9211 49653 9220
rect 49612 9017 49652 9211
rect 49323 8968 49324 9008
rect 49364 8968 49556 9008
rect 49611 9008 49653 9017
rect 49611 8968 49612 9008
rect 49652 8968 49653 9008
rect 49323 8959 49365 8968
rect 49611 8959 49653 8968
rect 49324 8924 49364 8959
rect 49324 8873 49364 8884
rect 48940 8800 49172 8840
rect 49419 8840 49461 8849
rect 49419 8800 49420 8840
rect 49460 8800 49461 8840
rect 48940 8681 48980 8800
rect 49419 8791 49461 8800
rect 49324 8756 49364 8765
rect 48939 8672 48981 8681
rect 48939 8632 48940 8672
rect 48980 8632 48981 8672
rect 48939 8623 48981 8632
rect 48940 8588 48980 8623
rect 48940 8538 48980 8548
rect 49324 8504 49364 8716
rect 49420 8756 49460 8791
rect 49420 8705 49460 8716
rect 49612 8756 49652 8959
rect 49708 8849 49748 9388
rect 49804 9378 49844 9463
rect 49900 8924 49940 11395
rect 49996 11360 50036 14920
rect 53163 11948 53205 11957
rect 53163 11908 53164 11948
rect 53204 11908 53205 11948
rect 53163 11899 53205 11908
rect 59691 11948 59733 11957
rect 59691 11908 59692 11948
rect 59732 11908 59733 11948
rect 59691 11899 59733 11908
rect 49996 11320 50132 11360
rect 50092 11024 50132 11320
rect 50092 10975 50132 10984
rect 50284 10781 50324 10866
rect 52107 10856 52149 10865
rect 52107 10816 52108 10856
rect 52148 10816 52149 10856
rect 52107 10807 52149 10816
rect 50283 10772 50325 10781
rect 50283 10732 50284 10772
rect 50324 10732 50325 10772
rect 50283 10723 50325 10732
rect 51243 10772 51285 10781
rect 51243 10732 51244 10772
rect 51284 10732 51285 10772
rect 51243 10723 51285 10732
rect 50288 10604 50656 10613
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50288 10555 50656 10564
rect 50283 10436 50325 10445
rect 50283 10396 50284 10436
rect 50324 10396 50325 10436
rect 50283 10387 50325 10396
rect 51147 10436 51189 10445
rect 51147 10396 51148 10436
rect 51188 10396 51189 10436
rect 51147 10387 51189 10396
rect 50284 10268 50324 10387
rect 50284 10219 50324 10228
rect 51148 9596 51188 10387
rect 51148 9547 51188 9556
rect 50288 9092 50656 9101
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50288 9043 50656 9052
rect 49707 8840 49749 8849
rect 49707 8800 49708 8840
rect 49748 8800 49749 8840
rect 49707 8791 49749 8800
rect 49612 8707 49652 8716
rect 49324 8464 49556 8504
rect 49048 8336 49416 8345
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49048 8287 49416 8296
rect 49516 8261 49556 8464
rect 49515 8252 49557 8261
rect 49515 8212 49516 8252
rect 49556 8212 49557 8252
rect 49515 8203 49557 8212
rect 49419 8168 49461 8177
rect 49419 8128 49420 8168
rect 49460 8128 49461 8168
rect 49419 8119 49461 8128
rect 49228 7916 49268 7925
rect 49131 7748 49173 7757
rect 49131 7708 49132 7748
rect 49172 7708 49173 7748
rect 49131 7699 49173 7708
rect 49036 7244 49076 7253
rect 48788 7204 49036 7244
rect 49132 7244 49172 7699
rect 49228 7589 49268 7876
rect 49420 7832 49460 8119
rect 49420 7783 49460 7792
rect 49516 7757 49556 8203
rect 49611 7916 49653 7925
rect 49900 7916 49940 8884
rect 50188 8840 50228 8849
rect 50228 8800 50516 8840
rect 50188 8791 50228 8800
rect 49995 8756 50037 8765
rect 50476 8756 50516 8800
rect 49995 8716 49996 8756
rect 50036 8716 50132 8756
rect 49995 8707 50037 8716
rect 49996 8622 50036 8707
rect 50092 7925 50132 8716
rect 50516 8716 50612 8756
rect 50476 8707 50516 8716
rect 50572 8000 50612 8716
rect 50956 8504 50996 8513
rect 50763 8252 50805 8261
rect 50763 8212 50764 8252
rect 50804 8212 50805 8252
rect 50763 8203 50805 8212
rect 50764 8168 50804 8203
rect 50764 8117 50804 8128
rect 50572 7951 50612 7960
rect 49611 7876 49612 7916
rect 49652 7876 49653 7916
rect 49611 7867 49653 7876
rect 49897 7876 49940 7916
rect 50091 7916 50133 7925
rect 50188 7916 50228 7925
rect 50091 7876 50092 7916
rect 50132 7876 50188 7916
rect 49515 7748 49557 7757
rect 49515 7708 49516 7748
rect 49556 7708 49557 7748
rect 49515 7699 49557 7708
rect 49612 7748 49652 7867
rect 49897 7832 49937 7876
rect 50091 7867 50133 7876
rect 49995 7832 50037 7841
rect 49897 7792 49940 7832
rect 49227 7580 49269 7589
rect 49227 7540 49228 7580
rect 49268 7540 49269 7580
rect 49227 7531 49269 7540
rect 49228 7244 49268 7253
rect 49132 7204 49228 7244
rect 48651 7160 48693 7169
rect 48651 7120 48652 7160
rect 48692 7120 48693 7160
rect 48651 7111 48693 7120
rect 48555 6908 48597 6917
rect 48555 6868 48556 6908
rect 48596 6868 48597 6908
rect 48555 6859 48597 6868
rect 48459 6824 48501 6833
rect 48459 6784 48460 6824
rect 48500 6784 48501 6824
rect 48459 6775 48501 6784
rect 48652 6656 48692 7111
rect 48748 6833 48788 7204
rect 49036 7195 49076 7204
rect 49228 7195 49268 7204
rect 49323 7244 49365 7253
rect 49323 7204 49324 7244
rect 49364 7204 49365 7244
rect 49323 7195 49365 7204
rect 49516 7244 49556 7253
rect 49612 7244 49652 7708
rect 49804 7706 49844 7715
rect 49900 7706 49940 7792
rect 49995 7792 49996 7832
rect 50036 7792 50037 7832
rect 49995 7783 50037 7792
rect 49844 7666 49940 7706
rect 49996 7698 50036 7783
rect 50092 7782 50132 7867
rect 49804 7657 49844 7666
rect 49900 7589 49940 7666
rect 49899 7580 49941 7589
rect 49899 7540 49900 7580
rect 49940 7540 49941 7580
rect 49899 7531 49941 7540
rect 49556 7204 49652 7244
rect 49708 7245 49748 7253
rect 49900 7245 49940 7531
rect 50092 7245 50132 7253
rect 49708 7244 50132 7245
rect 49748 7205 50092 7244
rect 49516 7195 49556 7204
rect 49708 7195 49748 7204
rect 50188 7244 50228 7876
rect 50288 7580 50656 7589
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50288 7531 50656 7540
rect 50956 7505 50996 8464
rect 51147 8252 51189 8261
rect 51147 8212 51148 8252
rect 51188 8212 51189 8252
rect 51147 8203 51189 8212
rect 50763 7496 50805 7505
rect 50763 7456 50764 7496
rect 50804 7456 50805 7496
rect 50763 7447 50805 7456
rect 50955 7496 50997 7505
rect 50955 7456 50956 7496
rect 50996 7456 51092 7496
rect 50955 7447 50997 7456
rect 50571 7412 50613 7421
rect 50571 7372 50572 7412
rect 50612 7372 50613 7412
rect 50571 7363 50613 7372
rect 50380 7244 50420 7253
rect 50572 7244 50612 7363
rect 50764 7253 50804 7447
rect 50188 7204 50380 7244
rect 50092 7195 50132 7204
rect 50380 7195 50420 7204
rect 50476 7204 50572 7244
rect 49036 7001 49076 7086
rect 49324 7001 49364 7195
rect 49035 6992 49077 7001
rect 49035 6952 49036 6992
rect 49076 6952 49077 6992
rect 49035 6943 49077 6952
rect 49323 6992 49365 7001
rect 49323 6952 49324 6992
rect 49364 6952 49365 6992
rect 49323 6943 49365 6952
rect 49516 6992 49556 7001
rect 48747 6824 48789 6833
rect 48747 6784 48748 6824
rect 48788 6784 48789 6824
rect 48747 6775 48789 6784
rect 49048 6824 49416 6833
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49048 6775 49416 6784
rect 48652 6607 48692 6616
rect 49036 6572 49076 6581
rect 48172 6355 48212 6364
rect 48940 6532 49036 6572
rect 47500 5599 47540 5608
rect 47596 6280 47732 6320
rect 47500 4892 47540 4903
rect 47500 4817 47540 4852
rect 47596 4892 47636 6280
rect 48076 6270 48116 6355
rect 47884 6236 47924 6245
rect 47884 5993 47924 6196
rect 47883 5984 47925 5993
rect 47883 5944 47884 5984
rect 47924 5944 47925 5984
rect 47883 5935 47925 5944
rect 48267 5900 48309 5909
rect 48267 5860 48268 5900
rect 48308 5860 48309 5900
rect 48267 5851 48309 5860
rect 47883 5648 47925 5657
rect 47883 5608 47884 5648
rect 47924 5608 47925 5648
rect 47883 5599 47925 5608
rect 48268 5648 48308 5851
rect 48651 5732 48693 5741
rect 48651 5692 48652 5732
rect 48692 5692 48693 5732
rect 48651 5683 48693 5692
rect 48268 5599 48308 5608
rect 47884 5514 47924 5599
rect 48652 5598 48692 5683
rect 47596 4843 47636 4852
rect 47692 5480 47732 5489
rect 47499 4808 47541 4817
rect 47499 4768 47500 4808
rect 47540 4768 47541 4808
rect 47499 4759 47541 4768
rect 47595 4304 47637 4313
rect 47595 4264 47596 4304
rect 47636 4264 47637 4304
rect 47595 4255 47637 4264
rect 47596 4170 47636 4255
rect 47499 3800 47541 3809
rect 47499 3760 47500 3800
rect 47540 3760 47541 3800
rect 47499 3751 47541 3760
rect 47308 3676 47444 3716
rect 47211 1112 47253 1121
rect 47211 1072 47212 1112
rect 47252 1072 47253 1112
rect 47211 1063 47253 1072
rect 47308 80 47348 3676
rect 47500 3380 47540 3751
rect 47403 3044 47445 3053
rect 47403 3004 47404 3044
rect 47444 3004 47445 3044
rect 47403 2995 47445 3004
rect 47404 2540 47444 2995
rect 47500 2969 47540 3340
rect 47499 2960 47541 2969
rect 47499 2920 47500 2960
rect 47540 2920 47541 2960
rect 47499 2911 47541 2920
rect 47404 2500 47540 2540
rect 47500 80 47540 2500
rect 47692 1289 47732 5440
rect 48076 5480 48116 5489
rect 48460 5480 48500 5489
rect 48116 5440 48308 5480
rect 48076 5431 48116 5440
rect 47788 4985 47828 4987
rect 47787 4976 47829 4985
rect 47787 4936 47788 4976
rect 47828 4936 47829 4976
rect 47787 4927 47829 4936
rect 47980 4976 48020 4985
rect 47788 4892 47828 4927
rect 47788 4843 47828 4852
rect 47787 4724 47829 4733
rect 47787 4684 47788 4724
rect 47828 4684 47829 4724
rect 47787 4675 47829 4684
rect 47788 4590 47828 4675
rect 47980 4565 48020 4936
rect 48172 4724 48212 4733
rect 47979 4556 48021 4565
rect 47979 4516 47980 4556
rect 48020 4516 48021 4556
rect 47979 4507 48021 4516
rect 48172 3557 48212 4684
rect 48268 3716 48308 5440
rect 48500 5440 48884 5480
rect 48460 5431 48500 5440
rect 48363 4976 48405 4985
rect 48363 4936 48364 4976
rect 48404 4936 48405 4976
rect 48363 4927 48405 4936
rect 48747 4976 48789 4985
rect 48747 4936 48748 4976
rect 48788 4936 48789 4976
rect 48747 4927 48789 4936
rect 48364 4842 48404 4927
rect 48748 4842 48788 4927
rect 48459 4724 48501 4733
rect 48459 4684 48460 4724
rect 48500 4684 48501 4724
rect 48459 4675 48501 4684
rect 48556 4724 48596 4733
rect 48596 4684 48692 4724
rect 48556 4675 48596 4684
rect 48460 4220 48500 4675
rect 48500 4180 48596 4220
rect 48460 4171 48500 4180
rect 48556 3725 48596 4180
rect 48555 3716 48597 3725
rect 48268 3676 48500 3716
rect 48171 3548 48213 3557
rect 48171 3508 48172 3548
rect 48212 3508 48213 3548
rect 48171 3499 48213 3508
rect 47979 3464 48021 3473
rect 47979 3424 47980 3464
rect 48020 3424 48021 3464
rect 47979 3415 48021 3424
rect 48364 3464 48404 3473
rect 47980 3330 48020 3415
rect 48172 3212 48212 3221
rect 48172 1625 48212 3172
rect 48364 2801 48404 3424
rect 48363 2792 48405 2801
rect 48363 2752 48364 2792
rect 48404 2752 48405 2792
rect 48363 2743 48405 2752
rect 48267 2624 48309 2633
rect 48267 2584 48268 2624
rect 48308 2584 48309 2624
rect 48267 2575 48309 2584
rect 48171 1616 48213 1625
rect 48171 1576 48172 1616
rect 48212 1576 48213 1616
rect 48171 1567 48213 1576
rect 47691 1280 47733 1289
rect 47691 1240 47692 1280
rect 47732 1240 47733 1280
rect 47691 1231 47733 1240
rect 48075 1280 48117 1289
rect 48075 1240 48076 1280
rect 48116 1240 48117 1280
rect 48075 1231 48117 1240
rect 47883 1196 47925 1205
rect 47883 1156 47884 1196
rect 47924 1156 47925 1196
rect 47883 1147 47925 1156
rect 47691 1112 47733 1121
rect 47691 1072 47692 1112
rect 47732 1072 47733 1112
rect 47691 1063 47733 1072
rect 47692 80 47732 1063
rect 47884 80 47924 1147
rect 48076 80 48116 1231
rect 48268 80 48308 2575
rect 48460 80 48500 3676
rect 48555 3676 48556 3716
rect 48596 3676 48597 3716
rect 48555 3667 48597 3676
rect 48556 3212 48596 3221
rect 48556 1541 48596 3172
rect 48652 3053 48692 4684
rect 48748 3464 48788 3473
rect 48748 3137 48788 3424
rect 48747 3128 48789 3137
rect 48747 3088 48748 3128
rect 48788 3088 48789 3128
rect 48747 3079 48789 3088
rect 48651 3044 48693 3053
rect 48651 3004 48652 3044
rect 48692 3004 48693 3044
rect 48651 2995 48693 3004
rect 48747 2708 48789 2717
rect 48747 2668 48748 2708
rect 48788 2668 48789 2708
rect 48747 2659 48789 2668
rect 48748 1616 48788 2659
rect 48652 1576 48788 1616
rect 48555 1532 48597 1541
rect 48555 1492 48556 1532
rect 48596 1492 48597 1532
rect 48555 1483 48597 1492
rect 48652 80 48692 1576
rect 48844 80 48884 5440
rect 48940 4985 48980 6532
rect 49036 6523 49076 6532
rect 49323 6404 49365 6413
rect 49516 6404 49556 6952
rect 49323 6364 49324 6404
rect 49364 6364 49556 6404
rect 50379 6404 50421 6413
rect 50379 6364 50380 6404
rect 50420 6364 50421 6404
rect 49323 6355 49365 6364
rect 50379 6355 50421 6364
rect 49324 6270 49364 6355
rect 50187 6320 50229 6329
rect 50187 6280 50188 6320
rect 50228 6280 50229 6320
rect 50187 6271 50229 6280
rect 49611 5732 49653 5741
rect 49611 5692 49612 5732
rect 49652 5692 49653 5732
rect 49611 5683 49653 5692
rect 49612 5598 49652 5683
rect 50092 5648 50132 5657
rect 50188 5648 50228 6271
rect 50380 6270 50420 6355
rect 50476 6236 50516 7204
rect 50572 7195 50612 7204
rect 50763 7244 50805 7253
rect 50763 7204 50764 7244
rect 50804 7204 50805 7244
rect 50763 7195 50805 7204
rect 50956 7244 50996 7253
rect 50667 6740 50709 6749
rect 50667 6700 50668 6740
rect 50708 6700 50709 6740
rect 50667 6691 50709 6700
rect 50668 6404 50708 6691
rect 50764 6413 50804 7195
rect 50859 6488 50901 6497
rect 50859 6448 50860 6488
rect 50900 6448 50901 6488
rect 50859 6439 50901 6448
rect 50668 6355 50708 6364
rect 50763 6404 50805 6413
rect 50763 6364 50764 6404
rect 50804 6364 50805 6404
rect 50763 6355 50805 6364
rect 50860 6404 50900 6439
rect 50860 6353 50900 6364
rect 50476 6187 50516 6196
rect 50288 6068 50656 6077
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50288 6019 50656 6028
rect 50956 5825 50996 7204
rect 51052 6329 51092 7456
rect 51148 6404 51188 8203
rect 51244 7916 51284 10723
rect 52108 10268 52148 10807
rect 52491 10520 52533 10529
rect 52491 10480 52492 10520
rect 52532 10480 52533 10520
rect 52491 10471 52533 10480
rect 53067 10520 53109 10529
rect 53067 10480 53068 10520
rect 53108 10480 53109 10520
rect 53067 10471 53109 10480
rect 52108 10219 52148 10228
rect 52107 9596 52149 9605
rect 52107 9556 52108 9596
rect 52148 9556 52149 9596
rect 52107 9547 52149 9556
rect 52299 9596 52341 9605
rect 52299 9556 52300 9596
rect 52340 9556 52341 9596
rect 52299 9547 52341 9556
rect 51436 9437 51476 9522
rect 52012 9437 52052 9522
rect 51340 9428 51380 9437
rect 51340 8261 51380 9388
rect 51435 9428 51477 9437
rect 51435 9388 51436 9428
rect 51476 9388 51477 9428
rect 51435 9379 51477 9388
rect 51819 9428 51861 9437
rect 51819 9388 51820 9428
rect 51860 9388 51861 9428
rect 51819 9379 51861 9388
rect 52011 9428 52053 9437
rect 52011 9388 52012 9428
rect 52052 9388 52053 9428
rect 52011 9379 52053 9388
rect 52108 9428 52148 9547
rect 52300 9462 52340 9547
rect 51435 9260 51477 9269
rect 51435 9220 51436 9260
rect 51476 9220 51477 9260
rect 51435 9211 51477 9220
rect 51436 9126 51476 9211
rect 51339 8252 51381 8261
rect 51339 8212 51340 8252
rect 51380 8212 51381 8252
rect 51339 8203 51381 8212
rect 51436 8084 51476 8093
rect 51476 8044 51668 8084
rect 51436 8035 51476 8044
rect 51339 8000 51381 8009
rect 51339 7960 51340 8000
rect 51380 7960 51381 8000
rect 51339 7951 51381 7960
rect 51244 7421 51284 7876
rect 51243 7412 51285 7421
rect 51243 7372 51244 7412
rect 51284 7372 51285 7412
rect 51243 7363 51285 7372
rect 51340 7412 51380 7951
rect 51340 7363 51380 7372
rect 51436 7916 51476 7925
rect 51436 7253 51476 7876
rect 51628 7916 51668 8044
rect 51820 7916 51860 9379
rect 52011 9260 52053 9269
rect 52011 9220 52012 9260
rect 52052 9220 52053 9260
rect 52011 9211 52053 9220
rect 51668 7876 51764 7916
rect 51628 7867 51668 7876
rect 51724 7664 51764 7876
rect 51860 7876 51956 7916
rect 51820 7867 51860 7876
rect 51724 7624 51860 7664
rect 51531 7412 51573 7421
rect 51531 7372 51532 7412
rect 51572 7372 51573 7412
rect 51531 7363 51573 7372
rect 51243 7244 51285 7253
rect 51243 7204 51244 7244
rect 51284 7204 51285 7244
rect 51243 7195 51285 7204
rect 51435 7244 51477 7253
rect 51435 7204 51436 7244
rect 51476 7204 51477 7244
rect 51435 7195 51477 7204
rect 51532 7244 51572 7363
rect 51244 7110 51284 7195
rect 51435 6824 51477 6833
rect 51435 6784 51436 6824
rect 51476 6784 51477 6824
rect 51435 6775 51477 6784
rect 51436 6656 51476 6775
rect 51436 6607 51476 6616
rect 51243 6572 51285 6581
rect 51243 6532 51244 6572
rect 51284 6532 51285 6572
rect 51243 6523 51285 6532
rect 51148 6355 51188 6364
rect 51244 6404 51284 6523
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51244 6355 51284 6364
rect 51436 6404 51476 6439
rect 51532 6413 51572 7204
rect 51627 7244 51669 7253
rect 51627 7204 51628 7244
rect 51668 7204 51669 7244
rect 51627 7195 51669 7204
rect 51724 7244 51764 7255
rect 51436 6353 51476 6364
rect 51531 6404 51573 6413
rect 51531 6364 51532 6404
rect 51572 6364 51573 6404
rect 51531 6355 51573 6364
rect 51628 6404 51668 7195
rect 51724 7169 51764 7204
rect 51820 7244 51860 7624
rect 51916 7421 51956 7876
rect 51915 7412 51957 7421
rect 51915 7372 51916 7412
rect 51956 7372 51957 7412
rect 51915 7363 51957 7372
rect 51820 7195 51860 7204
rect 51915 7244 51957 7253
rect 51915 7204 51916 7244
rect 51956 7204 51957 7244
rect 51915 7195 51957 7204
rect 52012 7244 52052 9211
rect 51723 7160 51765 7169
rect 51723 7120 51724 7160
rect 51764 7120 51765 7160
rect 51723 7111 51765 7120
rect 51819 7076 51861 7085
rect 51819 7036 51820 7076
rect 51860 7036 51861 7076
rect 51819 7027 51861 7036
rect 51820 6942 51860 7027
rect 51916 6656 51956 7195
rect 51916 6607 51956 6616
rect 52012 6497 52052 7204
rect 52108 7169 52148 9388
rect 52492 9428 52532 10471
rect 53068 10268 53108 10471
rect 53068 9605 53108 10228
rect 53067 9596 53109 9605
rect 53067 9556 53068 9596
rect 53108 9556 53109 9596
rect 53067 9547 53109 9556
rect 52492 9379 52532 9388
rect 52395 9344 52437 9353
rect 52395 9304 52396 9344
rect 52436 9304 52437 9344
rect 52395 9295 52437 9304
rect 52396 8840 52436 9295
rect 52587 9260 52629 9269
rect 52587 9220 52588 9260
rect 52628 9220 52629 9260
rect 52587 9211 52629 9220
rect 52588 8924 52628 9211
rect 52588 8875 52628 8884
rect 52396 8800 52532 8840
rect 52492 8756 52532 8800
rect 52588 8756 52628 8765
rect 52492 8716 52588 8756
rect 52588 8707 52628 8716
rect 52684 8756 52724 8767
rect 52684 8681 52724 8716
rect 52875 8756 52917 8765
rect 52875 8716 52876 8756
rect 52916 8716 52917 8756
rect 52875 8707 52917 8716
rect 52395 8672 52437 8681
rect 52395 8632 52396 8672
rect 52436 8632 52437 8672
rect 52395 8623 52437 8632
rect 52683 8672 52725 8681
rect 52683 8632 52684 8672
rect 52724 8632 52725 8672
rect 52683 8623 52725 8632
rect 52203 7412 52245 7421
rect 52203 7372 52204 7412
rect 52244 7372 52245 7412
rect 52203 7363 52245 7372
rect 52107 7160 52149 7169
rect 52107 7120 52108 7160
rect 52148 7120 52149 7160
rect 52107 7111 52149 7120
rect 52107 6992 52149 7001
rect 52107 6952 52108 6992
rect 52148 6952 52149 6992
rect 52204 6992 52244 7363
rect 52299 7244 52341 7253
rect 52299 7204 52300 7244
rect 52340 7204 52341 7244
rect 52299 7195 52341 7204
rect 52300 7110 52340 7195
rect 52204 6952 52340 6992
rect 52107 6943 52149 6952
rect 52108 6656 52148 6943
rect 52108 6607 52148 6616
rect 52300 6581 52340 6952
rect 52299 6572 52341 6581
rect 52299 6532 52300 6572
rect 52340 6532 52341 6572
rect 52299 6523 52341 6532
rect 52011 6488 52053 6497
rect 52011 6448 52012 6488
rect 52052 6448 52053 6488
rect 52011 6439 52053 6448
rect 51628 6355 51668 6364
rect 51915 6404 51957 6413
rect 51915 6364 51916 6404
rect 51956 6364 51957 6404
rect 51915 6355 51957 6364
rect 51051 6320 51093 6329
rect 51051 6280 51052 6320
rect 51092 6280 51093 6320
rect 51051 6271 51093 6280
rect 51916 6270 51956 6355
rect 52012 6320 52052 6439
rect 52300 6404 52340 6523
rect 52108 6390 52148 6399
rect 52300 6355 52340 6364
rect 52396 6404 52436 8623
rect 52876 8622 52916 8707
rect 52683 8252 52725 8261
rect 52683 8212 52684 8252
rect 52724 8212 52725 8252
rect 52683 8203 52725 8212
rect 52588 6992 52628 7003
rect 52588 6917 52628 6952
rect 52587 6908 52629 6917
rect 52587 6868 52588 6908
rect 52628 6868 52629 6908
rect 52587 6859 52629 6868
rect 52588 6656 52628 6665
rect 52684 6656 52724 8203
rect 52875 7580 52917 7589
rect 52875 7540 52876 7580
rect 52916 7540 52917 7580
rect 52875 7531 52917 7540
rect 52779 7160 52821 7169
rect 52779 7120 52780 7160
rect 52820 7120 52821 7160
rect 52779 7111 52821 7120
rect 52628 6616 52724 6656
rect 52588 6607 52628 6616
rect 52587 6488 52629 6497
rect 52587 6448 52588 6488
rect 52628 6448 52629 6488
rect 52587 6439 52629 6448
rect 52108 6320 52148 6350
rect 52012 6280 52148 6320
rect 51436 6236 51476 6245
rect 50955 5816 50997 5825
rect 50955 5776 50956 5816
rect 50996 5776 50997 5816
rect 50955 5767 50997 5776
rect 51436 5741 51476 6196
rect 51531 6236 51573 6245
rect 51531 6196 51532 6236
rect 51572 6196 51573 6236
rect 51531 6187 51573 6196
rect 51435 5732 51477 5741
rect 51435 5692 51436 5732
rect 51476 5692 51477 5732
rect 51435 5683 51477 5692
rect 50132 5608 50228 5648
rect 50092 5599 50132 5608
rect 49900 5480 49940 5489
rect 49048 5312 49416 5321
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49048 5263 49416 5272
rect 49035 5060 49077 5069
rect 49035 5020 49036 5060
rect 49076 5020 49172 5060
rect 49035 5011 49077 5020
rect 48939 4976 48981 4985
rect 48939 4936 48940 4976
rect 48980 4936 48981 4976
rect 48939 4927 48981 4936
rect 49132 4976 49172 5020
rect 49132 4927 49172 4936
rect 49516 4901 49556 4986
rect 49900 4901 49940 5440
rect 50475 4976 50517 4985
rect 50955 4976 50997 4985
rect 50475 4936 50476 4976
rect 50516 4936 50517 4976
rect 50475 4927 50517 4936
rect 50865 4936 50956 4976
rect 50996 4936 50997 4976
rect 49515 4892 49557 4901
rect 49515 4852 49516 4892
rect 49556 4852 49557 4892
rect 49515 4843 49557 4852
rect 49707 4892 49749 4901
rect 49707 4852 49708 4892
rect 49748 4852 49749 4892
rect 49707 4843 49749 4852
rect 49899 4892 49941 4901
rect 49899 4852 49900 4892
rect 49940 4852 49941 4892
rect 49899 4843 49941 4852
rect 50092 4892 50132 4901
rect 49612 4808 49652 4819
rect 49612 4733 49652 4768
rect 49708 4758 49748 4843
rect 49900 4758 49940 4843
rect 49995 4808 50037 4817
rect 49995 4768 49996 4808
rect 50036 4768 50037 4808
rect 49995 4759 50037 4768
rect 48940 4724 48980 4733
rect 48940 3641 48980 4684
rect 49227 4724 49269 4733
rect 49227 4684 49228 4724
rect 49268 4684 49269 4724
rect 49227 4675 49269 4684
rect 49324 4724 49364 4733
rect 49611 4724 49653 4733
rect 49364 4684 49556 4724
rect 49324 4675 49364 4684
rect 49035 4304 49077 4313
rect 49035 4264 49036 4304
rect 49076 4264 49077 4304
rect 49035 4255 49077 4264
rect 49036 4220 49076 4255
rect 49036 4169 49076 4180
rect 49228 4220 49268 4675
rect 49516 4472 49556 4684
rect 49611 4684 49612 4724
rect 49652 4684 49653 4724
rect 49611 4675 49653 4684
rect 49803 4724 49845 4733
rect 49803 4684 49804 4724
rect 49844 4684 49845 4724
rect 49803 4675 49845 4684
rect 49516 4432 49652 4472
rect 49516 4229 49556 4312
rect 49515 4220 49557 4229
rect 49268 4180 49364 4220
rect 49228 4171 49268 4180
rect 49228 3977 49268 4062
rect 49324 4052 49364 4180
rect 49515 4177 49516 4220
rect 49556 4177 49557 4220
rect 49515 4171 49557 4177
rect 49516 4168 49556 4171
rect 49516 4052 49556 4061
rect 49324 4012 49516 4052
rect 49516 4003 49556 4012
rect 49227 3968 49269 3977
rect 49227 3928 49228 3968
rect 49268 3928 49269 3968
rect 49227 3919 49269 3928
rect 49048 3800 49416 3809
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49048 3751 49416 3760
rect 49515 3800 49557 3809
rect 49515 3760 49516 3800
rect 49556 3760 49557 3800
rect 49515 3751 49557 3760
rect 48939 3632 48981 3641
rect 48939 3592 48940 3632
rect 48980 3592 48981 3632
rect 48939 3583 48981 3592
rect 49419 3632 49461 3641
rect 49419 3592 49420 3632
rect 49460 3592 49461 3632
rect 49419 3583 49461 3592
rect 49035 3548 49077 3557
rect 49035 3508 49036 3548
rect 49076 3508 49077 3548
rect 49035 3499 49077 3508
rect 48939 3212 48981 3221
rect 48939 3172 48940 3212
rect 48980 3172 48981 3212
rect 48939 3163 48981 3172
rect 48940 3078 48980 3163
rect 49036 80 49076 3499
rect 49131 3464 49173 3473
rect 49131 3424 49132 3464
rect 49172 3424 49173 3464
rect 49131 3415 49173 3424
rect 49132 3380 49172 3415
rect 49132 3329 49172 3340
rect 49228 3305 49268 3390
rect 49323 3380 49365 3389
rect 49323 3340 49324 3380
rect 49364 3340 49365 3380
rect 49323 3331 49365 3340
rect 49227 3296 49269 3305
rect 49227 3256 49228 3296
rect 49268 3256 49269 3296
rect 49227 3247 49269 3256
rect 49324 3246 49364 3331
rect 49227 3044 49269 3053
rect 49227 3004 49228 3044
rect 49268 3004 49269 3044
rect 49227 2995 49269 3004
rect 49228 80 49268 2995
rect 49420 80 49460 3583
rect 49516 3548 49556 3751
rect 49612 3716 49652 4432
rect 49804 4052 49844 4675
rect 49996 4472 50036 4759
rect 50092 4556 50132 4852
rect 50284 4892 50324 4901
rect 50187 4724 50229 4733
rect 50284 4724 50324 4852
rect 50476 4892 50516 4927
rect 50865 4905 50905 4936
rect 50955 4927 50997 4936
rect 50476 4841 50516 4852
rect 50668 4892 50708 4901
rect 50865 4856 50905 4865
rect 50380 4733 50420 4818
rect 50571 4808 50613 4817
rect 50668 4808 50708 4852
rect 50571 4768 50572 4808
rect 50612 4768 50708 4808
rect 50571 4759 50613 4768
rect 50187 4684 50188 4724
rect 50228 4684 50324 4724
rect 50379 4724 50421 4733
rect 50379 4684 50380 4724
rect 50420 4684 50421 4724
rect 50187 4675 50229 4684
rect 50379 4675 50421 4684
rect 50764 4724 50804 4733
rect 50187 4556 50229 4565
rect 50092 4516 50188 4556
rect 50228 4516 50229 4556
rect 50187 4507 50229 4516
rect 50288 4556 50656 4565
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50288 4507 50656 4516
rect 49996 4432 50132 4472
rect 49996 4229 50036 4314
rect 49995 4220 50037 4229
rect 49995 4180 49996 4220
rect 50036 4180 50037 4220
rect 49995 4171 50037 4180
rect 49996 4052 50036 4061
rect 49804 4012 49996 4052
rect 49996 4003 50036 4012
rect 49707 3968 49749 3977
rect 49707 3928 49708 3968
rect 49748 3928 49749 3968
rect 49707 3919 49749 3928
rect 49708 3834 49748 3919
rect 49899 3884 49941 3893
rect 49899 3844 49900 3884
rect 49940 3844 49941 3884
rect 49899 3835 49941 3844
rect 49612 3676 49748 3716
rect 49612 3548 49652 3557
rect 49516 3508 49612 3548
rect 49516 3389 49556 3508
rect 49612 3499 49652 3508
rect 49515 3380 49557 3389
rect 49515 3340 49516 3380
rect 49556 3340 49557 3380
rect 49515 3331 49557 3340
rect 49612 3380 49652 3391
rect 49612 3305 49652 3340
rect 49611 3296 49653 3305
rect 49611 3256 49612 3296
rect 49652 3256 49653 3296
rect 49611 3247 49653 3256
rect 49708 2372 49748 3676
rect 49804 3632 49844 3641
rect 49900 3632 49940 3835
rect 50092 3809 50132 4432
rect 50283 4136 50325 4145
rect 50283 4096 50284 4136
rect 50324 4096 50325 4136
rect 50283 4087 50325 4096
rect 50187 4052 50229 4061
rect 50187 4012 50188 4052
rect 50228 4012 50229 4052
rect 50187 4003 50229 4012
rect 50188 3918 50228 4003
rect 50091 3800 50133 3809
rect 50091 3760 50092 3800
rect 50132 3760 50133 3800
rect 50091 3751 50133 3760
rect 49844 3592 49940 3632
rect 49804 3583 49844 3592
rect 50092 3548 50132 3751
rect 50284 3716 50324 4087
rect 50092 3499 50132 3508
rect 50188 3676 50324 3716
rect 50668 3968 50708 3977
rect 50092 3380 50132 3389
rect 50188 3380 50228 3676
rect 50284 3548 50324 3557
rect 50324 3508 50516 3548
rect 50284 3499 50324 3508
rect 50476 3464 50516 3508
rect 50476 3415 50516 3424
rect 50132 3340 50228 3380
rect 50668 3380 50708 3928
rect 50764 3464 50804 4684
rect 50859 4724 50901 4733
rect 50859 4684 50860 4724
rect 50900 4684 50901 4724
rect 50859 4675 50901 4684
rect 50860 4136 50900 4675
rect 50956 4145 50996 4927
rect 51532 4220 51572 6187
rect 52108 5732 52148 6280
rect 52204 5732 52244 5741
rect 52108 5692 52204 5732
rect 52204 5683 52244 5692
rect 52396 5732 52436 6364
rect 52588 6404 52628 6439
rect 52588 6353 52628 6364
rect 52683 6404 52725 6413
rect 52683 6364 52684 6404
rect 52724 6364 52725 6404
rect 52683 6355 52725 6364
rect 52780 6404 52820 7111
rect 52876 6572 52916 7531
rect 53067 7244 53109 7253
rect 53067 7204 53068 7244
rect 53108 7204 53109 7244
rect 53067 7195 53109 7204
rect 52876 6532 53012 6572
rect 52780 6355 52820 6364
rect 52876 6404 52916 6415
rect 52491 6320 52533 6329
rect 52491 6280 52492 6320
rect 52532 6280 52533 6320
rect 52491 6271 52533 6280
rect 52396 5683 52436 5692
rect 52492 5732 52532 6271
rect 52588 6236 52628 6247
rect 52588 6161 52628 6196
rect 52587 6152 52629 6161
rect 52587 6112 52588 6152
rect 52628 6112 52629 6152
rect 52587 6103 52629 6112
rect 52492 5683 52532 5692
rect 52204 5480 52244 5491
rect 52204 5405 52244 5440
rect 52203 5396 52245 5405
rect 52203 5356 52204 5396
rect 52244 5356 52245 5396
rect 52203 5347 52245 5356
rect 52107 5060 52149 5069
rect 52107 5020 52108 5060
rect 52148 5020 52149 5060
rect 52107 5011 52149 5020
rect 51723 4892 51765 4901
rect 51723 4852 51724 4892
rect 51764 4852 51765 4892
rect 51723 4843 51765 4852
rect 51532 4171 51572 4180
rect 51724 4220 51764 4843
rect 52108 4388 52148 5011
rect 52395 4976 52437 4985
rect 52395 4936 52396 4976
rect 52436 4936 52437 4976
rect 52395 4927 52437 4936
rect 52396 4842 52436 4927
rect 52204 4724 52244 4733
rect 52244 4684 52340 4724
rect 52204 4675 52244 4684
rect 52203 4388 52245 4397
rect 52108 4348 52204 4388
rect 52244 4348 52245 4388
rect 52203 4339 52245 4348
rect 52012 4220 52052 4229
rect 51724 4180 52012 4220
rect 50860 4087 50900 4096
rect 50955 4136 50997 4145
rect 50955 4096 50956 4136
rect 50996 4096 50997 4136
rect 50955 4087 50997 4096
rect 51244 4136 51284 4147
rect 51244 4061 51284 4096
rect 51724 4136 51764 4180
rect 52012 4171 52052 4180
rect 52107 4220 52149 4229
rect 52107 4180 52108 4220
rect 52148 4180 52149 4220
rect 52107 4171 52149 4180
rect 52204 4220 52244 4339
rect 52204 4171 52244 4180
rect 51724 4087 51764 4096
rect 52108 4086 52148 4171
rect 51243 4052 51285 4061
rect 51243 4012 51244 4052
rect 51284 4012 51285 4052
rect 51243 4003 51285 4012
rect 51627 4052 51669 4061
rect 51627 4012 51628 4052
rect 51668 4012 51669 4052
rect 51627 4003 51669 4012
rect 51052 3968 51092 3977
rect 50956 3928 51052 3968
rect 50860 3464 50900 3473
rect 50764 3424 50860 3464
rect 50860 3415 50900 3424
rect 50668 3340 50804 3380
rect 50092 3331 50132 3340
rect 50764 3296 50804 3340
rect 50764 3256 50900 3296
rect 50187 3212 50229 3221
rect 50187 3172 50188 3212
rect 50228 3172 50229 3212
rect 50187 3163 50229 3172
rect 50668 3212 50708 3221
rect 50708 3172 50804 3212
rect 50668 3163 50708 3172
rect 49612 2332 49748 2372
rect 49612 80 49652 2332
rect 49803 1616 49845 1625
rect 49803 1576 49804 1616
rect 49844 1576 49845 1616
rect 49803 1567 49845 1576
rect 49804 80 49844 1567
rect 49995 1532 50037 1541
rect 49995 1492 49996 1532
rect 50036 1492 50037 1532
rect 49995 1483 50037 1492
rect 49996 80 50036 1483
rect 50188 80 50228 3163
rect 50288 3044 50656 3053
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50288 2995 50656 3004
rect 50475 2876 50517 2885
rect 50475 2836 50476 2876
rect 50516 2836 50517 2876
rect 50475 2827 50517 2836
rect 50476 440 50516 2827
rect 50571 2036 50613 2045
rect 50571 1996 50572 2036
rect 50612 1996 50613 2036
rect 50571 1987 50613 1996
rect 50380 400 50516 440
rect 50380 80 50420 400
rect 50572 80 50612 1987
rect 50764 80 50804 3172
rect 50860 2045 50900 3256
rect 50956 2885 50996 3928
rect 51052 3919 51092 3928
rect 51628 3918 51668 4003
rect 52203 3716 52245 3725
rect 52203 3676 52204 3716
rect 52244 3676 52245 3716
rect 52203 3667 52245 3676
rect 51435 3548 51477 3557
rect 51435 3508 51436 3548
rect 51476 3508 51477 3548
rect 51435 3499 51477 3508
rect 51436 3464 51476 3499
rect 51436 3413 51476 3424
rect 51819 3464 51861 3473
rect 51819 3424 51820 3464
rect 51860 3424 51861 3464
rect 51819 3415 51861 3424
rect 52204 3464 52244 3667
rect 52204 3415 52244 3424
rect 51820 3330 51860 3415
rect 51052 3212 51092 3221
rect 50955 2876 50997 2885
rect 50955 2836 50956 2876
rect 50996 2836 50997 2876
rect 50955 2827 50997 2836
rect 51052 2540 51092 3172
rect 51244 3212 51284 3221
rect 51244 2540 51284 3172
rect 51628 3212 51668 3221
rect 51628 2540 51668 3172
rect 50956 2500 51092 2540
rect 51148 2500 51284 2540
rect 51340 2500 51668 2540
rect 52012 3212 52052 3221
rect 50859 2036 50901 2045
rect 50859 1996 50860 2036
rect 50900 1996 50901 2036
rect 50859 1987 50901 1996
rect 50956 80 50996 2500
rect 51148 80 51188 2500
rect 51340 80 51380 2500
rect 51915 1700 51957 1709
rect 51915 1660 51916 1700
rect 51956 1660 51957 1700
rect 51915 1651 51957 1660
rect 51531 1616 51573 1625
rect 51531 1576 51532 1616
rect 51572 1576 51573 1616
rect 51531 1567 51573 1576
rect 51532 80 51572 1567
rect 51723 1280 51765 1289
rect 51723 1240 51724 1280
rect 51764 1240 51765 1280
rect 51723 1231 51765 1240
rect 51724 80 51764 1231
rect 51916 80 51956 1651
rect 52012 1625 52052 3172
rect 52300 2372 52340 4684
rect 52684 4388 52724 6355
rect 52876 6329 52916 6364
rect 52875 6320 52917 6329
rect 52875 6280 52876 6320
rect 52916 6280 52917 6320
rect 52875 6271 52917 6280
rect 52972 6152 53012 6532
rect 53068 6488 53108 7195
rect 53068 6439 53108 6448
rect 52876 6112 53012 6152
rect 52779 5144 52821 5153
rect 52779 5104 52780 5144
rect 52820 5104 52821 5144
rect 52779 5095 52821 5104
rect 52780 4892 52820 5095
rect 52876 4985 52916 6112
rect 53164 5648 53204 11899
rect 57675 10604 57717 10613
rect 57675 10564 57676 10604
rect 57716 10564 57717 10604
rect 57675 10555 57717 10564
rect 57964 10564 58196 10604
rect 57676 10436 57716 10555
rect 57676 10387 57716 10396
rect 56235 10352 56277 10361
rect 56235 10312 56236 10352
rect 56276 10312 56277 10352
rect 56235 10303 56277 10312
rect 57579 10352 57621 10361
rect 57579 10312 57580 10352
rect 57620 10312 57621 10352
rect 57579 10303 57621 10312
rect 53451 10100 53493 10109
rect 53451 10060 53452 10100
rect 53492 10060 53493 10100
rect 53451 10051 53493 10060
rect 53452 9428 53492 10051
rect 56236 9680 56276 10303
rect 57580 10268 57620 10303
rect 57580 10217 57620 10228
rect 57772 10268 57812 10277
rect 57964 10268 58004 10564
rect 58059 10436 58101 10445
rect 58059 10396 58060 10436
rect 58100 10396 58101 10436
rect 58059 10387 58101 10396
rect 57812 10228 58004 10268
rect 57772 10219 57812 10228
rect 57291 10100 57333 10109
rect 57291 10060 57292 10100
rect 57332 10060 57333 10100
rect 58060 10100 58100 10387
rect 58156 10361 58196 10564
rect 58155 10352 58197 10361
rect 58635 10352 58677 10361
rect 58155 10312 58156 10352
rect 58196 10312 58197 10352
rect 58155 10303 58197 10312
rect 58618 10312 58636 10352
rect 58676 10312 58677 10352
rect 58618 10303 58677 10312
rect 58827 10352 58869 10361
rect 58827 10312 58828 10352
rect 58868 10312 58869 10352
rect 58827 10303 58869 10312
rect 58156 10268 58196 10303
rect 58156 10219 58196 10228
rect 58618 10268 58658 10303
rect 58618 10219 58658 10228
rect 58828 10184 58868 10303
rect 58924 10268 58964 10277
rect 59116 10268 59156 10277
rect 58924 10184 58964 10228
rect 58828 10144 58964 10184
rect 59020 10228 59116 10268
rect 58156 10100 58196 10109
rect 58060 10060 58156 10100
rect 57291 10051 57333 10060
rect 58156 10051 58196 10060
rect 58443 10100 58485 10109
rect 58443 10060 58444 10100
rect 58484 10060 58485 10100
rect 58443 10051 58485 10060
rect 58635 10100 58677 10109
rect 58635 10060 58636 10100
rect 58676 10060 58677 10100
rect 58635 10051 58677 10060
rect 56236 9631 56276 9640
rect 56619 9680 56661 9689
rect 56619 9640 56620 9680
rect 56660 9640 56661 9680
rect 56619 9631 56661 9640
rect 55851 9596 55893 9605
rect 55851 9556 55852 9596
rect 55892 9556 55893 9596
rect 55851 9547 55893 9556
rect 55852 9462 55892 9547
rect 56620 9546 56660 9631
rect 53452 8765 53492 9388
rect 54795 9428 54837 9437
rect 54795 9388 54796 9428
rect 54836 9388 54837 9428
rect 54795 9379 54837 9388
rect 54988 9428 55028 9437
rect 54796 9294 54836 9379
rect 54892 9344 54932 9353
rect 54892 8924 54932 9304
rect 54796 8884 54932 8924
rect 53451 8756 53493 8765
rect 53451 8716 53452 8756
rect 53492 8716 53493 8756
rect 53451 8707 53493 8716
rect 54316 8756 54356 8767
rect 54316 8681 54356 8716
rect 54508 8756 54548 8765
rect 54796 8756 54836 8884
rect 54988 8849 55028 9388
rect 55659 9428 55701 9437
rect 55659 9388 55660 9428
rect 55700 9388 55701 9428
rect 55659 9379 55701 9388
rect 55756 9428 55796 9437
rect 55467 9092 55509 9101
rect 55467 9052 55468 9092
rect 55508 9052 55509 9092
rect 55467 9043 55509 9052
rect 55468 8924 55508 9043
rect 55468 8875 55508 8884
rect 54988 8840 55036 8849
rect 54988 8800 54995 8840
rect 55035 8800 55036 8840
rect 54994 8791 55036 8800
rect 54548 8716 54836 8756
rect 54508 8707 54548 8716
rect 54315 8672 54357 8681
rect 54315 8632 54316 8672
rect 54356 8632 54357 8672
rect 54315 8623 54357 8632
rect 54412 8672 54452 8681
rect 53835 8504 53877 8513
rect 53835 8464 53836 8504
rect 53876 8464 53877 8504
rect 53835 8455 53877 8464
rect 53355 6740 53397 6749
rect 53355 6700 53356 6740
rect 53396 6700 53397 6740
rect 53355 6691 53397 6700
rect 53260 6572 53300 6581
rect 53260 6329 53300 6532
rect 53356 6497 53396 6691
rect 53355 6488 53397 6497
rect 53355 6448 53356 6488
rect 53396 6448 53397 6488
rect 53355 6439 53397 6448
rect 53259 6320 53301 6329
rect 53259 6280 53260 6320
rect 53300 6280 53301 6320
rect 53259 6271 53301 6280
rect 53164 5599 53204 5608
rect 53163 5144 53205 5153
rect 53163 5104 53164 5144
rect 53204 5104 53205 5144
rect 53163 5095 53205 5104
rect 52875 4976 52917 4985
rect 52875 4936 52876 4976
rect 52916 4936 52917 4976
rect 52875 4927 52917 4936
rect 52780 4843 52820 4852
rect 52492 4348 52724 4388
rect 53164 4388 53204 5095
rect 53260 4733 53300 6271
rect 53356 5900 53396 6439
rect 53451 6152 53493 6161
rect 53451 6112 53452 6152
rect 53492 6112 53493 6152
rect 53451 6103 53493 6112
rect 53356 5851 53396 5860
rect 53259 4724 53301 4733
rect 53259 4684 53260 4724
rect 53300 4684 53301 4724
rect 53259 4675 53301 4684
rect 53259 4556 53301 4565
rect 53259 4516 53260 4556
rect 53300 4516 53301 4556
rect 53259 4507 53301 4516
rect 52395 4220 52437 4229
rect 52395 4180 52396 4220
rect 52436 4180 52437 4220
rect 52395 4171 52437 4180
rect 52396 4086 52436 4171
rect 52396 3968 52436 3977
rect 52396 3473 52436 3928
rect 52492 3725 52532 4348
rect 53164 4339 53204 4348
rect 52971 4304 53013 4313
rect 52971 4264 52972 4304
rect 53012 4264 53013 4304
rect 52971 4255 53013 4264
rect 52588 4220 52628 4229
rect 52588 4145 52628 4180
rect 52683 4220 52725 4229
rect 52683 4180 52684 4220
rect 52724 4180 52725 4220
rect 52683 4171 52725 4180
rect 52875 4220 52917 4229
rect 52875 4180 52876 4220
rect 52916 4180 52917 4220
rect 52875 4171 52917 4180
rect 52972 4220 53012 4255
rect 52587 4136 52629 4145
rect 52587 4096 52588 4136
rect 52628 4096 52629 4136
rect 52587 4087 52629 4096
rect 52491 3716 52533 3725
rect 52491 3676 52492 3716
rect 52532 3676 52533 3716
rect 52491 3667 52533 3676
rect 52491 3548 52533 3557
rect 52491 3508 52492 3548
rect 52532 3508 52533 3548
rect 52491 3499 52533 3508
rect 52395 3464 52437 3473
rect 52395 3424 52396 3464
rect 52436 3424 52437 3464
rect 52395 3415 52437 3424
rect 52492 3414 52532 3499
rect 52588 3380 52628 4087
rect 52684 3548 52724 4171
rect 52876 4052 52916 4171
rect 52972 4169 53012 4180
rect 52972 4052 53012 4061
rect 52876 4012 52972 4052
rect 52972 4003 53012 4012
rect 52779 3968 52821 3977
rect 52779 3928 52780 3968
rect 52820 3928 52821 3968
rect 52779 3919 52821 3928
rect 52684 3499 52724 3508
rect 52684 3380 52724 3389
rect 52588 3340 52684 3380
rect 52684 3331 52724 3340
rect 52108 2332 52340 2372
rect 52011 1616 52053 1625
rect 52011 1576 52012 1616
rect 52052 1576 52053 1616
rect 52011 1567 52053 1576
rect 52108 80 52148 2332
rect 52780 2036 52820 3919
rect 52875 3800 52917 3809
rect 52875 3760 52876 3800
rect 52916 3760 52917 3800
rect 52875 3751 52917 3760
rect 52684 1996 52820 2036
rect 52491 1784 52533 1793
rect 52491 1744 52492 1784
rect 52532 1744 52533 1784
rect 52491 1735 52533 1744
rect 52299 1616 52341 1625
rect 52299 1576 52300 1616
rect 52340 1576 52341 1616
rect 52299 1567 52341 1576
rect 52300 80 52340 1567
rect 52492 80 52532 1735
rect 52684 80 52724 1996
rect 52876 80 52916 3751
rect 53164 3464 53204 3473
rect 53260 3464 53300 4507
rect 53355 4220 53397 4229
rect 53355 4180 53356 4220
rect 53396 4180 53397 4220
rect 53355 4171 53397 4180
rect 53356 4086 53396 4171
rect 53356 3968 53396 3977
rect 53356 3725 53396 3928
rect 53355 3716 53397 3725
rect 53355 3676 53356 3716
rect 53396 3676 53397 3716
rect 53355 3667 53397 3676
rect 53204 3424 53300 3464
rect 53452 3464 53492 6103
rect 53739 5984 53781 5993
rect 53739 5944 53740 5984
rect 53780 5944 53781 5984
rect 53739 5935 53781 5944
rect 53740 5732 53780 5935
rect 53548 5692 53740 5732
rect 53548 4313 53588 5692
rect 53740 5683 53780 5692
rect 53644 4808 53684 4817
rect 53547 4304 53589 4313
rect 53547 4264 53548 4304
rect 53588 4264 53589 4304
rect 53547 4255 53589 4264
rect 53548 4220 53588 4255
rect 53548 4170 53588 4180
rect 53644 3893 53684 4768
rect 53739 3968 53781 3977
rect 53739 3928 53740 3968
rect 53780 3928 53781 3968
rect 53739 3919 53781 3928
rect 53643 3884 53685 3893
rect 53643 3844 53644 3884
rect 53684 3844 53685 3884
rect 53643 3835 53685 3844
rect 53740 3834 53780 3919
rect 53548 3464 53588 3473
rect 53452 3424 53548 3464
rect 53836 3464 53876 8455
rect 54412 8168 54452 8632
rect 54796 8588 54836 8716
rect 54892 8765 54932 8773
rect 54892 8764 54951 8765
rect 54932 8756 54951 8764
rect 54892 8716 54910 8724
rect 54950 8716 54951 8756
rect 54892 8715 54951 8716
rect 54909 8707 54951 8715
rect 55276 8756 55316 8765
rect 55316 8716 55412 8756
rect 55276 8707 55316 8716
rect 54910 8647 54950 8707
rect 54892 8588 54932 8597
rect 55276 8588 55316 8597
rect 54796 8548 54892 8588
rect 54932 8548 55276 8588
rect 54892 8539 54932 8548
rect 54699 8504 54741 8513
rect 54699 8464 54700 8504
rect 54740 8464 54741 8504
rect 54699 8455 54741 8464
rect 54700 8370 54740 8455
rect 54603 8336 54645 8345
rect 54603 8296 54604 8336
rect 54644 8296 54645 8336
rect 54603 8287 54645 8296
rect 54220 8128 54452 8168
rect 54604 8168 54644 8287
rect 53932 6404 53972 6413
rect 53932 5993 53972 6364
rect 54124 6404 54164 6413
rect 54124 6245 54164 6364
rect 54123 6236 54165 6245
rect 54123 6196 54124 6236
rect 54164 6196 54165 6236
rect 54123 6187 54165 6196
rect 53931 5984 53973 5993
rect 53931 5944 53932 5984
rect 53972 5944 53973 5984
rect 53931 5935 53973 5944
rect 53932 5741 53972 5826
rect 53931 5732 53973 5741
rect 53931 5692 53932 5732
rect 53972 5692 53973 5732
rect 53931 5683 53973 5692
rect 53932 5480 53972 5489
rect 53972 5440 54164 5480
rect 53932 5431 53972 5440
rect 54028 4892 54068 4901
rect 53931 4808 53973 4817
rect 53931 4768 53932 4808
rect 53972 4768 53973 4808
rect 53931 4759 53973 4768
rect 53932 4136 53972 4759
rect 54028 4649 54068 4852
rect 54027 4640 54069 4649
rect 54027 4600 54028 4640
rect 54068 4600 54069 4640
rect 54027 4591 54069 4600
rect 54124 4145 54164 5440
rect 53932 4087 53972 4096
rect 54123 4136 54165 4145
rect 54123 4096 54124 4136
rect 54164 4096 54165 4136
rect 54123 4087 54165 4096
rect 54027 3968 54069 3977
rect 54027 3928 54028 3968
rect 54068 3928 54069 3968
rect 54027 3919 54069 3928
rect 54124 3968 54164 3977
rect 53932 3464 53972 3473
rect 53836 3424 53932 3464
rect 53164 3415 53204 3424
rect 53548 3415 53588 3424
rect 53932 3415 53972 3424
rect 53643 3380 53685 3389
rect 53643 3340 53644 3380
rect 53684 3340 53685 3380
rect 53643 3331 53685 3340
rect 52972 3212 53012 3221
rect 52972 1289 53012 3172
rect 53356 3212 53396 3221
rect 53356 1709 53396 3172
rect 53451 3212 53493 3221
rect 53451 3172 53452 3212
rect 53492 3172 53493 3212
rect 53451 3163 53493 3172
rect 53355 1700 53397 1709
rect 53355 1660 53356 1700
rect 53396 1660 53397 1700
rect 53355 1651 53397 1660
rect 53067 1448 53109 1457
rect 53067 1408 53068 1448
rect 53108 1408 53109 1448
rect 53067 1399 53109 1408
rect 52971 1280 53013 1289
rect 52971 1240 52972 1280
rect 53012 1240 53013 1280
rect 52971 1231 53013 1240
rect 53068 80 53108 1399
rect 53259 1280 53301 1289
rect 53259 1240 53260 1280
rect 53300 1240 53301 1280
rect 53259 1231 53301 1240
rect 53260 80 53300 1231
rect 53452 80 53492 3163
rect 53644 80 53684 3331
rect 53740 3212 53780 3221
rect 53740 1625 53780 3172
rect 53739 1616 53781 1625
rect 53739 1576 53740 1616
rect 53780 1576 53781 1616
rect 53739 1567 53781 1576
rect 53835 1364 53877 1373
rect 53835 1324 53836 1364
rect 53876 1324 53877 1364
rect 53835 1315 53877 1324
rect 53836 80 53876 1315
rect 54028 80 54068 3919
rect 54124 3809 54164 3928
rect 54123 3800 54165 3809
rect 54123 3760 54124 3800
rect 54164 3760 54165 3800
rect 54123 3751 54165 3760
rect 54220 3464 54260 8128
rect 54604 8119 54644 8128
rect 54411 8000 54453 8009
rect 54411 7960 54412 8000
rect 54452 7960 54453 8000
rect 54411 7951 54453 7960
rect 54699 8000 54741 8009
rect 54699 7960 54700 8000
rect 54740 7960 54741 8000
rect 54699 7951 54741 7960
rect 54412 7866 54452 7951
rect 54604 7748 54644 7757
rect 54508 7708 54604 7748
rect 54315 7412 54357 7421
rect 54315 7372 54316 7412
rect 54356 7372 54357 7412
rect 54315 7363 54357 7372
rect 54316 7244 54356 7363
rect 54316 7195 54356 7204
rect 54508 7244 54548 7708
rect 54604 7699 54644 7708
rect 54508 7195 54548 7204
rect 54700 7076 54740 7951
rect 54795 7916 54837 7925
rect 54795 7876 54796 7916
rect 54836 7876 54837 7916
rect 54795 7867 54837 7876
rect 54988 7916 55028 8548
rect 55276 8539 55316 8548
rect 55372 7925 55412 8716
rect 54988 7867 55028 7876
rect 55371 7916 55413 7925
rect 55371 7876 55372 7916
rect 55412 7876 55413 7916
rect 55371 7867 55413 7876
rect 54508 7036 54740 7076
rect 54412 6992 54452 7001
rect 54412 6572 54452 6952
rect 54316 6532 54412 6572
rect 54316 6245 54356 6532
rect 54412 6523 54452 6532
rect 54412 6404 54452 6415
rect 54412 6329 54452 6364
rect 54411 6320 54453 6329
rect 54411 6280 54412 6320
rect 54452 6280 54453 6320
rect 54411 6271 54453 6280
rect 54315 6236 54357 6245
rect 54315 6196 54316 6236
rect 54356 6196 54357 6236
rect 54315 6187 54357 6196
rect 54316 5741 54356 6187
rect 54508 6152 54548 7036
rect 54796 6992 54836 7867
rect 54891 7748 54933 7757
rect 54891 7708 54892 7748
rect 54932 7708 54933 7748
rect 54891 7699 54933 7708
rect 54892 7614 54932 7699
rect 55372 7673 55412 7867
rect 55371 7664 55413 7673
rect 55371 7624 55372 7664
rect 55412 7624 55413 7664
rect 55371 7615 55413 7624
rect 54700 6952 54836 6992
rect 54700 6329 54740 6952
rect 55660 6833 55700 9379
rect 55756 7421 55796 9388
rect 55948 9428 55988 9439
rect 55948 9353 55988 9388
rect 56139 9428 56181 9437
rect 56139 9388 56140 9428
rect 56180 9388 56181 9428
rect 56139 9379 56181 9388
rect 56332 9428 56372 9439
rect 55947 9344 55989 9353
rect 55947 9304 55948 9344
rect 55988 9304 55989 9344
rect 55947 9295 55989 9304
rect 56140 9294 56180 9379
rect 56332 9353 56372 9388
rect 56524 9428 56564 9437
rect 56331 9344 56373 9353
rect 56331 9304 56332 9344
rect 56372 9304 56373 9344
rect 56331 9295 56373 9304
rect 56524 8840 56564 9388
rect 56716 9428 56756 9439
rect 56716 9353 56756 9388
rect 56715 9344 56757 9353
rect 56715 9304 56716 9344
rect 56756 9304 56757 9344
rect 56715 9295 56757 9304
rect 56140 8800 56564 8840
rect 56811 8840 56853 8849
rect 56811 8800 56812 8840
rect 56852 8800 56853 8840
rect 55947 8756 55989 8765
rect 55947 8716 55948 8756
rect 55988 8716 55989 8756
rect 55947 8707 55989 8716
rect 56140 8756 56180 8800
rect 56811 8791 56853 8800
rect 57195 8840 57237 8849
rect 57195 8800 57196 8840
rect 57236 8800 57237 8840
rect 57195 8791 57237 8800
rect 56812 8764 56852 8791
rect 55948 7916 55988 8707
rect 56043 8588 56085 8597
rect 56043 8548 56044 8588
rect 56084 8548 56085 8588
rect 56043 8539 56085 8548
rect 56044 8454 56084 8539
rect 56140 8513 56180 8716
rect 56332 8716 56660 8756
rect 56139 8504 56181 8513
rect 56139 8464 56140 8504
rect 56180 8464 56181 8504
rect 56139 8455 56181 8464
rect 56044 7916 56084 7925
rect 55948 7876 56044 7916
rect 56044 7867 56084 7876
rect 56139 7916 56181 7925
rect 56139 7876 56140 7916
rect 56180 7876 56181 7916
rect 56139 7867 56181 7876
rect 56236 7916 56276 7925
rect 56140 7782 56180 7867
rect 55851 7496 55893 7505
rect 55851 7456 55852 7496
rect 55892 7456 55893 7496
rect 55851 7447 55893 7456
rect 55755 7412 55797 7421
rect 55755 7372 55756 7412
rect 55796 7372 55797 7412
rect 55755 7363 55797 7372
rect 55659 6824 55701 6833
rect 55659 6784 55660 6824
rect 55700 6784 55701 6824
rect 55659 6775 55701 6784
rect 54988 6572 55028 6581
rect 54892 6532 54988 6572
rect 54795 6404 54837 6413
rect 54795 6364 54796 6404
rect 54836 6364 54837 6404
rect 54795 6355 54837 6364
rect 54699 6320 54741 6329
rect 54699 6280 54700 6320
rect 54740 6280 54741 6320
rect 54699 6271 54741 6280
rect 54412 6112 54548 6152
rect 54604 6236 54644 6245
rect 54315 5732 54357 5741
rect 54315 5692 54316 5732
rect 54356 5692 54357 5732
rect 54315 5683 54357 5692
rect 54316 5480 54356 5489
rect 54316 4565 54356 5440
rect 54315 4556 54357 4565
rect 54315 4516 54316 4556
rect 54356 4516 54357 4556
rect 54315 4507 54357 4516
rect 54316 4136 54356 4145
rect 54412 4136 54452 6112
rect 54604 5993 54644 6196
rect 54796 6236 54836 6355
rect 54892 6245 54932 6532
rect 54988 6523 55028 6532
rect 55179 6572 55221 6581
rect 55179 6532 55180 6572
rect 55220 6532 55221 6572
rect 55179 6523 55221 6532
rect 54987 6404 55029 6413
rect 54987 6364 54988 6404
rect 55028 6364 55029 6404
rect 54987 6355 55029 6364
rect 54796 6187 54836 6196
rect 54891 6236 54933 6245
rect 54891 6196 54892 6236
rect 54932 6196 54933 6236
rect 54891 6187 54933 6196
rect 54603 5984 54645 5993
rect 54603 5944 54604 5984
rect 54644 5944 54645 5984
rect 54603 5935 54645 5944
rect 54988 5741 55028 6355
rect 54507 5732 54549 5741
rect 54987 5732 55029 5741
rect 54507 5692 54508 5732
rect 54548 5692 54644 5732
rect 54507 5683 54549 5692
rect 54508 5598 54548 5683
rect 54507 4640 54549 4649
rect 54507 4600 54508 4640
rect 54548 4600 54549 4640
rect 54507 4591 54549 4600
rect 54508 4397 54548 4591
rect 54507 4388 54549 4397
rect 54507 4348 54508 4388
rect 54548 4348 54549 4388
rect 54507 4339 54549 4348
rect 54604 4220 54644 5692
rect 54987 5692 54988 5732
rect 55028 5692 55029 5732
rect 54987 5683 55029 5692
rect 54891 5648 54933 5657
rect 54891 5608 54892 5648
rect 54932 5608 54933 5648
rect 54891 5599 54933 5608
rect 54892 5514 54932 5599
rect 54604 4171 54644 4180
rect 54700 5480 54740 5489
rect 55084 5480 55124 5489
rect 54356 4096 54452 4136
rect 54316 4087 54356 4096
rect 54316 3464 54356 3473
rect 54220 3424 54316 3464
rect 54316 3415 54356 3424
rect 54124 3212 54164 3221
rect 54124 1793 54164 3172
rect 54604 3212 54644 3221
rect 54604 2801 54644 3172
rect 54603 2792 54645 2801
rect 54603 2752 54604 2792
rect 54644 2752 54645 2792
rect 54603 2743 54645 2752
rect 54700 2540 54740 5440
rect 54988 5440 55084 5480
rect 54988 5060 55028 5440
rect 55084 5431 55124 5440
rect 55180 5228 55220 6523
rect 55563 6404 55605 6413
rect 55372 6364 55508 6404
rect 55372 6161 55412 6364
rect 55468 6245 55508 6364
rect 55563 6364 55564 6404
rect 55604 6364 55605 6404
rect 55563 6355 55605 6364
rect 55756 6405 55796 6413
rect 55852 6405 55892 7447
rect 56139 7412 56181 7421
rect 56139 7372 56140 7412
rect 56180 7372 56181 7412
rect 56139 7363 56181 7372
rect 56044 6992 56084 7001
rect 55756 6404 55892 6405
rect 55796 6365 55892 6404
rect 55948 6952 56044 6992
rect 55756 6355 55796 6364
rect 55564 6270 55604 6355
rect 55467 6236 55509 6245
rect 55467 6196 55468 6236
rect 55508 6196 55509 6236
rect 55467 6187 55509 6196
rect 55371 6152 55413 6161
rect 55371 6112 55372 6152
rect 55412 6112 55413 6152
rect 55371 6103 55413 6112
rect 55659 6152 55701 6161
rect 55659 6112 55660 6152
rect 55700 6112 55701 6152
rect 55659 6103 55701 6112
rect 55275 6068 55317 6077
rect 55275 6028 55276 6068
rect 55316 6028 55317 6068
rect 55275 6019 55317 6028
rect 55276 5648 55316 6019
rect 55660 5732 55700 6103
rect 55851 5816 55893 5825
rect 55851 5776 55852 5816
rect 55892 5776 55893 5816
rect 55851 5767 55893 5776
rect 55660 5683 55700 5692
rect 55755 5732 55797 5741
rect 55755 5692 55756 5732
rect 55796 5692 55797 5732
rect 55755 5683 55797 5692
rect 55852 5732 55892 5767
rect 55276 5599 55316 5608
rect 55756 5598 55796 5683
rect 55852 5681 55892 5692
rect 55659 5564 55701 5573
rect 55659 5524 55660 5564
rect 55700 5524 55701 5564
rect 55659 5515 55701 5524
rect 55371 5312 55413 5321
rect 55371 5272 55372 5312
rect 55412 5272 55413 5312
rect 55371 5263 55413 5272
rect 54892 5020 55028 5060
rect 55084 5188 55220 5228
rect 54795 4892 54837 4901
rect 54795 4852 54796 4892
rect 54836 4852 54837 4892
rect 54795 4843 54837 4852
rect 54796 4229 54836 4843
rect 54795 4220 54837 4229
rect 54795 4180 54796 4220
rect 54836 4180 54837 4220
rect 54795 4171 54837 4180
rect 54795 4052 54837 4061
rect 54795 4012 54796 4052
rect 54836 4012 54837 4052
rect 54795 4003 54837 4012
rect 54796 3641 54836 4003
rect 54795 3632 54837 3641
rect 54795 3592 54796 3632
rect 54836 3592 54837 3632
rect 54795 3583 54837 3592
rect 54796 3548 54836 3583
rect 54796 3497 54836 3508
rect 54796 3380 54836 3391
rect 54796 3305 54836 3340
rect 54795 3296 54837 3305
rect 54795 3256 54796 3296
rect 54836 3256 54837 3296
rect 54795 3247 54837 3256
rect 54412 2500 54740 2540
rect 54123 1784 54165 1793
rect 54123 1744 54124 1784
rect 54164 1744 54165 1784
rect 54123 1735 54165 1744
rect 54219 1616 54261 1625
rect 54219 1576 54220 1616
rect 54260 1576 54261 1616
rect 54219 1567 54261 1576
rect 54220 80 54260 1567
rect 54412 80 54452 2500
rect 54603 2372 54645 2381
rect 54603 2332 54604 2372
rect 54644 2332 54645 2372
rect 54603 2323 54645 2332
rect 54604 80 54644 2323
rect 54892 860 54932 5020
rect 54988 4892 55028 4901
rect 54988 4313 55028 4852
rect 55084 4472 55124 5188
rect 55179 4892 55221 4901
rect 55179 4852 55180 4892
rect 55220 4852 55221 4892
rect 55179 4843 55221 4852
rect 55372 4892 55412 5263
rect 55180 4758 55220 4843
rect 55276 4724 55316 4733
rect 55084 4432 55220 4472
rect 55180 4388 55220 4432
rect 55276 4397 55316 4684
rect 55180 4339 55220 4348
rect 55275 4388 55317 4397
rect 55275 4348 55276 4388
rect 55316 4348 55317 4388
rect 55275 4339 55317 4348
rect 54987 4304 55029 4313
rect 54987 4264 54988 4304
rect 55028 4264 55029 4304
rect 54987 4255 55029 4264
rect 55084 4229 55124 4314
rect 55083 4220 55125 4229
rect 55083 4180 55084 4220
rect 55124 4180 55125 4220
rect 55083 4171 55125 4180
rect 55276 4220 55316 4229
rect 55372 4209 55412 4852
rect 55316 4180 55412 4209
rect 55276 4169 55412 4180
rect 54987 4136 55029 4145
rect 54987 4096 54988 4136
rect 55028 4096 55029 4136
rect 54987 4087 55029 4096
rect 54988 3305 55028 4087
rect 55275 3800 55317 3809
rect 55275 3760 55276 3800
rect 55316 3760 55317 3800
rect 55275 3751 55317 3760
rect 55276 3464 55316 3751
rect 55372 3641 55412 4169
rect 55564 4724 55604 4733
rect 55468 3968 55508 3977
rect 55371 3632 55413 3641
rect 55371 3592 55372 3632
rect 55412 3592 55413 3632
rect 55371 3583 55413 3592
rect 55276 3415 55316 3424
rect 55468 3389 55508 3928
rect 55467 3380 55509 3389
rect 55467 3340 55468 3380
rect 55508 3340 55509 3380
rect 55467 3331 55509 3340
rect 54987 3296 55029 3305
rect 54987 3256 54988 3296
rect 55028 3256 55029 3296
rect 54987 3247 55029 3256
rect 55275 3296 55317 3305
rect 55275 3256 55276 3296
rect 55316 3256 55317 3296
rect 55275 3247 55317 3256
rect 55084 3212 55124 3221
rect 54987 1532 55029 1541
rect 54987 1492 54988 1532
rect 55028 1492 55029 1532
rect 54987 1483 55029 1492
rect 54796 820 54932 860
rect 54796 80 54836 820
rect 54988 80 55028 1483
rect 55084 1457 55124 3172
rect 55276 2885 55316 3247
rect 55468 3212 55508 3221
rect 55275 2876 55317 2885
rect 55275 2836 55276 2876
rect 55316 2836 55317 2876
rect 55275 2827 55317 2836
rect 55371 2288 55413 2297
rect 55371 2248 55372 2288
rect 55412 2248 55413 2288
rect 55371 2239 55413 2248
rect 55179 1700 55221 1709
rect 55179 1660 55180 1700
rect 55220 1660 55221 1700
rect 55179 1651 55221 1660
rect 55083 1448 55125 1457
rect 55083 1408 55084 1448
rect 55124 1408 55125 1448
rect 55083 1399 55125 1408
rect 55180 80 55220 1651
rect 55372 80 55412 2239
rect 55468 1289 55508 3172
rect 55564 2540 55604 4684
rect 55660 4304 55700 5515
rect 55948 5144 55988 6952
rect 56044 6943 56084 6952
rect 56140 6908 56180 7363
rect 56236 7337 56276 7876
rect 56235 7328 56277 7337
rect 56235 7288 56236 7328
rect 56276 7288 56277 7328
rect 56235 7279 56277 7288
rect 56235 7160 56277 7169
rect 56235 7120 56236 7160
rect 56276 7120 56277 7160
rect 56235 7111 56277 7120
rect 56236 7026 56276 7111
rect 56140 6868 56276 6908
rect 56043 6824 56085 6833
rect 56043 6784 56044 6824
rect 56084 6784 56085 6824
rect 56043 6775 56085 6784
rect 56044 6404 56084 6775
rect 56044 6355 56084 6364
rect 56236 6404 56276 6868
rect 56236 6355 56276 6364
rect 56139 6320 56181 6329
rect 56139 6280 56140 6320
rect 56180 6280 56181 6320
rect 56139 6271 56181 6280
rect 56140 6186 56180 6271
rect 56332 6245 56372 8716
rect 56427 8588 56469 8597
rect 56427 8548 56428 8588
rect 56468 8548 56469 8588
rect 56427 8539 56469 8548
rect 56620 8588 56660 8716
rect 56812 8705 56852 8724
rect 57196 8764 57236 8791
rect 57196 8705 57236 8724
rect 56620 8539 56660 8548
rect 56715 8588 56757 8597
rect 56812 8588 56852 8597
rect 56715 8548 56716 8588
rect 56756 8548 56812 8588
rect 56715 8539 56757 8548
rect 56812 8539 56852 8548
rect 57003 8588 57045 8597
rect 57003 8548 57004 8588
rect 57044 8548 57045 8588
rect 57003 8539 57045 8548
rect 57195 8588 57237 8597
rect 57195 8548 57196 8588
rect 57236 8548 57237 8588
rect 57195 8539 57237 8548
rect 56428 7916 56468 8539
rect 56619 8084 56661 8093
rect 56619 8044 56620 8084
rect 56660 8044 56661 8084
rect 56619 8035 56661 8044
rect 56428 7867 56468 7876
rect 56620 7916 56660 8035
rect 56620 7867 56660 7876
rect 56812 7916 56852 7925
rect 56524 7748 56564 7757
rect 56524 7589 56564 7708
rect 56812 7673 56852 7876
rect 57004 7916 57044 8539
rect 57196 8454 57236 8539
rect 57004 7867 57044 7876
rect 56907 7748 56949 7757
rect 56907 7708 56908 7748
rect 56948 7708 56949 7748
rect 56907 7699 56949 7708
rect 56811 7664 56853 7673
rect 56811 7624 56812 7664
rect 56852 7624 56853 7664
rect 56811 7615 56853 7624
rect 56908 7614 56948 7699
rect 56523 7580 56565 7589
rect 56523 7540 56524 7580
rect 56564 7540 56565 7580
rect 56523 7531 56565 7540
rect 56620 7160 56660 7169
rect 56428 6992 56468 7001
rect 56331 6236 56373 6245
rect 56331 6196 56332 6236
rect 56372 6196 56373 6236
rect 56331 6187 56373 6196
rect 56139 6068 56181 6077
rect 56139 6028 56140 6068
rect 56180 6028 56181 6068
rect 56139 6019 56181 6028
rect 56140 5909 56180 6019
rect 56139 5900 56181 5909
rect 56139 5860 56140 5900
rect 56180 5860 56181 5900
rect 56139 5851 56181 5860
rect 56331 5900 56373 5909
rect 56331 5860 56332 5900
rect 56372 5860 56373 5900
rect 56331 5851 56373 5860
rect 56332 5732 56372 5851
rect 56332 5683 56372 5692
rect 56428 5144 56468 6952
rect 56523 6824 56565 6833
rect 56523 6784 56524 6824
rect 56564 6784 56565 6824
rect 56523 6775 56565 6784
rect 56524 6413 56564 6775
rect 56620 6581 56660 7120
rect 57196 7160 57236 7169
rect 57004 6992 57044 7001
rect 57044 6952 57140 6992
rect 57004 6943 57044 6952
rect 57100 6581 57140 6952
rect 57196 6917 57236 7120
rect 57195 6908 57237 6917
rect 57195 6868 57196 6908
rect 57236 6868 57237 6908
rect 57195 6859 57237 6868
rect 57292 6581 57332 10051
rect 57964 10016 58004 10025
rect 58004 9976 58100 10016
rect 57964 9967 58004 9976
rect 57675 8756 57717 8765
rect 57675 8716 57676 8756
rect 57716 8716 57717 8756
rect 57675 8707 57717 8716
rect 57387 8504 57429 8513
rect 57387 8464 57388 8504
rect 57428 8464 57429 8504
rect 57387 8455 57429 8464
rect 57388 8370 57428 8455
rect 57676 7916 57716 8707
rect 57771 8420 57813 8429
rect 57771 8380 57772 8420
rect 57812 8380 57813 8420
rect 57771 8371 57813 8380
rect 57772 8177 57812 8371
rect 57771 8168 57813 8177
rect 57771 8128 57772 8168
rect 57812 8128 57813 8168
rect 57771 8119 57813 8128
rect 57676 7673 57716 7876
rect 57867 7916 57909 7925
rect 57867 7876 57868 7916
rect 57908 7876 57909 7916
rect 57867 7867 57909 7876
rect 57868 7782 57908 7867
rect 57772 7748 57812 7757
rect 57675 7664 57717 7673
rect 57675 7624 57676 7664
rect 57716 7624 57717 7664
rect 57675 7615 57717 7624
rect 57772 7589 57812 7708
rect 57771 7580 57813 7589
rect 57771 7540 57772 7580
rect 57812 7540 57813 7580
rect 57771 7531 57813 7540
rect 57867 6992 57909 7001
rect 57867 6952 57868 6992
rect 57908 6952 57909 6992
rect 57867 6943 57909 6952
rect 57675 6908 57717 6917
rect 57675 6868 57676 6908
rect 57716 6868 57717 6908
rect 57675 6859 57717 6868
rect 56619 6572 56661 6581
rect 57004 6572 57044 6581
rect 56619 6532 56620 6572
rect 56660 6532 56661 6572
rect 56619 6523 56661 6532
rect 56716 6532 57004 6572
rect 56523 6404 56565 6413
rect 56523 6364 56524 6404
rect 56564 6364 56565 6404
rect 56523 6355 56565 6364
rect 56716 6404 56756 6532
rect 57004 6523 57044 6532
rect 57099 6572 57141 6581
rect 57099 6532 57100 6572
rect 57140 6532 57141 6572
rect 57099 6523 57141 6532
rect 57291 6572 57333 6581
rect 57291 6532 57292 6572
rect 57332 6532 57333 6572
rect 57291 6523 57333 6532
rect 57483 6488 57525 6497
rect 57483 6448 57484 6488
rect 57524 6448 57525 6488
rect 57483 6439 57525 6448
rect 56524 5909 56564 6355
rect 56716 6329 56756 6364
rect 57003 6404 57045 6413
rect 57003 6364 57004 6404
rect 57044 6364 57045 6404
rect 57003 6355 57045 6364
rect 57388 6404 57428 6415
rect 56620 6320 56660 6329
rect 56620 6161 56660 6280
rect 56715 6320 56757 6329
rect 56715 6280 56716 6320
rect 56756 6280 56757 6320
rect 56715 6271 56757 6280
rect 57004 6270 57044 6355
rect 57388 6329 57428 6364
rect 57484 6354 57524 6439
rect 57579 6404 57621 6413
rect 57579 6364 57580 6404
rect 57620 6364 57621 6404
rect 57579 6355 57621 6364
rect 57387 6320 57429 6329
rect 57387 6280 57388 6320
rect 57428 6280 57429 6320
rect 57387 6271 57429 6280
rect 57580 6270 57620 6355
rect 57195 6236 57237 6245
rect 57195 6196 57196 6236
rect 57236 6196 57237 6236
rect 57195 6187 57237 6196
rect 56619 6152 56661 6161
rect 56619 6112 56620 6152
rect 56660 6112 56661 6152
rect 56619 6103 56661 6112
rect 57196 6102 57236 6187
rect 57676 6077 57716 6859
rect 57868 6497 57908 6943
rect 57867 6488 57909 6497
rect 57867 6448 57868 6488
rect 57908 6448 57909 6488
rect 57867 6439 57909 6448
rect 57964 6488 58004 6497
rect 57964 6245 58004 6448
rect 57772 6236 57812 6245
rect 57675 6068 57717 6077
rect 57675 6028 57676 6068
rect 57716 6028 57717 6068
rect 57675 6019 57717 6028
rect 56812 5909 56852 5994
rect 56523 5900 56565 5909
rect 56811 5900 56853 5909
rect 56523 5860 56524 5900
rect 56564 5860 56660 5900
rect 56523 5851 56565 5860
rect 56620 5816 56660 5860
rect 56811 5860 56812 5900
rect 56852 5860 56853 5900
rect 56811 5851 56853 5860
rect 57676 5825 57716 5835
rect 57675 5816 57717 5825
rect 56620 5776 56756 5816
rect 56524 5732 56564 5741
rect 56716 5732 56756 5776
rect 57675 5776 57676 5816
rect 57716 5776 57717 5816
rect 57675 5767 57717 5776
rect 56564 5692 56660 5732
rect 56524 5683 56564 5692
rect 56523 5564 56565 5573
rect 56523 5524 56524 5564
rect 56564 5524 56565 5564
rect 56523 5515 56565 5524
rect 56524 5430 56564 5515
rect 55852 5104 55988 5144
rect 56236 5104 56468 5144
rect 55756 4976 55796 4985
rect 55756 4565 55796 4936
rect 55852 4724 55892 5104
rect 55948 4901 55988 4986
rect 55947 4892 55989 4901
rect 55947 4852 55948 4892
rect 55988 4852 55989 4892
rect 55947 4843 55989 4852
rect 56140 4892 56180 4901
rect 56044 4808 56084 4817
rect 55852 4684 55988 4724
rect 55755 4556 55797 4565
rect 55755 4516 55756 4556
rect 55796 4516 55797 4556
rect 55755 4507 55797 4516
rect 55660 4264 55796 4304
rect 55659 4136 55701 4145
rect 55659 4096 55660 4136
rect 55700 4096 55701 4136
rect 55659 4087 55701 4096
rect 55660 4002 55700 4087
rect 55660 3464 55700 3473
rect 55756 3464 55796 4264
rect 55851 3968 55893 3977
rect 55851 3928 55852 3968
rect 55892 3928 55893 3968
rect 55851 3919 55893 3928
rect 55852 3834 55892 3919
rect 55700 3424 55796 3464
rect 55660 3415 55700 3424
rect 55851 3212 55893 3221
rect 55851 3172 55852 3212
rect 55892 3172 55893 3212
rect 55851 3163 55893 3172
rect 55852 3078 55892 3163
rect 55564 2500 55796 2540
rect 55756 2381 55796 2500
rect 55755 2372 55797 2381
rect 55755 2332 55756 2372
rect 55796 2332 55797 2372
rect 55755 2323 55797 2332
rect 55467 1280 55509 1289
rect 55467 1240 55468 1280
rect 55508 1240 55509 1280
rect 55467 1231 55509 1240
rect 55755 776 55797 785
rect 55755 736 55756 776
rect 55796 736 55797 776
rect 55755 727 55797 736
rect 55563 272 55605 281
rect 55563 232 55564 272
rect 55604 232 55605 272
rect 55563 223 55605 232
rect 55564 80 55604 223
rect 55756 80 55796 727
rect 55948 80 55988 4684
rect 56044 4472 56084 4768
rect 56140 4640 56180 4852
rect 56236 4724 56276 5104
rect 56332 4901 56372 4986
rect 56428 4979 56468 4985
rect 56620 4979 56660 5692
rect 56716 5683 56756 5692
rect 56907 5732 56949 5741
rect 57292 5732 57332 5741
rect 56907 5692 56908 5732
rect 56948 5692 57044 5732
rect 56907 5683 56949 5692
rect 56908 5598 56948 5683
rect 56716 5060 56756 5069
rect 56716 4985 56756 5020
rect 56908 4985 56948 5070
rect 56428 4976 56660 4979
rect 56468 4939 56660 4976
rect 56428 4927 56468 4936
rect 56331 4892 56373 4901
rect 56331 4852 56332 4892
rect 56372 4852 56373 4892
rect 56331 4843 56373 4852
rect 56524 4871 56564 4880
rect 56524 4733 56564 4831
rect 56620 4817 56660 4939
rect 56714 4976 56756 4985
rect 56714 4936 56715 4976
rect 56755 4936 56756 4976
rect 56714 4927 56756 4936
rect 56907 4976 56949 4985
rect 56907 4936 56908 4976
rect 56948 4936 56949 4976
rect 56907 4927 56949 4936
rect 57004 4892 57044 5692
rect 57196 5692 57292 5732
rect 57100 5480 57140 5489
rect 57100 5237 57140 5440
rect 57099 5228 57141 5237
rect 57099 5188 57100 5228
rect 57140 5188 57141 5228
rect 57099 5179 57141 5188
rect 57100 4892 57140 4901
rect 57004 4852 57100 4892
rect 57196 4892 57236 5692
rect 57292 5683 57332 5692
rect 57387 5732 57429 5741
rect 57387 5692 57388 5732
rect 57428 5692 57429 5732
rect 57387 5683 57429 5692
rect 57676 5740 57716 5767
rect 57676 5691 57716 5700
rect 57292 5590 57332 5599
rect 57292 5321 57332 5550
rect 57388 5480 57428 5683
rect 57676 5564 57716 5573
rect 57658 5524 57676 5564
rect 57658 5515 57716 5524
rect 57658 5480 57698 5515
rect 57388 5440 57698 5480
rect 57291 5312 57333 5321
rect 57291 5272 57292 5312
rect 57332 5272 57333 5312
rect 57291 5263 57333 5272
rect 57483 5060 57525 5069
rect 57483 5020 57484 5060
rect 57524 5020 57525 5060
rect 57483 5011 57525 5020
rect 57292 4892 57332 4901
rect 57484 4892 57524 5011
rect 57196 4852 57292 4892
rect 57100 4843 57140 4852
rect 56619 4808 56661 4817
rect 56619 4768 56620 4808
rect 56660 4768 56661 4808
rect 56619 4759 56661 4768
rect 56523 4724 56565 4733
rect 56236 4684 56372 4724
rect 56140 4600 56276 4640
rect 56236 4481 56276 4600
rect 56235 4472 56277 4481
rect 56044 4432 56180 4472
rect 56043 4304 56085 4313
rect 56043 4264 56044 4304
rect 56084 4264 56085 4304
rect 56043 4255 56085 4264
rect 56044 4136 56084 4255
rect 56044 4087 56084 4096
rect 56140 4061 56180 4432
rect 56235 4432 56236 4472
rect 56276 4432 56277 4472
rect 56235 4423 56277 4432
rect 56139 4052 56181 4061
rect 56139 4012 56140 4052
rect 56180 4012 56181 4052
rect 56139 4003 56181 4012
rect 56043 3632 56085 3641
rect 56043 3592 56044 3632
rect 56084 3592 56085 3632
rect 56043 3583 56085 3592
rect 56044 3464 56084 3583
rect 56044 3415 56084 3424
rect 56236 3212 56276 3221
rect 56236 1373 56276 3172
rect 56235 1364 56277 1373
rect 56235 1324 56236 1364
rect 56276 1324 56277 1364
rect 56235 1315 56277 1324
rect 56139 1028 56181 1037
rect 56139 988 56140 1028
rect 56180 988 56181 1028
rect 56139 979 56181 988
rect 56140 80 56180 979
rect 56332 80 56372 4684
rect 56523 4684 56524 4724
rect 56564 4684 56565 4724
rect 56523 4675 56565 4684
rect 56524 4229 56564 4314
rect 56523 4220 56565 4229
rect 56523 4180 56524 4220
rect 56564 4180 56565 4220
rect 56523 4171 56565 4180
rect 56523 4052 56565 4061
rect 56523 4012 56524 4052
rect 56564 4012 56565 4052
rect 56620 4052 56660 4759
rect 57292 4733 57332 4852
rect 57388 4852 57484 4892
rect 57099 4724 57141 4733
rect 57196 4724 57236 4733
rect 57099 4684 57100 4724
rect 57140 4684 57196 4724
rect 57099 4675 57141 4684
rect 57196 4675 57236 4684
rect 57291 4724 57333 4733
rect 57291 4684 57292 4724
rect 57332 4684 57333 4724
rect 57291 4675 57333 4684
rect 56715 4472 56757 4481
rect 56715 4432 56716 4472
rect 56756 4432 56757 4472
rect 56715 4423 56757 4432
rect 57003 4472 57045 4481
rect 57003 4432 57004 4472
rect 57044 4432 57045 4472
rect 57003 4423 57045 4432
rect 56716 4388 56756 4423
rect 56716 4337 56756 4348
rect 57004 4220 57044 4423
rect 57100 4229 57140 4248
rect 57099 4220 57141 4229
rect 57044 4180 57100 4220
rect 57140 4180 57141 4220
rect 57292 4220 57332 4675
rect 57388 4481 57428 4852
rect 57484 4843 57524 4852
rect 57675 4892 57717 4901
rect 57675 4852 57676 4892
rect 57716 4852 57717 4892
rect 57675 4843 57717 4852
rect 57580 4724 57620 4733
rect 57580 4481 57620 4684
rect 57387 4472 57429 4481
rect 57387 4432 57388 4472
rect 57428 4432 57429 4472
rect 57387 4423 57429 4432
rect 57579 4472 57621 4481
rect 57579 4432 57580 4472
rect 57620 4432 57621 4472
rect 57579 4423 57621 4432
rect 57580 4220 57620 4229
rect 57292 4207 57527 4220
rect 57292 4180 57580 4207
rect 57004 4171 57044 4180
rect 57099 4171 57141 4180
rect 57487 4167 57620 4180
rect 57495 4078 57535 4167
rect 57004 4052 57332 4078
rect 56620 4012 57004 4052
rect 57044 4038 57332 4052
rect 56523 4003 56565 4012
rect 57004 4003 57044 4012
rect 56427 3968 56469 3977
rect 56427 3928 56428 3968
rect 56468 3928 56469 3968
rect 56427 3919 56469 3928
rect 56428 3464 56468 3919
rect 56524 3918 56564 4003
rect 57196 3968 57236 3977
rect 57196 3632 57236 3928
rect 57195 3592 57236 3632
rect 57195 3548 57235 3592
rect 57292 3548 57332 4038
rect 57484 4038 57535 4078
rect 57579 4052 57621 4061
rect 57676 4052 57716 4843
rect 57387 3968 57429 3977
rect 57387 3928 57388 3968
rect 57428 3928 57429 3968
rect 57387 3919 57429 3928
rect 57388 3834 57428 3919
rect 57195 3508 57236 3548
rect 56428 3415 56468 3424
rect 56812 3464 56852 3473
rect 56812 3221 56852 3424
rect 56907 3464 56949 3473
rect 56907 3424 56908 3464
rect 56948 3424 56949 3464
rect 56907 3415 56949 3424
rect 56620 3212 56660 3221
rect 56620 1625 56660 3172
rect 56811 3212 56853 3221
rect 56811 3172 56812 3212
rect 56852 3172 56853 3212
rect 56811 3163 56853 3172
rect 56715 1784 56757 1793
rect 56715 1744 56716 1784
rect 56756 1744 56757 1784
rect 56715 1735 56757 1744
rect 56619 1616 56661 1625
rect 56619 1576 56620 1616
rect 56660 1576 56661 1616
rect 56619 1567 56661 1576
rect 56523 1112 56565 1121
rect 56523 1072 56524 1112
rect 56564 1072 56565 1112
rect 56523 1063 56565 1072
rect 56524 80 56564 1063
rect 56716 80 56756 1735
rect 56908 80 56948 3415
rect 57196 3389 57236 3508
rect 57292 3499 57332 3508
rect 57195 3380 57237 3389
rect 57195 3340 57196 3380
rect 57236 3340 57237 3380
rect 57195 3331 57237 3340
rect 57292 3380 57332 3389
rect 57484 3380 57524 4038
rect 57579 4012 57580 4052
rect 57620 4012 57716 4052
rect 57579 4003 57621 4012
rect 57580 3918 57620 4003
rect 57772 3632 57812 6196
rect 57963 6236 58005 6245
rect 57963 6196 57964 6236
rect 58004 6196 58005 6236
rect 57963 6187 58005 6196
rect 58060 6068 58100 9976
rect 58444 9966 58484 10051
rect 58636 9689 58676 10051
rect 58635 9680 58677 9689
rect 58635 9640 58636 9680
rect 58676 9640 58677 9680
rect 58635 9631 58677 9640
rect 58732 9605 58772 9690
rect 58731 9596 58773 9605
rect 58731 9556 58732 9596
rect 58772 9556 58773 9596
rect 58731 9547 58773 9556
rect 58155 9428 58197 9437
rect 58155 9388 58156 9428
rect 58196 9388 58197 9428
rect 58155 9379 58197 9388
rect 58732 9428 58772 9437
rect 58828 9428 58868 10144
rect 59020 10109 59060 10228
rect 59116 10219 59156 10228
rect 59019 10100 59061 10109
rect 59019 10060 59020 10100
rect 59060 10060 59061 10100
rect 59019 10051 59061 10060
rect 59116 10016 59156 10025
rect 59116 9437 59156 9976
rect 59403 9680 59445 9689
rect 59403 9640 59404 9680
rect 59444 9640 59445 9680
rect 59403 9631 59445 9640
rect 59211 9596 59253 9605
rect 59211 9556 59212 9596
rect 59252 9556 59253 9596
rect 59211 9547 59253 9556
rect 59020 9428 59060 9437
rect 58772 9388 59020 9428
rect 57964 6028 58100 6068
rect 57867 5564 57909 5573
rect 57867 5524 57868 5564
rect 57908 5524 57909 5564
rect 57867 5515 57909 5524
rect 57868 5430 57908 5515
rect 57867 5312 57909 5321
rect 57867 5272 57868 5312
rect 57908 5272 57909 5312
rect 57867 5263 57909 5272
rect 57868 5144 57908 5263
rect 57868 5095 57908 5104
rect 57964 4985 58004 6028
rect 58060 5480 58100 5489
rect 58060 5060 58100 5440
rect 58156 5321 58196 9379
rect 58540 9260 58580 9269
rect 58580 9220 58676 9260
rect 58540 9211 58580 9220
rect 58443 8084 58485 8093
rect 58443 8044 58444 8084
rect 58484 8044 58485 8084
rect 58443 8035 58485 8044
rect 58347 8000 58389 8009
rect 58347 7960 58348 8000
rect 58388 7960 58389 8000
rect 58347 7951 58389 7960
rect 58251 7916 58293 7925
rect 58251 7876 58252 7916
rect 58292 7876 58293 7916
rect 58251 7867 58293 7876
rect 58252 7076 58292 7867
rect 58348 7866 58388 7951
rect 58444 7916 58484 8035
rect 58444 7867 58484 7876
rect 58347 7664 58389 7673
rect 58347 7624 58348 7664
rect 58388 7624 58389 7664
rect 58347 7615 58389 7624
rect 58348 7244 58388 7615
rect 58348 7195 58388 7204
rect 58348 7076 58388 7085
rect 58252 7036 58348 7076
rect 58348 7027 58388 7036
rect 58539 6992 58581 7001
rect 58539 6952 58540 6992
rect 58580 6952 58581 6992
rect 58539 6943 58581 6952
rect 58540 6858 58580 6943
rect 58251 6404 58293 6413
rect 58251 6364 58252 6404
rect 58292 6364 58293 6404
rect 58251 6355 58293 6364
rect 58443 6404 58485 6413
rect 58443 6364 58444 6404
rect 58484 6364 58485 6404
rect 58636 6404 58676 9220
rect 58732 8924 58772 9388
rect 59020 9379 59060 9388
rect 59115 9428 59157 9437
rect 59115 9388 59116 9428
rect 59156 9388 59157 9428
rect 59115 9379 59157 9388
rect 59212 9428 59252 9547
rect 59212 9379 59252 9388
rect 59404 9428 59444 9631
rect 59404 9379 59444 9388
rect 59595 9428 59637 9437
rect 59595 9388 59596 9428
rect 59636 9388 59637 9428
rect 59595 9379 59637 9388
rect 59596 9294 59636 9379
rect 58732 8875 58772 8884
rect 59116 9260 59156 9269
rect 58924 8765 58964 8796
rect 58923 8756 58965 8765
rect 58923 8716 58924 8756
rect 58964 8716 58965 8756
rect 58923 8707 58965 8716
rect 58924 8672 58964 8707
rect 58924 8252 58964 8632
rect 58924 8212 59060 8252
rect 58731 8168 58773 8177
rect 58731 8128 58732 8168
rect 58772 8128 58773 8168
rect 58731 8119 58773 8128
rect 58732 8034 58772 8119
rect 58924 8084 58964 8093
rect 58828 8044 58924 8084
rect 58828 7925 58868 8044
rect 58924 8035 58964 8044
rect 58827 7916 58869 7925
rect 58827 7876 58828 7916
rect 58868 7876 58869 7916
rect 58827 7867 58869 7876
rect 58924 7916 58964 7925
rect 59020 7916 59060 8212
rect 58964 7876 59060 7916
rect 58827 7748 58869 7757
rect 58827 7708 58828 7748
rect 58868 7708 58869 7748
rect 58827 7699 58869 7708
rect 58828 6488 58868 7699
rect 58828 6439 58868 6448
rect 58924 6413 58964 7876
rect 58923 6404 58965 6413
rect 58636 6364 58772 6404
rect 58443 6355 58485 6364
rect 58252 5732 58292 6355
rect 58444 6270 58484 6355
rect 58636 6236 58676 6245
rect 58292 5692 58388 5732
rect 58252 5683 58292 5692
rect 58252 5564 58292 5575
rect 58252 5489 58292 5524
rect 58251 5480 58293 5489
rect 58251 5440 58252 5480
rect 58292 5440 58293 5480
rect 58251 5431 58293 5440
rect 58155 5312 58197 5321
rect 58155 5272 58156 5312
rect 58196 5272 58197 5312
rect 58155 5263 58197 5272
rect 58060 5020 58196 5060
rect 57963 4976 58005 4985
rect 57963 4936 57964 4976
rect 58004 4936 58005 4976
rect 57963 4927 58005 4936
rect 57868 4892 57908 4903
rect 57868 4817 57908 4852
rect 58060 4892 58100 4901
rect 57867 4808 57909 4817
rect 57867 4768 57868 4808
rect 57908 4768 57909 4808
rect 57867 4759 57909 4768
rect 58060 4733 58100 4852
rect 58059 4724 58101 4733
rect 58059 4684 58060 4724
rect 58100 4684 58101 4724
rect 58059 4675 58101 4684
rect 57963 4220 58005 4229
rect 57963 4180 57964 4220
rect 58004 4180 58005 4220
rect 57963 4171 58005 4180
rect 57964 4086 58004 4171
rect 58059 4136 58101 4145
rect 58059 4096 58060 4136
rect 58100 4096 58101 4136
rect 58059 4087 58101 4096
rect 57772 3592 57908 3632
rect 57771 3464 57813 3473
rect 57771 3424 57772 3464
rect 57812 3424 57813 3464
rect 57771 3415 57813 3424
rect 57332 3340 57524 3380
rect 57292 3331 57332 3340
rect 57772 3330 57812 3415
rect 57099 3212 57141 3221
rect 57099 3172 57100 3212
rect 57140 3172 57141 3212
rect 57099 3163 57141 3172
rect 57580 3212 57620 3221
rect 57100 3078 57140 3163
rect 57099 2792 57141 2801
rect 57099 2752 57100 2792
rect 57140 2752 57141 2792
rect 57099 2743 57141 2752
rect 57100 80 57140 2743
rect 57291 2204 57333 2213
rect 57291 2164 57292 2204
rect 57332 2164 57333 2204
rect 57291 2155 57333 2164
rect 57292 80 57332 2155
rect 57483 1616 57525 1625
rect 57483 1576 57484 1616
rect 57524 1576 57525 1616
rect 57483 1567 57525 1576
rect 57484 80 57524 1567
rect 57580 1541 57620 3172
rect 57868 2801 57908 3592
rect 57964 3212 58004 3221
rect 57867 2792 57909 2801
rect 57867 2752 57868 2792
rect 57908 2752 57909 2792
rect 57867 2743 57909 2752
rect 57675 2708 57717 2717
rect 57675 2668 57676 2708
rect 57716 2668 57717 2708
rect 57675 2659 57717 2668
rect 57579 1532 57621 1541
rect 57579 1492 57580 1532
rect 57620 1492 57621 1532
rect 57579 1483 57621 1492
rect 57676 80 57716 2659
rect 57964 1709 58004 3172
rect 58060 2456 58100 4087
rect 58156 3641 58196 5020
rect 58251 4892 58293 4901
rect 58251 4852 58252 4892
rect 58292 4852 58293 4892
rect 58348 4892 58388 5692
rect 58540 5480 58580 5489
rect 58444 4901 58484 4986
rect 58443 4892 58485 4901
rect 58348 4852 58444 4892
rect 58484 4852 58485 4892
rect 58251 4843 58293 4852
rect 58443 4843 58485 4852
rect 58252 4758 58292 4843
rect 58348 4724 58388 4733
rect 58348 4313 58388 4684
rect 58443 4724 58485 4733
rect 58443 4684 58444 4724
rect 58484 4684 58485 4724
rect 58443 4675 58485 4684
rect 58444 4565 58484 4675
rect 58443 4556 58485 4565
rect 58443 4516 58444 4556
rect 58484 4516 58485 4556
rect 58443 4507 58485 4516
rect 58347 4304 58389 4313
rect 58347 4264 58348 4304
rect 58388 4264 58389 4304
rect 58347 4255 58389 4264
rect 58540 4145 58580 5440
rect 58636 4892 58676 6196
rect 58732 5816 58772 6364
rect 58923 6364 58924 6404
rect 58964 6364 58965 6404
rect 58923 6355 58965 6364
rect 59116 6329 59156 9220
rect 59500 9260 59540 9269
rect 59212 8756 59252 8765
rect 59212 8093 59252 8716
rect 59307 8504 59349 8513
rect 59307 8464 59308 8504
rect 59348 8464 59349 8504
rect 59307 8455 59349 8464
rect 59211 8084 59253 8093
rect 59211 8044 59212 8084
rect 59252 8044 59253 8084
rect 59211 8035 59253 8044
rect 59212 7244 59252 7253
rect 59212 6833 59252 7204
rect 59308 6992 59348 8455
rect 59500 8093 59540 9220
rect 59595 9092 59637 9101
rect 59595 9052 59596 9092
rect 59636 9052 59637 9092
rect 59595 9043 59637 9052
rect 59499 8084 59541 8093
rect 59499 8044 59500 8084
rect 59540 8044 59541 8084
rect 59499 8035 59541 8044
rect 59500 7916 59540 7925
rect 59500 7673 59540 7876
rect 59499 7664 59541 7673
rect 59499 7624 59500 7664
rect 59540 7624 59541 7664
rect 59499 7615 59541 7624
rect 59596 7496 59636 9043
rect 59692 8849 59732 11899
rect 60940 11360 60980 14920
rect 64168 11360 64536 11369
rect 60940 11320 61076 11360
rect 61036 10940 61076 11320
rect 64208 11320 64250 11360
rect 64290 11320 64332 11360
rect 64372 11320 64414 11360
rect 64454 11320 64496 11360
rect 71884 11360 71924 14920
rect 79288 11360 79656 11369
rect 71884 11320 72020 11360
rect 64168 11311 64536 11320
rect 61036 10891 61076 10900
rect 61228 10940 61268 10949
rect 60075 10436 60117 10445
rect 60075 10396 60076 10436
rect 60116 10396 60117 10436
rect 60075 10387 60117 10396
rect 60363 10436 60405 10445
rect 60363 10396 60364 10436
rect 60404 10396 60405 10436
rect 60363 10387 60405 10396
rect 59884 10268 59924 10277
rect 59788 10228 59884 10268
rect 59788 9428 59828 10228
rect 59884 10219 59924 10228
rect 60076 10268 60116 10387
rect 60076 10219 60116 10228
rect 60268 10268 60308 10277
rect 60075 10100 60117 10109
rect 60075 10060 60076 10100
rect 60116 10060 60117 10100
rect 60075 10051 60117 10060
rect 60076 9966 60116 10051
rect 59883 9680 59925 9689
rect 59883 9640 59884 9680
rect 59924 9640 59925 9680
rect 59883 9631 59925 9640
rect 59884 9596 59924 9631
rect 59884 9545 59924 9556
rect 59883 9428 59925 9437
rect 59788 9388 59884 9428
rect 59924 9388 59925 9428
rect 60268 9428 60308 10228
rect 60364 9596 60404 10387
rect 60460 10268 60500 10277
rect 60460 10184 60500 10228
rect 60460 10144 60596 10184
rect 60556 10100 60596 10144
rect 60556 10060 60884 10100
rect 60460 10016 60500 10025
rect 60500 9976 60692 10016
rect 60460 9967 60500 9976
rect 60459 9764 60501 9773
rect 60459 9724 60460 9764
rect 60500 9724 60501 9764
rect 60459 9715 60501 9724
rect 60364 9547 60404 9556
rect 60363 9428 60405 9437
rect 60268 9388 60364 9428
rect 60404 9388 60405 9428
rect 59883 9379 59925 9388
rect 60363 9379 60405 9388
rect 59884 9101 59924 9379
rect 60076 9260 60116 9269
rect 60116 9220 60308 9260
rect 60076 9211 60116 9220
rect 59883 9092 59925 9101
rect 59883 9052 59884 9092
rect 59924 9052 59925 9092
rect 59883 9043 59925 9052
rect 60171 9092 60213 9101
rect 60171 9052 60172 9092
rect 60212 9052 60213 9092
rect 60171 9043 60213 9052
rect 59691 8840 59733 8849
rect 59691 8800 59692 8840
rect 59732 8800 59733 8840
rect 59691 8791 59733 8800
rect 60075 8756 60117 8765
rect 60075 8716 60076 8756
rect 60116 8716 60117 8756
rect 60075 8707 60117 8716
rect 60076 8622 60116 8707
rect 60172 8168 60212 9043
rect 60172 8119 60212 8128
rect 59980 8000 60020 8009
rect 59500 7456 59636 7496
rect 59692 7916 59732 7925
rect 59980 7916 60020 7960
rect 59732 7876 60020 7916
rect 59403 7412 59445 7421
rect 59403 7372 59404 7412
rect 59444 7372 59445 7412
rect 59403 7363 59445 7372
rect 59404 7244 59444 7363
rect 59500 7261 59540 7456
rect 59692 7421 59732 7876
rect 59883 7748 59925 7757
rect 59883 7708 59884 7748
rect 59924 7708 59925 7748
rect 59883 7699 59925 7708
rect 59691 7412 59733 7421
rect 59788 7412 59828 7421
rect 59691 7372 59692 7412
rect 59732 7372 59788 7412
rect 59691 7363 59733 7372
rect 59788 7363 59828 7372
rect 59500 7221 59636 7261
rect 59404 7195 59444 7204
rect 59308 6952 59540 6992
rect 59211 6824 59253 6833
rect 59211 6784 59212 6824
rect 59252 6784 59253 6824
rect 59211 6775 59253 6784
rect 59307 6656 59349 6665
rect 59307 6616 59308 6656
rect 59348 6616 59349 6656
rect 59307 6607 59349 6616
rect 59308 6522 59348 6607
rect 59115 6320 59157 6329
rect 59115 6280 59116 6320
rect 59156 6280 59157 6320
rect 59115 6271 59157 6280
rect 59115 5984 59157 5993
rect 59115 5944 59116 5984
rect 59156 5944 59157 5984
rect 59115 5935 59157 5944
rect 58732 5776 59060 5816
rect 58732 5648 58772 5657
rect 58732 5153 58772 5608
rect 58924 5480 58964 5489
rect 58731 5144 58773 5153
rect 58731 5104 58732 5144
rect 58772 5104 58773 5144
rect 58731 5095 58773 5104
rect 58828 4976 58868 4985
rect 58636 4852 58772 4892
rect 58636 4724 58676 4733
rect 58539 4136 58581 4145
rect 58539 4096 58540 4136
rect 58580 4096 58581 4136
rect 58539 4087 58581 4096
rect 58539 3884 58581 3893
rect 58539 3844 58540 3884
rect 58580 3844 58581 3884
rect 58539 3835 58581 3844
rect 58251 3800 58293 3809
rect 58251 3760 58252 3800
rect 58292 3760 58293 3800
rect 58251 3751 58293 3760
rect 58155 3632 58197 3641
rect 58155 3592 58156 3632
rect 58196 3592 58197 3632
rect 58155 3583 58197 3592
rect 58155 3464 58197 3473
rect 58155 3424 58156 3464
rect 58196 3424 58197 3464
rect 58155 3415 58197 3424
rect 58156 3330 58196 3415
rect 58060 2416 58196 2456
rect 58059 2288 58101 2297
rect 58059 2248 58060 2288
rect 58100 2248 58101 2288
rect 58059 2239 58101 2248
rect 57963 1700 58005 1709
rect 57963 1660 57964 1700
rect 58004 1660 58005 1700
rect 57963 1651 58005 1660
rect 57867 1448 57909 1457
rect 57867 1408 57868 1448
rect 57908 1408 57909 1448
rect 57867 1399 57909 1408
rect 57868 80 57908 1399
rect 58060 80 58100 2239
rect 58156 2213 58196 2416
rect 58155 2204 58197 2213
rect 58155 2164 58156 2204
rect 58196 2164 58197 2204
rect 58155 2155 58197 2164
rect 58252 80 58292 3751
rect 58540 3464 58580 3835
rect 58540 3415 58580 3424
rect 58348 3212 58388 3221
rect 58348 281 58388 3172
rect 58443 2204 58485 2213
rect 58443 2164 58444 2204
rect 58484 2164 58485 2204
rect 58443 2155 58485 2164
rect 58347 272 58389 281
rect 58347 232 58348 272
rect 58388 232 58389 272
rect 58347 223 58389 232
rect 58444 80 58484 2155
rect 58636 1448 58676 4684
rect 58732 3809 58772 4852
rect 58828 4397 58868 4936
rect 58827 4388 58869 4397
rect 58827 4348 58828 4388
rect 58868 4348 58869 4388
rect 58827 4339 58869 4348
rect 58827 4220 58869 4229
rect 58827 4180 58828 4220
rect 58868 4180 58869 4220
rect 58827 4171 58869 4180
rect 58828 4086 58868 4171
rect 58731 3800 58773 3809
rect 58731 3760 58732 3800
rect 58772 3760 58773 3800
rect 58731 3751 58773 3760
rect 58924 3632 58964 5440
rect 59020 4901 59060 5776
rect 59116 5648 59156 5935
rect 59116 5599 59156 5608
rect 59500 5648 59540 6952
rect 59596 6161 59636 7221
rect 59787 7244 59829 7253
rect 59787 7204 59788 7244
rect 59828 7204 59829 7244
rect 59787 7195 59829 7204
rect 59788 7110 59828 7195
rect 59787 6992 59829 7001
rect 59787 6952 59788 6992
rect 59828 6952 59829 6992
rect 59787 6943 59829 6952
rect 59595 6152 59637 6161
rect 59595 6112 59596 6152
rect 59636 6112 59637 6152
rect 59595 6103 59637 6112
rect 59788 5648 59828 6943
rect 59884 6404 59924 7699
rect 60268 7412 60308 9220
rect 60364 9101 60404 9379
rect 60363 9092 60405 9101
rect 60363 9052 60364 9092
rect 60404 9052 60405 9092
rect 60363 9043 60405 9052
rect 60460 8849 60500 9715
rect 60652 9344 60692 9976
rect 60844 9605 60884 10060
rect 60843 9596 60885 9605
rect 60843 9556 60844 9596
rect 60884 9556 60885 9596
rect 60843 9547 60885 9556
rect 60843 9428 60885 9437
rect 60843 9388 60844 9428
rect 60884 9388 60885 9428
rect 60843 9379 60885 9388
rect 60652 9304 60788 9344
rect 60556 9260 60596 9269
rect 60596 9220 60692 9260
rect 60556 9211 60596 9220
rect 60459 8840 60501 8849
rect 60459 8800 60460 8840
rect 60500 8800 60501 8840
rect 60459 8791 60501 8800
rect 60555 8420 60597 8429
rect 60555 8380 60556 8420
rect 60596 8380 60597 8420
rect 60555 8371 60597 8380
rect 60556 7421 60596 8371
rect 60652 7589 60692 9220
rect 60651 7580 60693 7589
rect 60651 7540 60652 7580
rect 60692 7540 60693 7580
rect 60651 7531 60693 7540
rect 60748 7505 60788 9304
rect 60844 9294 60884 9379
rect 61036 9260 61076 9269
rect 61076 9220 61172 9260
rect 61036 9211 61076 9220
rect 60843 8756 60885 8765
rect 60843 8716 60844 8756
rect 60884 8716 60885 8756
rect 60843 8707 60885 8716
rect 60747 7496 60789 7505
rect 60747 7456 60748 7496
rect 60788 7456 60789 7496
rect 60747 7447 60789 7456
rect 60172 7372 60308 7412
rect 60363 7412 60405 7421
rect 60555 7412 60597 7421
rect 60363 7372 60364 7412
rect 60404 7372 60500 7412
rect 59979 7244 60021 7253
rect 59979 7204 59980 7244
rect 60020 7204 60021 7244
rect 59979 7195 60021 7204
rect 60076 7244 60116 7253
rect 59980 7110 60020 7195
rect 59979 6992 60021 7001
rect 59979 6952 59980 6992
rect 60020 6952 60021 6992
rect 59979 6943 60021 6952
rect 59884 6355 59924 6364
rect 59884 5648 59924 5657
rect 59788 5608 59884 5648
rect 59500 5599 59540 5608
rect 59884 5599 59924 5608
rect 59308 5480 59348 5489
rect 59692 5480 59732 5489
rect 59211 4976 59253 4985
rect 59211 4936 59212 4976
rect 59252 4936 59253 4976
rect 59211 4927 59253 4936
rect 59019 4892 59061 4901
rect 59019 4852 59020 4892
rect 59060 4852 59061 4892
rect 59019 4843 59061 4852
rect 59212 4842 59252 4927
rect 58828 3592 58964 3632
rect 59020 4724 59060 4733
rect 58540 1408 58676 1448
rect 58732 3212 58772 3221
rect 58540 1037 58580 1408
rect 58635 1280 58677 1289
rect 58635 1240 58636 1280
rect 58676 1240 58677 1280
rect 58635 1231 58677 1240
rect 58539 1028 58581 1037
rect 58539 988 58540 1028
rect 58580 988 58581 1028
rect 58539 979 58581 988
rect 58636 80 58676 1231
rect 58732 785 58772 3172
rect 58828 2717 58868 3592
rect 58924 3464 58964 3473
rect 58924 3137 58964 3424
rect 58923 3128 58965 3137
rect 58923 3088 58924 3128
rect 58964 3088 58965 3128
rect 58923 3079 58965 3088
rect 58827 2708 58869 2717
rect 58827 2668 58828 2708
rect 58868 2668 58869 2708
rect 58827 2659 58869 2668
rect 58827 2540 58869 2549
rect 59020 2540 59060 4684
rect 59115 4724 59157 4733
rect 59115 4684 59116 4724
rect 59156 4684 59157 4724
rect 59115 4675 59157 4684
rect 58827 2500 58828 2540
rect 58868 2500 58869 2540
rect 58827 2491 58869 2500
rect 58924 2500 59060 2540
rect 58731 776 58773 785
rect 58731 736 58732 776
rect 58772 736 58773 776
rect 58731 727 58773 736
rect 58828 80 58868 2491
rect 58924 1121 58964 2500
rect 59019 2372 59061 2381
rect 59019 2332 59020 2372
rect 59060 2332 59061 2372
rect 59019 2323 59061 2332
rect 58923 1112 58965 1121
rect 58923 1072 58924 1112
rect 58964 1072 58965 1112
rect 58923 1063 58965 1072
rect 59020 80 59060 2323
rect 59116 2213 59156 4675
rect 59212 4220 59252 4229
rect 59212 3557 59252 4180
rect 59211 3548 59253 3557
rect 59211 3508 59212 3548
rect 59252 3508 59253 3548
rect 59211 3499 59253 3508
rect 59308 2297 59348 5440
rect 59596 5440 59692 5480
rect 59499 5312 59541 5321
rect 59499 5272 59500 5312
rect 59540 5272 59541 5312
rect 59499 5263 59541 5272
rect 59403 4976 59445 4985
rect 59403 4936 59404 4976
rect 59444 4936 59445 4976
rect 59403 4927 59445 4936
rect 59404 4229 59444 4927
rect 59500 4313 59540 5263
rect 59499 4304 59541 4313
rect 59499 4264 59500 4304
rect 59540 4264 59541 4304
rect 59499 4255 59541 4264
rect 59403 4220 59445 4229
rect 59403 4180 59404 4220
rect 59444 4180 59445 4220
rect 59403 4171 59445 4180
rect 59500 3380 59540 4255
rect 59500 3331 59540 3340
rect 59499 3212 59541 3221
rect 59499 3172 59500 3212
rect 59540 3172 59541 3212
rect 59499 3163 59541 3172
rect 59500 3078 59540 3163
rect 59499 2624 59541 2633
rect 59596 2624 59636 5440
rect 59692 5431 59732 5440
rect 59787 5480 59829 5489
rect 59787 5440 59788 5480
rect 59828 5440 59829 5480
rect 59787 5431 59829 5440
rect 59691 4976 59733 4985
rect 59691 4936 59692 4976
rect 59732 4936 59733 4976
rect 59691 4927 59733 4936
rect 59692 4892 59732 4927
rect 59692 4841 59732 4852
rect 59692 4724 59732 4733
rect 59692 3641 59732 4684
rect 59691 3632 59733 3641
rect 59691 3592 59692 3632
rect 59732 3592 59733 3632
rect 59691 3583 59733 3592
rect 59692 3380 59732 3389
rect 59692 3221 59732 3340
rect 59691 3212 59733 3221
rect 59691 3172 59692 3212
rect 59732 3172 59733 3212
rect 59691 3163 59733 3172
rect 59499 2584 59500 2624
rect 59540 2584 59636 2624
rect 59499 2575 59541 2584
rect 59788 2540 59828 5431
rect 59884 4892 59924 4901
rect 59884 4229 59924 4852
rect 59883 4220 59925 4229
rect 59883 4180 59884 4220
rect 59924 4180 59925 4220
rect 59883 4171 59925 4180
rect 59980 2717 60020 6943
rect 60076 6413 60116 7204
rect 60075 6404 60117 6413
rect 60075 6364 60076 6404
rect 60116 6364 60117 6404
rect 60075 6355 60117 6364
rect 60075 5480 60117 5489
rect 60075 5440 60076 5480
rect 60116 5440 60117 5480
rect 60075 5431 60117 5440
rect 60076 5346 60116 5431
rect 60172 5069 60212 7372
rect 60363 7363 60405 7372
rect 60460 7328 60500 7372
rect 60555 7372 60556 7412
rect 60596 7372 60597 7412
rect 60555 7363 60597 7372
rect 60844 7412 60884 8707
rect 60844 7363 60884 7372
rect 60267 7244 60309 7253
rect 60267 7204 60268 7244
rect 60308 7204 60309 7244
rect 60267 7195 60309 7204
rect 60364 7244 60410 7253
rect 60409 7204 60410 7244
rect 60364 7195 60410 7204
rect 60268 6824 60308 7195
rect 60369 7114 60409 7195
rect 60268 6784 60404 6824
rect 60267 6656 60309 6665
rect 60267 6616 60268 6656
rect 60308 6616 60309 6656
rect 60267 6607 60309 6616
rect 60268 6404 60308 6607
rect 60268 6355 60308 6364
rect 60364 6329 60404 6784
rect 60460 6413 60500 7288
rect 60556 7278 60596 7363
rect 60651 7244 60693 7253
rect 60651 7204 60652 7244
rect 60692 7204 60693 7244
rect 60651 7195 60693 7204
rect 60555 6992 60597 7001
rect 60555 6952 60556 6992
rect 60596 6952 60597 6992
rect 60555 6943 60597 6952
rect 60556 6858 60596 6943
rect 60459 6404 60501 6413
rect 60459 6364 60460 6404
rect 60500 6364 60501 6404
rect 60459 6355 60501 6364
rect 60363 6320 60405 6329
rect 60363 6280 60364 6320
rect 60404 6280 60405 6320
rect 60363 6271 60405 6280
rect 60555 6320 60597 6329
rect 60555 6280 60556 6320
rect 60596 6280 60597 6320
rect 60555 6271 60597 6280
rect 60556 6186 60596 6271
rect 60363 6152 60405 6161
rect 60363 6112 60364 6152
rect 60404 6112 60405 6152
rect 60363 6103 60405 6112
rect 60268 5648 60308 5659
rect 60268 5573 60308 5608
rect 60267 5564 60309 5573
rect 60267 5524 60268 5564
rect 60308 5524 60309 5564
rect 60267 5515 60309 5524
rect 60171 5060 60213 5069
rect 60171 5020 60172 5060
rect 60212 5020 60213 5060
rect 60171 5011 60213 5020
rect 60364 4976 60404 6103
rect 60652 6068 60692 7195
rect 61036 7160 61076 7169
rect 61036 7001 61076 7120
rect 61035 6992 61077 7001
rect 61035 6952 61036 6992
rect 61076 6952 61077 6992
rect 61035 6943 61077 6952
rect 61035 6656 61077 6665
rect 61035 6616 61036 6656
rect 61076 6616 61077 6656
rect 61035 6607 61077 6616
rect 60747 6572 60789 6581
rect 60747 6532 60748 6572
rect 60788 6532 60789 6572
rect 60747 6523 60789 6532
rect 60748 6236 60788 6523
rect 61036 6404 61076 6607
rect 61036 6355 61076 6364
rect 60748 6187 60788 6196
rect 60652 6028 60788 6068
rect 60651 5648 60693 5657
rect 60651 5608 60652 5648
rect 60692 5608 60693 5648
rect 60651 5599 60693 5608
rect 60652 5514 60692 5599
rect 60364 4927 60404 4936
rect 60460 5480 60500 5489
rect 60075 4892 60117 4901
rect 60075 4852 60076 4892
rect 60116 4852 60117 4892
rect 60075 4843 60117 4852
rect 60076 4061 60116 4843
rect 60171 4724 60213 4733
rect 60171 4684 60172 4724
rect 60212 4684 60213 4724
rect 60171 4675 60213 4684
rect 60172 4590 60212 4675
rect 60460 4472 60500 5440
rect 60748 4976 60788 6028
rect 61132 5657 61172 9220
rect 61228 8597 61268 10900
rect 61323 10940 61365 10949
rect 61323 10900 61324 10940
rect 61364 10900 61365 10940
rect 61323 10891 61365 10900
rect 71980 10940 72020 11320
rect 79328 11320 79370 11360
rect 79410 11320 79452 11360
rect 79492 11320 79534 11360
rect 79574 11320 79616 11360
rect 82828 11360 82868 14920
rect 93772 11957 93812 14920
rect 93771 11948 93813 11957
rect 93771 11908 93772 11948
rect 93812 11908 93813 11948
rect 93771 11899 93813 11908
rect 94408 11360 94776 11369
rect 82828 11320 82964 11360
rect 79288 11311 79656 11320
rect 71980 10891 72020 10900
rect 72172 10940 72212 10949
rect 82924 10940 82964 11320
rect 94448 11320 94490 11360
rect 94530 11320 94572 11360
rect 94612 11320 94654 11360
rect 94694 11320 94736 11360
rect 94408 11311 94776 11320
rect 72212 10900 72404 10940
rect 72172 10891 72212 10900
rect 61227 8588 61269 8597
rect 61227 8548 61228 8588
rect 61268 8548 61269 8588
rect 61227 8539 61269 8548
rect 61227 8420 61269 8429
rect 61227 8380 61228 8420
rect 61268 8380 61269 8420
rect 61227 8371 61269 8380
rect 61228 6572 61268 8371
rect 61324 6581 61364 10891
rect 68427 10688 68469 10697
rect 68427 10648 68428 10688
rect 68468 10648 68469 10688
rect 68427 10639 68469 10648
rect 65408 10604 65776 10613
rect 65448 10564 65490 10604
rect 65530 10564 65572 10604
rect 65612 10564 65654 10604
rect 65694 10564 65736 10604
rect 65408 10555 65776 10564
rect 68428 10268 68468 10639
rect 69771 10436 69813 10445
rect 69771 10396 69772 10436
rect 69812 10396 69813 10436
rect 69771 10387 69813 10396
rect 71307 10436 71349 10445
rect 71307 10396 71308 10436
rect 71348 10396 71349 10436
rect 71307 10387 71349 10396
rect 68428 10219 68468 10228
rect 69579 10268 69621 10277
rect 69579 10228 69580 10268
rect 69620 10228 69621 10268
rect 69579 10219 69621 10228
rect 69772 10268 69812 10387
rect 69772 10219 69812 10228
rect 71308 10268 71348 10387
rect 71308 10219 71348 10228
rect 71500 10268 71540 10277
rect 71540 10228 71636 10268
rect 71500 10219 71540 10228
rect 69580 10134 69620 10219
rect 69099 10100 69141 10109
rect 69099 10060 69100 10100
rect 69140 10060 69141 10100
rect 69099 10051 69141 10060
rect 69100 9966 69140 10051
rect 71404 10016 71444 10025
rect 64168 9848 64536 9857
rect 64208 9808 64250 9848
rect 64290 9808 64332 9848
rect 64372 9808 64414 9848
rect 64454 9808 64496 9848
rect 64168 9799 64536 9808
rect 67947 9596 67989 9605
rect 67947 9556 67948 9596
rect 67988 9556 67989 9596
rect 67947 9547 67989 9556
rect 66891 9512 66933 9521
rect 66891 9472 66892 9512
rect 66932 9472 66933 9512
rect 66891 9463 66933 9472
rect 62092 9428 62132 9437
rect 62092 9017 62132 9388
rect 65163 9428 65205 9437
rect 65163 9388 65164 9428
rect 65204 9388 65205 9428
rect 65163 9379 65205 9388
rect 66124 9428 66164 9437
rect 62956 9344 62996 9353
rect 62956 9017 62996 9304
rect 65164 9294 65204 9379
rect 63723 9260 63765 9269
rect 63723 9220 63724 9260
rect 63764 9220 63765 9260
rect 63723 9211 63765 9220
rect 62091 9008 62133 9017
rect 62091 8968 62092 9008
rect 62132 8968 62133 9008
rect 62091 8959 62133 8968
rect 62955 9008 62997 9017
rect 62955 8968 62956 9008
rect 62996 8968 62997 9008
rect 62955 8959 62997 8968
rect 62091 8336 62133 8345
rect 62091 8296 62092 8336
rect 62132 8296 62133 8336
rect 62091 8287 62133 8296
rect 62092 8009 62132 8287
rect 63627 8252 63669 8261
rect 63627 8212 63628 8252
rect 63668 8212 63669 8252
rect 63627 8203 63669 8212
rect 62091 8000 62133 8009
rect 62091 7960 62092 8000
rect 62132 7960 62133 8000
rect 62091 7951 62133 7960
rect 61707 7412 61749 7421
rect 61707 7372 61708 7412
rect 61748 7372 61749 7412
rect 61707 7363 61749 7372
rect 61804 7412 61844 7421
rect 62092 7412 62132 7951
rect 62667 7916 62709 7925
rect 62667 7876 62668 7916
rect 62708 7876 62709 7916
rect 62667 7867 62709 7876
rect 63628 7916 63668 8203
rect 63628 7867 63668 7876
rect 62668 7782 62708 7867
rect 62379 7580 62421 7589
rect 62379 7540 62380 7580
rect 62420 7540 62421 7580
rect 62379 7531 62421 7540
rect 61844 7372 62036 7412
rect 61804 7363 61844 7372
rect 61708 7244 61748 7363
rect 61899 7244 61941 7253
rect 61708 7204 61844 7244
rect 61228 6523 61268 6532
rect 61323 6572 61365 6581
rect 61323 6532 61324 6572
rect 61364 6532 61365 6572
rect 61323 6523 61365 6532
rect 61228 6404 61268 6413
rect 61324 6404 61364 6523
rect 61268 6364 61364 6404
rect 61804 6404 61844 7204
rect 61899 7204 61900 7244
rect 61940 7204 61941 7244
rect 61899 7195 61941 7204
rect 61900 7110 61940 7195
rect 61899 6572 61941 6581
rect 61899 6532 61900 6572
rect 61940 6532 61941 6572
rect 61899 6523 61941 6532
rect 61900 6413 61940 6523
rect 61228 6355 61268 6364
rect 61804 6355 61844 6364
rect 61899 6404 61941 6413
rect 61899 6364 61900 6404
rect 61940 6364 61941 6404
rect 61899 6355 61941 6364
rect 61996 6404 62036 7372
rect 62092 7363 62132 7372
rect 62187 7244 62229 7253
rect 62187 7204 62188 7244
rect 62228 7204 62229 7244
rect 62187 7195 62229 7204
rect 61419 6320 61461 6329
rect 61419 6280 61420 6320
rect 61460 6280 61461 6320
rect 61419 6271 61461 6280
rect 61227 6236 61269 6245
rect 61227 6196 61228 6236
rect 61268 6196 61269 6236
rect 61227 6187 61269 6196
rect 61228 5741 61268 6187
rect 61323 5984 61365 5993
rect 61323 5944 61324 5984
rect 61364 5944 61365 5984
rect 61323 5935 61365 5944
rect 61324 5900 61364 5935
rect 61324 5849 61364 5860
rect 61227 5732 61269 5741
rect 61227 5692 61228 5732
rect 61268 5692 61269 5732
rect 61227 5683 61269 5692
rect 61324 5732 61364 5741
rect 61420 5732 61460 6271
rect 61900 6270 61940 6355
rect 61996 5993 62036 6364
rect 62092 6404 62132 6415
rect 62092 6329 62132 6364
rect 62091 6320 62133 6329
rect 62091 6280 62092 6320
rect 62132 6280 62133 6320
rect 62091 6271 62133 6280
rect 61803 5984 61845 5993
rect 61803 5944 61804 5984
rect 61844 5944 61845 5984
rect 61803 5935 61845 5944
rect 61995 5984 62037 5993
rect 61995 5944 61996 5984
rect 62036 5944 62037 5984
rect 61995 5935 62037 5944
rect 61364 5692 61460 5732
rect 61324 5683 61364 5692
rect 61131 5648 61173 5657
rect 61131 5608 61132 5648
rect 61172 5608 61173 5648
rect 61131 5599 61173 5608
rect 61228 5598 61268 5683
rect 61804 5648 61844 5935
rect 61804 5599 61844 5608
rect 61996 5732 62036 5741
rect 62188 5732 62228 7195
rect 62284 6572 62324 6581
rect 62284 6413 62324 6532
rect 62283 6404 62325 6413
rect 62283 6364 62284 6404
rect 62324 6364 62325 6404
rect 62283 6355 62325 6364
rect 62036 5692 62228 5732
rect 61899 5564 61941 5573
rect 61899 5524 61900 5564
rect 61940 5524 61941 5564
rect 61899 5515 61941 5524
rect 61036 5480 61076 5489
rect 61076 5440 61364 5480
rect 60939 5228 60981 5237
rect 60939 5188 60940 5228
rect 60980 5188 60981 5228
rect 60939 5179 60981 5188
rect 60748 4927 60788 4936
rect 60364 4432 60500 4472
rect 60556 4724 60596 4733
rect 60171 4304 60213 4313
rect 60171 4264 60172 4304
rect 60212 4264 60213 4304
rect 60171 4255 60213 4264
rect 60172 4220 60212 4255
rect 60172 4169 60212 4180
rect 60075 4052 60117 4061
rect 60075 4012 60076 4052
rect 60116 4012 60117 4052
rect 60075 4003 60117 4012
rect 60076 3380 60116 4003
rect 60268 3557 60308 3642
rect 60267 3548 60309 3557
rect 60267 3508 60268 3548
rect 60308 3508 60309 3548
rect 60267 3499 60309 3508
rect 60076 3331 60116 3340
rect 60268 3380 60308 3389
rect 60268 3221 60308 3340
rect 60267 3212 60309 3221
rect 60267 3172 60268 3212
rect 60308 3172 60309 3212
rect 60267 3163 60309 3172
rect 59979 2708 60021 2717
rect 59979 2668 59980 2708
rect 60020 2668 60021 2708
rect 59979 2659 60021 2668
rect 60364 2549 60404 4432
rect 60460 4218 60500 4303
rect 60459 4209 60501 4218
rect 60459 4169 60460 4209
rect 60500 4169 60501 4209
rect 60459 4160 60501 4169
rect 60459 4052 60501 4061
rect 60459 4012 60460 4052
rect 60500 4012 60501 4052
rect 60459 4003 60501 4012
rect 60460 3918 60500 4003
rect 60556 3632 60596 4684
rect 60652 4220 60692 4229
rect 60652 4061 60692 4180
rect 60940 4220 60980 5179
rect 60940 4171 60980 4180
rect 61036 4220 61076 5440
rect 61324 4892 61364 5440
rect 61900 5430 61940 5515
rect 61996 5405 62036 5692
rect 62380 5648 62420 7531
rect 63051 7244 63093 7253
rect 63051 7204 63052 7244
rect 63092 7204 63093 7244
rect 63051 7195 63093 7204
rect 62475 7160 62517 7169
rect 62475 7120 62476 7160
rect 62516 7120 62517 7160
rect 62475 7111 62517 7120
rect 62476 6656 62516 7111
rect 63052 7110 63092 7195
rect 62476 6607 62516 6616
rect 62667 6404 62709 6413
rect 62667 6364 62668 6404
rect 62708 6364 62709 6404
rect 62667 6355 62709 6364
rect 62956 6404 62996 6413
rect 62668 6270 62708 6355
rect 62764 6236 62804 6245
rect 62956 6236 62996 6364
rect 63147 6404 63189 6413
rect 63147 6364 63148 6404
rect 63188 6364 63189 6404
rect 63147 6355 63189 6364
rect 62804 6196 62996 6236
rect 63052 6320 63092 6329
rect 62476 5648 62516 5657
rect 62380 5608 62476 5648
rect 62476 5599 62516 5608
rect 62284 5480 62324 5489
rect 61995 5396 62037 5405
rect 61995 5356 61996 5396
rect 62036 5356 62037 5396
rect 61995 5347 62037 5356
rect 61803 5228 61845 5237
rect 61803 5188 61804 5228
rect 61844 5188 61845 5228
rect 61803 5179 61845 5188
rect 61804 5144 61844 5179
rect 62284 5144 62324 5440
rect 62667 5480 62709 5489
rect 62667 5440 62668 5480
rect 62708 5440 62709 5480
rect 62667 5431 62709 5440
rect 62668 5346 62708 5431
rect 62764 5405 62804 6196
rect 62860 5648 62900 5657
rect 63052 5648 63092 6280
rect 63148 6270 63188 6355
rect 63244 5648 63284 5657
rect 63052 5608 63188 5648
rect 62763 5396 62805 5405
rect 62763 5356 62764 5396
rect 62804 5356 62805 5396
rect 62763 5347 62805 5356
rect 62860 5237 62900 5608
rect 62955 5564 62997 5573
rect 62955 5524 62956 5564
rect 62996 5524 62997 5564
rect 62955 5515 62997 5524
rect 62859 5228 62901 5237
rect 62859 5188 62860 5228
rect 62900 5188 62901 5228
rect 62859 5179 62901 5188
rect 61804 5093 61844 5104
rect 61900 5104 62324 5144
rect 61900 4976 61940 5104
rect 62956 5069 62996 5515
rect 63052 5480 63092 5489
rect 62763 5060 62805 5069
rect 62763 5020 62764 5060
rect 62804 5020 62805 5060
rect 62763 5011 62805 5020
rect 62955 5060 62997 5069
rect 62955 5020 62956 5060
rect 62996 5020 62997 5060
rect 62955 5011 62997 5020
rect 61804 4936 61940 4976
rect 62764 4976 62804 5011
rect 61708 4892 61748 4901
rect 61364 4852 61708 4892
rect 61324 4843 61364 4852
rect 61708 4843 61748 4852
rect 61228 4724 61268 4733
rect 61228 4565 61268 4684
rect 61516 4724 61556 4733
rect 61227 4556 61269 4565
rect 61227 4516 61228 4556
rect 61268 4516 61269 4556
rect 61227 4507 61269 4516
rect 61227 4388 61269 4397
rect 61227 4348 61228 4388
rect 61268 4348 61269 4388
rect 61227 4339 61269 4348
rect 61228 4254 61268 4339
rect 61036 4171 61076 4180
rect 60651 4052 60693 4061
rect 60651 4012 60652 4052
rect 60692 4012 60693 4052
rect 60651 4003 60693 4012
rect 61420 3968 61460 3977
rect 60651 3800 60693 3809
rect 60651 3760 60652 3800
rect 60692 3760 60693 3800
rect 60651 3751 60693 3760
rect 60460 3592 60596 3632
rect 59596 2500 59828 2540
rect 59979 2540 60021 2549
rect 59979 2500 59980 2540
rect 60020 2500 60021 2540
rect 59307 2288 59349 2297
rect 59307 2248 59308 2288
rect 59348 2248 59349 2288
rect 59307 2239 59349 2248
rect 59115 2204 59157 2213
rect 59115 2164 59116 2204
rect 59156 2164 59157 2204
rect 59115 2155 59157 2164
rect 59403 2036 59445 2045
rect 59403 1996 59404 2036
rect 59444 1996 59445 2036
rect 59403 1987 59445 1996
rect 59211 1112 59253 1121
rect 59211 1072 59212 1112
rect 59252 1072 59253 1112
rect 59211 1063 59253 1072
rect 59212 80 59252 1063
rect 59404 80 59444 1987
rect 59596 80 59636 2500
rect 59979 2491 60021 2500
rect 60363 2540 60405 2549
rect 60363 2500 60364 2540
rect 60404 2500 60405 2540
rect 60363 2491 60405 2500
rect 59787 1196 59829 1205
rect 59787 1156 59788 1196
rect 59828 1156 59829 1196
rect 59787 1147 59829 1156
rect 59788 80 59828 1147
rect 59980 80 60020 2491
rect 60460 2381 60500 3592
rect 60556 3212 60596 3221
rect 60459 2372 60501 2381
rect 60459 2332 60460 2372
rect 60500 2332 60501 2372
rect 60459 2323 60501 2332
rect 60363 1868 60405 1877
rect 60363 1828 60364 1868
rect 60404 1828 60405 1868
rect 60363 1819 60405 1828
rect 60171 860 60213 869
rect 60171 820 60172 860
rect 60212 820 60213 860
rect 60171 811 60213 820
rect 60172 80 60212 811
rect 60364 80 60404 1819
rect 60556 1793 60596 3172
rect 60555 1784 60597 1793
rect 60555 1744 60556 1784
rect 60596 1744 60597 1784
rect 60555 1735 60597 1744
rect 60652 1616 60692 3751
rect 61131 3716 61173 3725
rect 61131 3676 61132 3716
rect 61172 3676 61173 3716
rect 61131 3667 61173 3676
rect 60747 3464 60789 3473
rect 60747 3424 60748 3464
rect 60788 3424 60789 3464
rect 60747 3415 60789 3424
rect 61132 3464 61172 3667
rect 61227 3548 61269 3557
rect 61227 3508 61228 3548
rect 61268 3508 61269 3548
rect 61227 3499 61269 3508
rect 61132 3415 61172 3424
rect 60748 3330 60788 3415
rect 60747 3212 60789 3221
rect 60747 3172 60748 3212
rect 60788 3172 60789 3212
rect 60747 3163 60789 3172
rect 60940 3212 60980 3221
rect 60556 1576 60692 1616
rect 60556 80 60596 1576
rect 60748 80 60788 3163
rect 60940 1625 60980 3172
rect 61228 2885 61268 3499
rect 61324 3212 61364 3221
rect 61227 2876 61269 2885
rect 61227 2836 61228 2876
rect 61268 2836 61269 2876
rect 61227 2827 61269 2836
rect 61131 2456 61173 2465
rect 61131 2416 61132 2456
rect 61172 2416 61173 2456
rect 61131 2407 61173 2416
rect 60939 1616 60981 1625
rect 60939 1576 60940 1616
rect 60980 1576 60981 1616
rect 60939 1567 60981 1576
rect 60939 1028 60981 1037
rect 60939 988 60940 1028
rect 60980 988 60981 1028
rect 60939 979 60981 988
rect 60940 80 60980 979
rect 61132 80 61172 2407
rect 61324 1457 61364 3172
rect 61420 2045 61460 3928
rect 61516 3725 61556 4684
rect 61611 4724 61653 4733
rect 61611 4684 61612 4724
rect 61652 4684 61653 4724
rect 61611 4675 61653 4684
rect 61612 4136 61652 4675
rect 61804 4136 61844 4936
rect 62764 4925 62804 4936
rect 62092 4892 62132 4901
rect 61900 4871 61940 4880
rect 61900 4565 61940 4831
rect 61899 4556 61941 4565
rect 61899 4516 61900 4556
rect 61940 4516 61941 4556
rect 61899 4507 61941 4516
rect 61612 4087 61652 4096
rect 61708 4096 61844 4136
rect 61995 4136 62037 4145
rect 61995 4096 61996 4136
rect 62036 4096 62037 4136
rect 61515 3716 61557 3725
rect 61515 3676 61516 3716
rect 61556 3676 61557 3716
rect 61515 3667 61557 3676
rect 61516 3464 61556 3473
rect 61516 3053 61556 3424
rect 61708 3380 61748 4096
rect 61995 4087 62037 4096
rect 61996 4002 62036 4087
rect 61612 3340 61748 3380
rect 61804 3968 61844 3977
rect 61515 3044 61557 3053
rect 61515 3004 61516 3044
rect 61556 3004 61557 3044
rect 61515 2995 61557 3004
rect 61612 2540 61652 3340
rect 61516 2500 61652 2540
rect 61708 3212 61748 3221
rect 61419 2036 61461 2045
rect 61419 1996 61420 2036
rect 61460 1996 61461 2036
rect 61419 1987 61461 1996
rect 61323 1448 61365 1457
rect 61323 1408 61324 1448
rect 61364 1408 61365 1448
rect 61323 1399 61365 1408
rect 61323 944 61365 953
rect 61323 904 61324 944
rect 61364 904 61365 944
rect 61323 895 61365 904
rect 61324 80 61364 895
rect 61516 80 61556 2500
rect 61611 2204 61653 2213
rect 61611 2164 61612 2204
rect 61652 2164 61653 2204
rect 61611 2155 61653 2164
rect 61612 1112 61652 2155
rect 61708 1289 61748 3172
rect 61804 3137 61844 3928
rect 62092 3893 62132 4852
rect 62284 4892 62324 4901
rect 62284 4229 62324 4852
rect 62572 4724 62612 4733
rect 62859 4724 62901 4733
rect 62612 4684 62708 4724
rect 62572 4675 62612 4684
rect 62475 4556 62517 4565
rect 62475 4516 62476 4556
rect 62516 4516 62517 4556
rect 62475 4507 62517 4516
rect 62379 4472 62421 4481
rect 62379 4432 62380 4472
rect 62420 4432 62421 4472
rect 62379 4423 62421 4432
rect 62283 4220 62325 4229
rect 62283 4180 62284 4220
rect 62324 4180 62325 4220
rect 62283 4171 62325 4180
rect 62380 4136 62420 4423
rect 62380 4087 62420 4096
rect 62188 3968 62228 3977
rect 62228 3928 62420 3968
rect 62188 3919 62228 3928
rect 62091 3884 62133 3893
rect 62091 3844 62092 3884
rect 62132 3844 62133 3884
rect 62091 3835 62133 3844
rect 62283 3548 62325 3557
rect 62283 3508 62284 3548
rect 62324 3508 62325 3548
rect 62283 3499 62325 3508
rect 61900 3464 61940 3473
rect 62284 3464 62324 3499
rect 61940 3451 61953 3464
rect 61940 3424 62228 3451
rect 61900 3415 62228 3424
rect 61913 3411 62228 3415
rect 62284 3413 62324 3424
rect 62188 3296 62228 3411
rect 62188 3256 62324 3296
rect 62092 3212 62132 3221
rect 61803 3128 61845 3137
rect 61803 3088 61804 3128
rect 61844 3088 61845 3128
rect 61803 3079 61845 3088
rect 61995 3128 62037 3137
rect 61995 3088 61996 3128
rect 62036 3088 62037 3128
rect 61995 3079 62037 3088
rect 61899 2876 61941 2885
rect 61899 2836 61900 2876
rect 61940 2836 61941 2876
rect 61899 2827 61941 2836
rect 61707 1280 61749 1289
rect 61707 1240 61708 1280
rect 61748 1240 61749 1280
rect 61707 1231 61749 1240
rect 61612 1072 61748 1112
rect 61708 80 61748 1072
rect 61900 80 61940 2827
rect 61996 1205 62036 3079
rect 61995 1196 62037 1205
rect 61995 1156 61996 1196
rect 62036 1156 62037 1196
rect 61995 1147 62037 1156
rect 62092 1121 62132 3172
rect 62187 3128 62229 3137
rect 62187 3088 62188 3128
rect 62228 3088 62229 3128
rect 62187 3079 62229 3088
rect 62091 1112 62133 1121
rect 62091 1072 62092 1112
rect 62132 1072 62133 1112
rect 62091 1063 62133 1072
rect 62188 944 62228 3079
rect 62284 2969 62324 3256
rect 62283 2960 62325 2969
rect 62283 2920 62284 2960
rect 62324 2920 62325 2960
rect 62283 2911 62325 2920
rect 62283 2372 62325 2381
rect 62283 2332 62284 2372
rect 62324 2332 62325 2372
rect 62283 2323 62325 2332
rect 62092 904 62228 944
rect 62092 80 62132 904
rect 62284 80 62324 2323
rect 62380 869 62420 3928
rect 62379 860 62421 869
rect 62379 820 62380 860
rect 62420 820 62421 860
rect 62379 811 62421 820
rect 62476 80 62516 4507
rect 62572 3968 62612 3977
rect 62572 3809 62612 3928
rect 62571 3800 62613 3809
rect 62571 3760 62572 3800
rect 62612 3760 62613 3800
rect 62571 3751 62613 3760
rect 62571 3380 62613 3389
rect 62571 3340 62572 3380
rect 62612 3340 62613 3380
rect 62571 3331 62613 3340
rect 62572 3246 62612 3331
rect 62668 2465 62708 4684
rect 62859 4684 62860 4724
rect 62900 4684 62901 4724
rect 62859 4675 62901 4684
rect 62763 4640 62805 4649
rect 62763 4600 62764 4640
rect 62804 4600 62805 4640
rect 62763 4591 62805 4600
rect 62764 4136 62804 4591
rect 62764 4087 62804 4096
rect 62763 3380 62805 3389
rect 62763 3340 62764 3380
rect 62804 3340 62805 3380
rect 62763 3331 62805 3340
rect 62764 3246 62804 3331
rect 62667 2456 62709 2465
rect 62667 2416 62668 2456
rect 62708 2416 62709 2456
rect 62667 2407 62709 2416
rect 62667 1196 62709 1205
rect 62667 1156 62668 1196
rect 62708 1156 62709 1196
rect 62667 1147 62709 1156
rect 62668 80 62708 1147
rect 62860 80 62900 4675
rect 63052 4565 63092 5440
rect 63051 4556 63093 4565
rect 63051 4516 63052 4556
rect 63092 4516 63093 4556
rect 63051 4507 63093 4516
rect 63051 3884 63093 3893
rect 63051 3844 63052 3884
rect 63092 3844 63093 3884
rect 63051 3835 63093 3844
rect 63052 3380 63092 3835
rect 62956 3340 63092 3380
rect 62956 3044 62996 3340
rect 63148 3305 63188 5608
rect 63244 5489 63284 5608
rect 63531 5648 63573 5657
rect 63531 5608 63532 5648
rect 63572 5608 63573 5648
rect 63531 5599 63573 5608
rect 63628 5648 63668 5657
rect 63724 5648 63764 9211
rect 66124 9101 66164 9388
rect 65408 9092 65776 9101
rect 65448 9052 65490 9092
rect 65530 9052 65572 9092
rect 65612 9052 65654 9092
rect 65694 9052 65736 9092
rect 65408 9043 65776 9052
rect 66123 9092 66165 9101
rect 66123 9052 66124 9092
rect 66164 9052 66165 9092
rect 66123 9043 66165 9052
rect 64011 8840 64053 8849
rect 64011 8800 64012 8840
rect 64052 8800 64053 8840
rect 64011 8791 64053 8800
rect 64012 7916 64052 8791
rect 64971 8672 65013 8681
rect 64971 8632 64972 8672
rect 65012 8632 65013 8672
rect 64971 8623 65013 8632
rect 64168 8336 64536 8345
rect 64208 8296 64250 8336
rect 64290 8296 64332 8336
rect 64372 8296 64414 8336
rect 64454 8296 64496 8336
rect 64168 8287 64536 8296
rect 64683 8084 64725 8093
rect 64683 8044 64684 8084
rect 64724 8044 64725 8084
rect 64683 8035 64725 8044
rect 64012 7867 64052 7876
rect 64011 7328 64053 7337
rect 64011 7288 64012 7328
rect 64052 7288 64053 7328
rect 64011 7279 64053 7288
rect 64012 7244 64052 7279
rect 64012 7193 64052 7204
rect 64491 7244 64533 7253
rect 64491 7204 64492 7244
rect 64532 7204 64533 7244
rect 64491 7195 64533 7204
rect 64684 7244 64724 8035
rect 64972 7916 65012 8623
rect 66411 8168 66453 8177
rect 66411 8128 66412 8168
rect 66452 8128 66453 8168
rect 66411 8119 66453 8128
rect 64972 7867 65012 7876
rect 65259 7916 65301 7925
rect 65259 7876 65260 7916
rect 65300 7876 65301 7916
rect 65259 7867 65301 7876
rect 66220 7916 66260 7925
rect 65260 7782 65300 7867
rect 65835 7832 65877 7841
rect 65835 7792 65836 7832
rect 65876 7792 65877 7832
rect 65835 7783 65877 7792
rect 65408 7580 65776 7589
rect 65448 7540 65490 7580
rect 65530 7540 65572 7580
rect 65612 7540 65654 7580
rect 65694 7540 65736 7580
rect 65408 7531 65776 7540
rect 64684 7195 64724 7204
rect 64972 7244 65012 7253
rect 64492 7110 64532 7195
rect 64011 7076 64053 7085
rect 64011 7036 64012 7076
rect 64052 7036 64053 7076
rect 64011 7027 64053 7036
rect 64012 6404 64052 7027
rect 64972 6917 65012 7204
rect 65164 7244 65204 7253
rect 64971 6908 65013 6917
rect 64971 6868 64972 6908
rect 65012 6868 65013 6908
rect 64971 6859 65013 6868
rect 65164 6833 65204 7204
rect 64168 6824 64536 6833
rect 64208 6784 64250 6824
rect 64290 6784 64332 6824
rect 64372 6784 64414 6824
rect 64454 6784 64496 6824
rect 64168 6775 64536 6784
rect 65163 6824 65205 6833
rect 65163 6784 65164 6824
rect 65204 6784 65205 6824
rect 65163 6775 65205 6784
rect 64779 6488 64821 6497
rect 64779 6448 64780 6488
rect 64820 6448 64821 6488
rect 64779 6439 64821 6448
rect 64012 6355 64052 6364
rect 64780 6329 64820 6439
rect 64972 6404 65012 6415
rect 64972 6329 65012 6364
rect 65259 6404 65301 6413
rect 65259 6364 65260 6404
rect 65300 6364 65301 6404
rect 65259 6355 65301 6364
rect 64779 6320 64821 6329
rect 64779 6280 64780 6320
rect 64820 6280 64821 6320
rect 64779 6271 64821 6280
rect 64971 6320 65013 6329
rect 64971 6280 64972 6320
rect 65012 6280 65013 6320
rect 64971 6271 65013 6280
rect 65260 6270 65300 6355
rect 65067 6152 65109 6161
rect 65067 6112 65068 6152
rect 65108 6112 65109 6152
rect 65067 6103 65109 6112
rect 63915 5900 63957 5909
rect 63915 5860 63916 5900
rect 63956 5860 63957 5900
rect 63915 5851 63957 5860
rect 65068 5900 65108 6103
rect 65408 6068 65776 6077
rect 65448 6028 65490 6068
rect 65530 6028 65572 6068
rect 65612 6028 65654 6068
rect 65694 6028 65736 6068
rect 65408 6019 65776 6028
rect 65259 5984 65301 5993
rect 65259 5944 65260 5984
rect 65300 5944 65301 5984
rect 65259 5935 65301 5944
rect 65068 5851 65108 5860
rect 63668 5608 63764 5648
rect 63628 5599 63668 5608
rect 63243 5480 63285 5489
rect 63436 5480 63476 5489
rect 63243 5440 63244 5480
rect 63284 5440 63285 5480
rect 63243 5431 63285 5440
rect 63340 5440 63436 5480
rect 63243 4892 63285 4901
rect 63243 4852 63244 4892
rect 63284 4852 63285 4892
rect 63243 4843 63285 4852
rect 63244 4758 63284 4843
rect 63340 3893 63380 5440
rect 63436 5431 63476 5440
rect 63435 4892 63477 4901
rect 63435 4852 63436 4892
rect 63476 4852 63477 4892
rect 63435 4843 63477 4852
rect 63436 4758 63476 4843
rect 63532 4808 63572 5599
rect 63820 5564 63860 5573
rect 63532 4768 63668 4808
rect 63531 4472 63573 4481
rect 63531 4432 63532 4472
rect 63572 4432 63573 4472
rect 63531 4423 63573 4432
rect 63435 4388 63477 4397
rect 63435 4348 63436 4388
rect 63476 4348 63477 4388
rect 63435 4339 63477 4348
rect 63436 4220 63476 4339
rect 63436 4171 63476 4180
rect 63339 3884 63381 3893
rect 63339 3844 63340 3884
rect 63380 3844 63381 3884
rect 63339 3835 63381 3844
rect 63532 3632 63572 4423
rect 63628 4207 63668 4768
rect 63724 4724 63764 4733
rect 63724 4481 63764 4684
rect 63723 4472 63765 4481
rect 63723 4432 63724 4472
rect 63764 4432 63765 4472
rect 63723 4423 63765 4432
rect 63628 4167 63764 4207
rect 63627 4052 63669 4061
rect 63627 4012 63628 4052
rect 63668 4012 63669 4052
rect 63627 4003 63669 4012
rect 63628 3918 63668 4003
rect 63340 3592 63572 3632
rect 63243 3464 63285 3473
rect 63243 3424 63244 3464
rect 63284 3424 63285 3464
rect 63243 3415 63285 3424
rect 63244 3330 63284 3415
rect 63147 3296 63189 3305
rect 63147 3256 63148 3296
rect 63188 3256 63189 3296
rect 63147 3247 63189 3256
rect 63052 3212 63092 3221
rect 63052 3128 63092 3172
rect 63052 3088 63284 3128
rect 62956 3004 63092 3044
rect 63052 80 63092 3004
rect 63244 1877 63284 3088
rect 63340 2381 63380 3592
rect 63628 3464 63668 3473
rect 63724 3464 63764 4167
rect 63668 3424 63764 3464
rect 63628 3415 63668 3424
rect 63820 3380 63860 5524
rect 63916 4976 63956 5851
rect 64587 5732 64629 5741
rect 64587 5692 64588 5732
rect 64628 5692 64629 5732
rect 64587 5683 64629 5692
rect 64011 5648 64053 5657
rect 64011 5608 64012 5648
rect 64052 5608 64053 5648
rect 64011 5599 64053 5608
rect 64012 5514 64052 5599
rect 64588 5598 64628 5683
rect 64168 5312 64536 5321
rect 64208 5272 64250 5312
rect 64290 5272 64332 5312
rect 64372 5272 64414 5312
rect 64454 5272 64496 5312
rect 64168 5263 64536 5272
rect 64011 5228 64053 5237
rect 64011 5188 64012 5228
rect 64052 5188 64053 5228
rect 64011 5179 64053 5188
rect 63916 4927 63956 4936
rect 63915 3548 63957 3557
rect 63915 3508 63916 3548
rect 63956 3508 63957 3548
rect 63915 3499 63957 3508
rect 63724 3340 63860 3380
rect 63531 3296 63573 3305
rect 63724 3296 63764 3340
rect 63531 3256 63532 3296
rect 63572 3256 63573 3296
rect 63531 3247 63573 3256
rect 63628 3256 63764 3296
rect 63435 3212 63477 3221
rect 63435 3172 63436 3212
rect 63476 3172 63477 3212
rect 63435 3163 63477 3172
rect 63436 3078 63476 3163
rect 63339 2372 63381 2381
rect 63339 2332 63340 2372
rect 63380 2332 63381 2372
rect 63339 2323 63381 2332
rect 63532 2036 63572 3247
rect 63436 1996 63572 2036
rect 63243 1868 63285 1877
rect 63243 1828 63244 1868
rect 63284 1828 63285 1868
rect 63243 1819 63285 1828
rect 63243 1700 63285 1709
rect 63243 1660 63244 1700
rect 63284 1660 63285 1700
rect 63243 1651 63285 1660
rect 63244 80 63284 1651
rect 63436 80 63476 1996
rect 63628 80 63668 3256
rect 63820 3212 63860 3221
rect 63724 3172 63820 3212
rect 63724 1037 63764 3172
rect 63820 3163 63860 3172
rect 63916 3137 63956 3499
rect 64012 3464 64052 5179
rect 64779 5060 64821 5069
rect 64779 5020 64780 5060
rect 64820 5020 64821 5060
rect 64779 5011 64821 5020
rect 64300 4976 64340 4985
rect 64107 4724 64149 4733
rect 64107 4684 64108 4724
rect 64148 4684 64149 4724
rect 64107 4675 64149 4684
rect 64108 4590 64148 4675
rect 64203 4472 64245 4481
rect 64203 4432 64204 4472
rect 64244 4432 64245 4472
rect 64203 4423 64245 4432
rect 64204 4304 64244 4423
rect 64300 4397 64340 4936
rect 64395 4976 64437 4985
rect 64395 4936 64396 4976
rect 64436 4936 64437 4976
rect 64395 4927 64437 4936
rect 64587 4976 64629 4985
rect 64587 4936 64588 4976
rect 64628 4936 64629 4976
rect 64587 4927 64629 4936
rect 64396 4733 64436 4927
rect 64395 4724 64437 4733
rect 64395 4684 64396 4724
rect 64436 4684 64437 4724
rect 64395 4675 64437 4684
rect 64299 4388 64341 4397
rect 64299 4348 64300 4388
rect 64340 4348 64341 4388
rect 64299 4339 64341 4348
rect 64204 4255 64244 4264
rect 64588 4229 64628 4927
rect 64780 4892 64820 5011
rect 64780 4843 64820 4852
rect 64780 4229 64820 4314
rect 64587 4220 64629 4229
rect 64779 4220 64821 4229
rect 64587 4180 64588 4220
rect 64628 4180 64629 4220
rect 64587 4171 64629 4180
rect 64684 4180 64780 4220
rect 64820 4180 64821 4220
rect 64588 4086 64628 4171
rect 64587 3968 64629 3977
rect 64587 3928 64588 3968
rect 64628 3928 64629 3968
rect 64587 3919 64629 3928
rect 64168 3800 64536 3809
rect 64208 3760 64250 3800
rect 64290 3760 64332 3800
rect 64372 3760 64414 3800
rect 64454 3760 64496 3800
rect 64168 3751 64536 3760
rect 64396 3464 64436 3473
rect 64012 3415 64052 3424
rect 64300 3424 64396 3464
rect 64204 3212 64244 3221
rect 63915 3128 63957 3137
rect 63915 3088 63916 3128
rect 63956 3088 63957 3128
rect 63915 3079 63957 3088
rect 63915 2960 63957 2969
rect 63915 2920 63916 2960
rect 63956 2920 63957 2960
rect 63915 2911 63957 2920
rect 63819 2792 63861 2801
rect 63819 2752 63820 2792
rect 63860 2752 63861 2792
rect 63819 2743 63861 2752
rect 63723 1028 63765 1037
rect 63723 988 63724 1028
rect 63764 988 63765 1028
rect 63723 979 63765 988
rect 63820 80 63860 2743
rect 63916 2717 63956 2911
rect 63915 2708 63957 2717
rect 63915 2668 63916 2708
rect 63956 2668 63957 2708
rect 63915 2659 63957 2668
rect 64204 2540 64244 3172
rect 64300 2969 64340 3424
rect 64396 3415 64436 3424
rect 64588 3380 64628 3919
rect 64684 3893 64724 4180
rect 64779 4171 64821 4180
rect 65260 4136 65300 5935
rect 65451 5564 65493 5573
rect 65451 5524 65452 5564
rect 65492 5524 65493 5564
rect 65451 5515 65493 5524
rect 65452 5060 65492 5515
rect 65452 5011 65492 5020
rect 65408 4556 65776 4565
rect 65448 4516 65490 4556
rect 65530 4516 65572 4556
rect 65612 4516 65654 4556
rect 65694 4516 65736 4556
rect 65408 4507 65776 4516
rect 65836 4388 65876 7783
rect 66220 7673 66260 7876
rect 66219 7664 66261 7673
rect 66219 7624 66220 7664
rect 66260 7624 66261 7664
rect 66219 7615 66261 7624
rect 66219 7160 66261 7169
rect 66219 7120 66220 7160
rect 66260 7120 66261 7160
rect 66219 7111 66261 7120
rect 66220 6404 66260 7111
rect 66220 6355 66260 6364
rect 66412 6404 66452 8119
rect 66795 7244 66837 7253
rect 66795 7204 66796 7244
rect 66836 7204 66837 7244
rect 66795 7195 66837 7204
rect 66796 7110 66836 7195
rect 66603 6488 66645 6497
rect 66603 6448 66604 6488
rect 66644 6448 66645 6488
rect 66603 6439 66645 6448
rect 66412 6355 66452 6364
rect 66604 6404 66644 6439
rect 66604 6353 66644 6364
rect 66411 5732 66453 5741
rect 66411 5692 66412 5732
rect 66452 5692 66453 5732
rect 66411 5683 66453 5692
rect 66124 4976 66164 4985
rect 66028 4936 66124 4976
rect 65260 4087 65300 4096
rect 65548 4348 65876 4388
rect 65932 4724 65972 4733
rect 64779 4052 64821 4061
rect 64779 4012 64780 4052
rect 64820 4012 64821 4052
rect 64779 4003 64821 4012
rect 64780 3918 64820 4003
rect 65068 3968 65108 3977
rect 65452 3968 65492 3977
rect 64683 3884 64725 3893
rect 64683 3844 64684 3884
rect 64724 3844 64725 3884
rect 64683 3835 64725 3844
rect 64875 3884 64917 3893
rect 64875 3844 64876 3884
rect 64916 3844 64917 3884
rect 64875 3835 64917 3844
rect 64779 3800 64821 3809
rect 64779 3760 64780 3800
rect 64820 3760 64821 3800
rect 64779 3751 64821 3760
rect 64780 3632 64820 3751
rect 64492 3340 64628 3380
rect 64684 3592 64820 3632
rect 64395 3212 64437 3221
rect 64395 3172 64396 3212
rect 64436 3172 64437 3212
rect 64395 3163 64437 3172
rect 64299 2960 64341 2969
rect 64299 2920 64300 2960
rect 64340 2920 64341 2960
rect 64299 2911 64341 2920
rect 64108 2500 64244 2540
rect 64011 1280 64053 1289
rect 64011 1240 64012 1280
rect 64052 1240 64053 1280
rect 64011 1231 64053 1240
rect 64012 80 64052 1231
rect 64108 953 64148 2500
rect 64396 2213 64436 3163
rect 64395 2204 64437 2213
rect 64395 2164 64396 2204
rect 64436 2164 64437 2204
rect 64395 2155 64437 2164
rect 64492 2036 64532 3340
rect 64587 3212 64629 3221
rect 64587 3172 64588 3212
rect 64628 3172 64629 3212
rect 64587 3163 64629 3172
rect 64588 3078 64628 3163
rect 64587 2876 64629 2885
rect 64587 2836 64588 2876
rect 64628 2836 64629 2876
rect 64587 2827 64629 2836
rect 64396 1996 64532 2036
rect 64203 1616 64245 1625
rect 64203 1576 64204 1616
rect 64244 1576 64245 1616
rect 64203 1567 64245 1576
rect 64107 944 64149 953
rect 64107 904 64108 944
rect 64148 904 64149 944
rect 64107 895 64149 904
rect 64204 80 64244 1567
rect 64396 80 64436 1996
rect 64588 80 64628 2827
rect 64684 1205 64724 3592
rect 64780 3464 64820 3473
rect 64780 3305 64820 3424
rect 64779 3296 64821 3305
rect 64779 3256 64780 3296
rect 64820 3256 64821 3296
rect 64779 3247 64821 3256
rect 64876 2036 64916 3835
rect 64971 3716 65013 3725
rect 65068 3716 65108 3928
rect 64971 3676 64972 3716
rect 65012 3676 65108 3716
rect 65164 3928 65452 3968
rect 64971 3667 65013 3676
rect 65164 3632 65204 3928
rect 65452 3919 65492 3928
rect 65259 3800 65301 3809
rect 65451 3800 65493 3809
rect 65259 3760 65260 3800
rect 65300 3760 65396 3800
rect 65259 3751 65301 3760
rect 65068 3592 65204 3632
rect 65356 3632 65396 3760
rect 65451 3760 65452 3800
rect 65492 3760 65493 3800
rect 65451 3751 65493 3760
rect 64971 3548 65013 3557
rect 64971 3508 64972 3548
rect 65012 3508 65013 3548
rect 64971 3499 65013 3508
rect 64972 3414 65012 3499
rect 64971 2960 65013 2969
rect 64971 2920 64972 2960
rect 65012 2920 65013 2960
rect 64971 2911 65013 2920
rect 64780 1996 64916 2036
rect 64683 1196 64725 1205
rect 64683 1156 64684 1196
rect 64724 1156 64725 1196
rect 64683 1147 64725 1156
rect 64780 80 64820 1996
rect 64972 80 65012 2911
rect 65068 1289 65108 3592
rect 65356 3583 65396 3592
rect 65163 3464 65205 3473
rect 65163 3424 65164 3464
rect 65204 3424 65205 3464
rect 65163 3415 65205 3424
rect 65164 3330 65204 3415
rect 65452 3212 65492 3751
rect 65548 3464 65588 4348
rect 65643 4220 65685 4229
rect 65643 4180 65644 4220
rect 65684 4180 65685 4220
rect 65643 4171 65685 4180
rect 65644 4136 65684 4171
rect 65644 4085 65684 4096
rect 65835 3968 65877 3977
rect 65835 3928 65836 3968
rect 65876 3928 65877 3968
rect 65835 3919 65877 3928
rect 65836 3834 65876 3919
rect 65932 3809 65972 4684
rect 66028 4397 66068 4936
rect 66124 4927 66164 4936
rect 66316 4724 66356 4733
rect 66124 4684 66316 4724
rect 66027 4388 66069 4397
rect 66027 4348 66028 4388
rect 66068 4348 66069 4388
rect 66027 4339 66069 4348
rect 66027 4136 66069 4145
rect 66027 4096 66028 4136
rect 66068 4096 66069 4136
rect 66027 4087 66069 4096
rect 66028 4002 66068 4087
rect 65931 3800 65973 3809
rect 65931 3760 65932 3800
rect 65972 3760 65973 3800
rect 65931 3751 65973 3760
rect 66124 3632 66164 4684
rect 66316 4675 66356 4684
rect 66412 4304 66452 5683
rect 66507 5480 66549 5489
rect 66796 5480 66836 5489
rect 66507 5440 66508 5480
rect 66548 5440 66549 5480
rect 66507 5431 66549 5440
rect 66604 5440 66796 5480
rect 66508 4976 66548 5431
rect 66508 4927 66548 4936
rect 66412 4264 66548 4304
rect 66411 4136 66453 4145
rect 66411 4096 66412 4136
rect 66452 4096 66453 4136
rect 66411 4087 66453 4096
rect 66220 3977 66260 4062
rect 66412 4002 66452 4087
rect 66219 3968 66261 3977
rect 66219 3928 66220 3968
rect 66260 3928 66261 3968
rect 66219 3919 66261 3928
rect 66219 3716 66261 3725
rect 66219 3676 66220 3716
rect 66260 3676 66261 3716
rect 66219 3667 66261 3676
rect 65548 3415 65588 3424
rect 65836 3592 66164 3632
rect 65740 3221 65780 3306
rect 65260 3172 65492 3212
rect 65739 3212 65781 3221
rect 65739 3172 65740 3212
rect 65780 3172 65781 3212
rect 65260 2372 65300 3172
rect 65739 3163 65781 3172
rect 65408 3044 65776 3053
rect 65448 3004 65490 3044
rect 65530 3004 65572 3044
rect 65612 3004 65654 3044
rect 65694 3004 65736 3044
rect 65408 2995 65776 3004
rect 65355 2624 65397 2633
rect 65355 2584 65356 2624
rect 65396 2584 65397 2624
rect 65355 2575 65397 2584
rect 65164 2332 65300 2372
rect 65067 1280 65109 1289
rect 65067 1240 65068 1280
rect 65108 1240 65109 1280
rect 65067 1231 65109 1240
rect 65164 80 65204 2332
rect 65356 80 65396 2575
rect 65836 2372 65876 3592
rect 65931 3464 65973 3473
rect 65931 3424 65932 3464
rect 65972 3424 65973 3464
rect 65931 3415 65973 3424
rect 65932 3330 65972 3415
rect 66027 3212 66069 3221
rect 66027 3172 66028 3212
rect 66068 3172 66069 3212
rect 66027 3163 66069 3172
rect 66124 3212 66164 3221
rect 65931 2708 65973 2717
rect 65931 2668 65932 2708
rect 65972 2668 65973 2708
rect 65931 2659 65973 2668
rect 65548 2332 65876 2372
rect 65548 80 65588 2332
rect 65932 1448 65972 2659
rect 66028 1709 66068 3163
rect 66124 2801 66164 3172
rect 66123 2792 66165 2801
rect 66123 2752 66124 2792
rect 66164 2752 66165 2792
rect 66123 2743 66165 2752
rect 66220 2372 66260 3667
rect 66315 3548 66357 3557
rect 66315 3508 66316 3548
rect 66356 3508 66357 3548
rect 66315 3499 66357 3508
rect 66316 3464 66356 3499
rect 66316 3413 66356 3424
rect 66508 3389 66548 4264
rect 66507 3380 66549 3389
rect 66507 3340 66508 3380
rect 66548 3340 66549 3380
rect 66507 3331 66549 3340
rect 66315 3212 66357 3221
rect 66508 3212 66548 3221
rect 66315 3172 66316 3212
rect 66356 3172 66357 3212
rect 66315 3163 66357 3172
rect 66412 3172 66508 3212
rect 66124 2332 66260 2372
rect 66027 1700 66069 1709
rect 66027 1660 66028 1700
rect 66068 1660 66069 1700
rect 66027 1651 66069 1660
rect 65740 1408 65972 1448
rect 65740 80 65780 1408
rect 65931 1280 65973 1289
rect 65931 1240 65932 1280
rect 65972 1240 65973 1280
rect 65931 1231 65973 1240
rect 65932 80 65972 1231
rect 66124 80 66164 2332
rect 66316 80 66356 3163
rect 66412 1625 66452 3172
rect 66508 3163 66548 3172
rect 66507 2792 66549 2801
rect 66507 2752 66508 2792
rect 66548 2752 66549 2792
rect 66507 2743 66549 2752
rect 66411 1616 66453 1625
rect 66411 1576 66412 1616
rect 66452 1576 66453 1616
rect 66411 1567 66453 1576
rect 66508 80 66548 2743
rect 66604 2540 66644 5440
rect 66796 5431 66836 5440
rect 66892 4976 66932 9463
rect 66987 8756 67029 8765
rect 66987 8716 66988 8756
rect 67028 8716 67029 8756
rect 66987 8707 67029 8716
rect 67179 8756 67221 8765
rect 67179 8716 67180 8756
rect 67220 8716 67221 8756
rect 67179 8707 67221 8716
rect 66988 8622 67028 8707
rect 67180 8622 67220 8707
rect 67851 8000 67893 8009
rect 67851 7960 67852 8000
rect 67892 7960 67893 8000
rect 67851 7951 67893 7960
rect 67179 7916 67221 7925
rect 67179 7876 67180 7916
rect 67220 7876 67221 7916
rect 67179 7867 67221 7876
rect 67372 7916 67412 7925
rect 67180 7782 67220 7867
rect 67372 7757 67412 7876
rect 67659 7916 67701 7925
rect 67659 7876 67660 7916
rect 67700 7876 67701 7916
rect 67659 7867 67701 7876
rect 67852 7916 67892 7951
rect 67660 7782 67700 7867
rect 67852 7865 67892 7876
rect 67371 7748 67413 7757
rect 67371 7708 67372 7748
rect 67412 7708 67413 7748
rect 67371 7699 67413 7708
rect 66988 7244 67028 7253
rect 67948 7244 67988 9547
rect 70540 9428 70580 9437
rect 70059 9260 70101 9269
rect 70059 9220 70060 9260
rect 70100 9220 70101 9260
rect 70059 9211 70101 9220
rect 68715 8924 68757 8933
rect 68715 8884 68716 8924
rect 68756 8884 68757 8924
rect 68715 8875 68757 8884
rect 68716 7916 68756 8875
rect 70060 8840 70100 9211
rect 70540 9185 70580 9388
rect 70731 9428 70773 9437
rect 70731 9388 70732 9428
rect 70772 9388 70773 9428
rect 70731 9379 70773 9388
rect 70732 9294 70772 9379
rect 70539 9176 70581 9185
rect 70539 9136 70540 9176
rect 70580 9136 70581 9176
rect 70539 9127 70581 9136
rect 71211 9176 71253 9185
rect 71211 9136 71212 9176
rect 71252 9136 71253 9176
rect 71211 9127 71253 9136
rect 70060 8791 70100 8800
rect 70252 8884 70580 8924
rect 69964 8756 70004 8765
rect 69964 7925 70004 8716
rect 70155 8756 70197 8765
rect 70155 8716 70156 8756
rect 70196 8716 70197 8756
rect 70155 8707 70197 8716
rect 70156 8622 70196 8707
rect 70252 8084 70292 8884
rect 70540 8840 70580 8884
rect 70540 8791 70580 8800
rect 70923 8840 70965 8849
rect 70923 8800 70924 8840
rect 70964 8800 70965 8840
rect 70923 8791 70965 8800
rect 70060 8044 70292 8084
rect 70444 8756 70484 8765
rect 68716 7867 68756 7876
rect 68907 7916 68949 7925
rect 68907 7876 68908 7916
rect 68948 7876 68949 7916
rect 68907 7867 68949 7876
rect 69771 7916 69813 7925
rect 69771 7876 69772 7916
rect 69812 7876 69813 7916
rect 69771 7867 69813 7876
rect 69963 7916 70005 7925
rect 69963 7876 69964 7916
rect 70004 7876 70005 7916
rect 69963 7867 70005 7876
rect 68908 7782 68948 7867
rect 69772 7589 69812 7867
rect 69868 7832 69908 7841
rect 69771 7580 69813 7589
rect 69771 7540 69772 7580
rect 69812 7540 69813 7580
rect 69771 7531 69813 7540
rect 66988 7085 67028 7204
rect 67852 7204 67988 7244
rect 68043 7244 68085 7253
rect 68236 7244 68276 7255
rect 68043 7204 68044 7244
rect 68084 7204 68180 7244
rect 66987 7076 67029 7085
rect 66987 7036 66988 7076
rect 67028 7036 67029 7076
rect 66987 7027 67029 7036
rect 67083 6908 67125 6917
rect 67083 6868 67084 6908
rect 67124 6868 67125 6908
rect 67083 6859 67125 6868
rect 67084 6413 67124 6859
rect 67179 6572 67221 6581
rect 67179 6532 67180 6572
rect 67220 6532 67221 6572
rect 67179 6523 67221 6532
rect 67276 6572 67316 6581
rect 67316 6532 67604 6572
rect 67276 6523 67316 6532
rect 67083 6404 67125 6413
rect 67083 6364 67084 6404
rect 67124 6364 67125 6404
rect 67083 6355 67125 6364
rect 67180 6404 67220 6523
rect 67180 6355 67220 6364
rect 67371 6404 67413 6413
rect 67371 6364 67372 6404
rect 67412 6364 67413 6404
rect 67371 6355 67413 6364
rect 67372 6270 67412 6355
rect 67276 5732 67316 5741
rect 66987 5648 67029 5657
rect 66987 5608 66988 5648
rect 67028 5608 67029 5648
rect 66987 5599 67029 5608
rect 66988 5514 67028 5599
rect 66892 4927 66932 4936
rect 67179 4976 67221 4985
rect 67179 4936 67180 4976
rect 67220 4936 67221 4976
rect 67179 4927 67221 4936
rect 67180 4892 67220 4927
rect 67276 4892 67316 5692
rect 67468 5732 67508 6532
rect 67564 6404 67604 6532
rect 67564 6355 67604 6364
rect 67755 6404 67797 6413
rect 67755 6364 67756 6404
rect 67796 6364 67797 6404
rect 67755 6355 67797 6364
rect 67756 6270 67796 6355
rect 67852 5984 67892 7204
rect 68043 7195 68085 7204
rect 68044 7110 68084 7195
rect 67947 7076 67989 7085
rect 67947 7036 67948 7076
rect 67988 7036 67989 7076
rect 67947 7027 67989 7036
rect 67948 6236 67988 7027
rect 68043 6824 68085 6833
rect 68043 6784 68044 6824
rect 68084 6784 68085 6824
rect 68043 6775 68085 6784
rect 68044 6404 68084 6775
rect 68140 6413 68180 7204
rect 68236 7169 68276 7204
rect 68524 7244 68564 7253
rect 68715 7244 68757 7253
rect 69004 7244 69044 7253
rect 68564 7204 68660 7244
rect 68524 7195 68564 7204
rect 68235 7160 68277 7169
rect 68235 7120 68236 7160
rect 68276 7120 68277 7160
rect 68235 7111 68277 7120
rect 68236 6992 68276 7001
rect 68524 6992 68564 7001
rect 68276 6952 68372 6992
rect 68236 6943 68276 6952
rect 68044 6355 68084 6364
rect 68139 6404 68181 6413
rect 68236 6404 68276 6413
rect 68139 6364 68140 6404
rect 68180 6364 68236 6404
rect 68139 6355 68181 6364
rect 68236 6355 68276 6364
rect 68140 6236 68180 6245
rect 67948 6196 68084 6236
rect 67468 5683 67508 5692
rect 67756 5944 67892 5984
rect 67660 5480 67700 5489
rect 67468 5440 67660 5480
rect 67372 4901 67412 4986
rect 67371 4892 67413 4901
rect 67276 4852 67372 4892
rect 67412 4852 67413 4892
rect 67180 4841 67220 4852
rect 67371 4843 67413 4852
rect 66891 4808 66933 4817
rect 66891 4768 66892 4808
rect 66932 4768 66933 4808
rect 66891 4759 66933 4768
rect 66700 4724 66740 4733
rect 66700 3725 66740 4684
rect 66892 4481 66932 4759
rect 67276 4724 67316 4733
rect 67180 4684 67276 4724
rect 66891 4472 66933 4481
rect 67180 4472 67220 4684
rect 67276 4675 67316 4684
rect 66891 4432 66892 4472
rect 66932 4432 66933 4472
rect 66891 4423 66933 4432
rect 66988 4432 67220 4472
rect 66892 4220 66932 4423
rect 66892 4171 66932 4180
rect 66699 3716 66741 3725
rect 66699 3676 66700 3716
rect 66740 3676 66741 3716
rect 66699 3667 66741 3676
rect 66700 3464 66740 3475
rect 66988 3473 67028 4432
rect 67468 4313 67508 5440
rect 67660 5431 67700 5440
rect 67563 5312 67605 5321
rect 67563 5272 67564 5312
rect 67604 5272 67605 5312
rect 67563 5263 67605 5272
rect 67564 5144 67604 5263
rect 67756 5237 67796 5944
rect 67851 5816 67893 5825
rect 67851 5776 67852 5816
rect 67892 5776 67893 5816
rect 67851 5767 67893 5776
rect 67852 5648 67892 5767
rect 68044 5741 68084 6196
rect 68043 5732 68085 5741
rect 68043 5692 68044 5732
rect 68084 5692 68085 5732
rect 68043 5683 68085 5692
rect 68140 5657 68180 6196
rect 68235 6236 68277 6245
rect 68235 6196 68236 6236
rect 68276 6196 68277 6236
rect 68235 6187 68277 6196
rect 67852 5599 67892 5608
rect 68139 5648 68181 5657
rect 68139 5608 68140 5648
rect 68180 5608 68181 5648
rect 68139 5599 68181 5608
rect 67755 5228 67797 5237
rect 67755 5188 67756 5228
rect 67796 5188 67797 5228
rect 67755 5179 67797 5188
rect 67948 5144 67988 5153
rect 67564 5095 67604 5104
rect 67852 5104 67948 5144
rect 67659 5060 67701 5069
rect 67659 5020 67660 5060
rect 67700 5020 67701 5060
rect 67659 5011 67701 5020
rect 67564 4892 67604 4901
rect 67564 4649 67604 4852
rect 67563 4640 67605 4649
rect 67563 4600 67564 4640
rect 67604 4600 67605 4640
rect 67563 4591 67605 4600
rect 67083 4304 67125 4313
rect 67275 4304 67317 4313
rect 67083 4264 67084 4304
rect 67124 4264 67125 4304
rect 67083 4255 67125 4264
rect 67180 4264 67276 4304
rect 67316 4264 67317 4304
rect 67084 4220 67124 4255
rect 67084 4169 67124 4180
rect 67084 4052 67124 4061
rect 67084 3809 67124 4012
rect 67083 3800 67125 3809
rect 67083 3760 67084 3800
rect 67124 3760 67125 3800
rect 67083 3751 67125 3760
rect 66700 3389 66740 3424
rect 66987 3464 67029 3473
rect 66987 3424 66988 3464
rect 67028 3424 67029 3464
rect 66987 3415 67029 3424
rect 67084 3464 67124 3475
rect 67084 3389 67124 3424
rect 66699 3380 66741 3389
rect 66699 3340 66700 3380
rect 66740 3340 66741 3380
rect 66699 3331 66741 3340
rect 67083 3380 67125 3389
rect 67083 3340 67084 3380
rect 67124 3340 67125 3380
rect 67083 3331 67125 3340
rect 66892 3212 66932 3221
rect 66796 3172 66892 3212
rect 66796 2885 66836 3172
rect 66892 3163 66932 3172
rect 66795 2876 66837 2885
rect 66795 2836 66796 2876
rect 66836 2836 66837 2876
rect 66795 2827 66837 2836
rect 66987 2876 67029 2885
rect 66987 2836 66988 2876
rect 67028 2836 67029 2876
rect 66987 2827 67029 2836
rect 66604 2500 66740 2540
rect 66700 80 66740 2500
rect 66988 1616 67028 2827
rect 67180 2540 67220 4264
rect 67275 4255 67317 4264
rect 67467 4304 67509 4313
rect 67467 4264 67468 4304
rect 67508 4264 67509 4304
rect 67467 4255 67509 4264
rect 67564 4136 67604 4145
rect 67660 4136 67700 5011
rect 67755 4892 67797 4901
rect 67755 4852 67756 4892
rect 67796 4852 67797 4892
rect 67755 4843 67797 4852
rect 67756 4640 67796 4843
rect 67852 4724 67892 5104
rect 67948 5095 67988 5104
rect 68043 5144 68085 5153
rect 68043 5104 68044 5144
rect 68084 5104 68085 5144
rect 68043 5095 68085 5104
rect 67948 4985 67988 4987
rect 67947 4976 67989 4985
rect 67947 4936 67948 4976
rect 67988 4936 67989 4976
rect 67947 4927 67989 4936
rect 67948 4892 67988 4927
rect 67948 4843 67988 4852
rect 68044 4871 68084 5095
rect 68140 4985 68180 5000
rect 68139 4976 68181 4985
rect 68139 4936 68140 4976
rect 68180 4936 68181 4976
rect 68139 4927 68181 4936
rect 68140 4905 68180 4927
rect 68044 4831 68094 4871
rect 68140 4856 68180 4865
rect 68054 4808 68094 4831
rect 68054 4768 68180 4808
rect 67852 4684 68084 4724
rect 67756 4600 67988 4640
rect 67755 4472 67797 4481
rect 67755 4432 67756 4472
rect 67796 4432 67797 4472
rect 67755 4423 67797 4432
rect 67756 4220 67796 4423
rect 67948 4313 67988 4600
rect 67947 4304 67989 4313
rect 67947 4264 67948 4304
rect 67988 4264 67989 4304
rect 67947 4255 67989 4264
rect 67756 4171 67796 4180
rect 67948 4220 67988 4255
rect 68044 4229 68084 4684
rect 68140 4339 68180 4768
rect 68140 4229 68185 4339
rect 67948 4170 67988 4180
rect 68043 4220 68085 4229
rect 68043 4180 68044 4220
rect 68084 4180 68085 4220
rect 68043 4171 68085 4180
rect 68140 4220 68186 4229
rect 68185 4180 68186 4220
rect 68140 4171 68186 4180
rect 67604 4096 67700 4136
rect 67564 4087 67604 4096
rect 67372 3968 67412 3977
rect 67276 3212 67316 3221
rect 67276 2969 67316 3172
rect 67275 2960 67317 2969
rect 67275 2920 67276 2960
rect 67316 2920 67317 2960
rect 67275 2911 67317 2920
rect 67180 2500 67316 2540
rect 66988 1576 67124 1616
rect 66891 1364 66933 1373
rect 66891 1324 66892 1364
rect 66932 1324 66933 1364
rect 66891 1315 66933 1324
rect 66892 80 66932 1315
rect 67084 80 67124 1576
rect 67276 80 67316 2500
rect 67372 1289 67412 3928
rect 67756 3968 67796 3979
rect 68140 3977 68180 4062
rect 67756 3893 67796 3928
rect 68139 3968 68181 3977
rect 68139 3928 68140 3968
rect 68180 3928 68181 3968
rect 68139 3919 68181 3928
rect 67755 3884 67797 3893
rect 67755 3844 67756 3884
rect 67796 3844 67797 3884
rect 67755 3835 67797 3844
rect 67851 3800 67893 3809
rect 67851 3760 67852 3800
rect 67892 3760 67893 3800
rect 67851 3751 67893 3760
rect 67467 3464 67509 3473
rect 67467 3424 67468 3464
rect 67508 3424 67509 3464
rect 67467 3415 67509 3424
rect 67852 3464 67892 3751
rect 68139 3716 68181 3725
rect 68139 3676 68140 3716
rect 68180 3676 68181 3716
rect 68139 3667 68181 3676
rect 67852 3415 67892 3424
rect 67468 3330 67508 3415
rect 67660 3212 67700 3221
rect 67660 2633 67700 3172
rect 68044 3212 68084 3221
rect 68044 2717 68084 3172
rect 68043 2708 68085 2717
rect 68043 2668 68044 2708
rect 68084 2668 68085 2708
rect 68043 2659 68085 2668
rect 67659 2624 67701 2633
rect 67659 2584 67660 2624
rect 67700 2584 67701 2624
rect 67659 2575 67701 2584
rect 68140 2372 68180 3667
rect 68236 3632 68276 6187
rect 68332 5993 68372 6952
rect 68428 6952 68524 6992
rect 68620 6992 68660 7204
rect 68715 7204 68716 7244
rect 68756 7204 68757 7244
rect 68715 7195 68757 7204
rect 68908 7204 69004 7244
rect 68716 7110 68756 7195
rect 68620 6952 68756 6992
rect 68331 5984 68373 5993
rect 68331 5944 68332 5984
rect 68372 5944 68373 5984
rect 68331 5935 68373 5944
rect 68332 5741 68372 5826
rect 68331 5732 68373 5741
rect 68331 5692 68332 5732
rect 68372 5692 68373 5732
rect 68331 5683 68373 5692
rect 68331 5480 68373 5489
rect 68331 5440 68332 5480
rect 68372 5440 68373 5480
rect 68331 5431 68373 5440
rect 68332 5346 68372 5431
rect 68428 5069 68468 6952
rect 68524 6943 68564 6952
rect 68619 6656 68661 6665
rect 68619 6616 68620 6656
rect 68660 6616 68661 6656
rect 68619 6607 68661 6616
rect 68523 6404 68565 6413
rect 68523 6364 68524 6404
rect 68564 6364 68565 6404
rect 68523 6355 68565 6364
rect 68620 6404 68660 6607
rect 68620 6355 68660 6364
rect 68524 5732 68564 6355
rect 68716 6161 68756 6952
rect 68811 6572 68853 6581
rect 68811 6532 68812 6572
rect 68852 6532 68853 6572
rect 68811 6523 68853 6532
rect 68812 6404 68852 6523
rect 68812 6355 68852 6364
rect 68908 6329 68948 7204
rect 69004 7195 69044 7204
rect 69195 7244 69237 7253
rect 69195 7204 69196 7244
rect 69236 7204 69237 7244
rect 69195 7195 69237 7204
rect 69004 6992 69044 7001
rect 68907 6320 68949 6329
rect 68907 6280 68908 6320
rect 68948 6280 68949 6320
rect 68907 6271 68949 6280
rect 68908 6161 68948 6271
rect 68715 6152 68757 6161
rect 68715 6112 68716 6152
rect 68756 6112 68757 6152
rect 68715 6103 68757 6112
rect 68907 6152 68949 6161
rect 68907 6112 68908 6152
rect 68948 6112 68949 6152
rect 68907 6103 68949 6112
rect 68716 5993 68756 6103
rect 68715 5984 68757 5993
rect 68715 5944 68716 5984
rect 68756 5944 68757 5984
rect 68715 5935 68757 5944
rect 68716 5732 68756 5741
rect 68564 5692 68716 5732
rect 68524 5683 68564 5692
rect 68716 5683 68756 5692
rect 68908 5732 68948 5743
rect 68908 5657 68948 5692
rect 68812 5648 68852 5657
rect 68427 5060 68469 5069
rect 68427 5020 68428 5060
rect 68468 5020 68469 5060
rect 68427 5011 68469 5020
rect 68332 4892 68372 4903
rect 68332 4817 68372 4852
rect 68523 4892 68565 4901
rect 68523 4852 68524 4892
rect 68564 4852 68565 4892
rect 68523 4843 68565 4852
rect 68331 4808 68373 4817
rect 68331 4768 68332 4808
rect 68372 4768 68373 4808
rect 68331 4759 68373 4768
rect 68524 4758 68564 4843
rect 68812 4817 68852 5608
rect 68907 5648 68949 5657
rect 68907 5608 68908 5648
rect 68948 5608 68949 5648
rect 68907 5599 68949 5608
rect 69004 5480 69044 6952
rect 69099 6488 69141 6497
rect 69099 6448 69100 6488
rect 69140 6448 69141 6488
rect 69099 6439 69141 6448
rect 69100 6404 69140 6439
rect 69196 6404 69236 7195
rect 69675 6572 69717 6581
rect 69675 6532 69676 6572
rect 69716 6532 69717 6572
rect 69675 6523 69717 6532
rect 69292 6404 69332 6413
rect 69484 6404 69524 6413
rect 69196 6364 69292 6404
rect 69332 6364 69484 6404
rect 69100 6353 69140 6364
rect 69292 6355 69332 6364
rect 69484 6355 69524 6364
rect 69676 6404 69716 6523
rect 69676 6355 69716 6364
rect 69868 6320 69908 7792
rect 69964 7782 70004 7867
rect 70060 6908 70100 8044
rect 70347 8000 70389 8009
rect 70347 7960 70348 8000
rect 70388 7960 70389 8000
rect 70347 7951 70389 7960
rect 70155 7916 70197 7925
rect 70155 7876 70156 7916
rect 70196 7876 70197 7916
rect 70155 7867 70197 7876
rect 70348 7916 70388 7951
rect 70444 7916 70484 8716
rect 70636 8756 70676 8767
rect 70636 8681 70676 8716
rect 70828 8756 70868 8765
rect 70635 8672 70677 8681
rect 70635 8632 70636 8672
rect 70676 8632 70677 8672
rect 70635 8623 70677 8632
rect 70731 8084 70773 8093
rect 70731 8044 70732 8084
rect 70772 8044 70773 8084
rect 70731 8035 70773 8044
rect 70539 7916 70581 7925
rect 70444 7876 70540 7916
rect 70580 7876 70581 7916
rect 70156 7782 70196 7867
rect 70348 7865 70388 7876
rect 70539 7867 70581 7876
rect 70732 7916 70772 8035
rect 70828 7916 70868 8716
rect 70924 8706 70964 8791
rect 71020 8756 71060 8765
rect 71020 8597 71060 8716
rect 71019 8588 71061 8597
rect 71019 8548 71020 8588
rect 71060 8548 71061 8588
rect 71019 8539 71061 8548
rect 71115 8252 71157 8261
rect 71115 8212 71116 8252
rect 71156 8212 71157 8252
rect 71115 8203 71157 8212
rect 70923 7916 70965 7925
rect 70828 7876 70924 7916
rect 70964 7876 70965 7916
rect 70732 7867 70772 7876
rect 70923 7867 70965 7876
rect 71116 7916 71156 8203
rect 71116 7867 71156 7876
rect 70251 7832 70293 7841
rect 70251 7792 70252 7832
rect 70292 7792 70293 7832
rect 70251 7783 70293 7792
rect 70252 7698 70292 7783
rect 70540 7265 70580 7867
rect 70540 7216 70580 7225
rect 70636 7832 70676 7841
rect 70636 7160 70676 7792
rect 70924 7782 70964 7867
rect 71020 7832 71060 7841
rect 70731 7748 70773 7757
rect 70731 7708 70732 7748
rect 70772 7708 70773 7748
rect 70731 7699 70773 7708
rect 70732 7244 70772 7699
rect 70732 7195 70772 7204
rect 70540 7120 70676 7160
rect 70060 6868 70196 6908
rect 70059 6740 70101 6749
rect 70059 6700 70060 6740
rect 70100 6700 70101 6740
rect 70059 6691 70101 6700
rect 69868 6280 70004 6320
rect 69195 6236 69237 6245
rect 69195 6196 69196 6236
rect 69236 6196 69237 6236
rect 69195 6187 69237 6196
rect 69387 6236 69429 6245
rect 69387 6196 69388 6236
rect 69428 6196 69429 6236
rect 69387 6187 69429 6196
rect 69580 6236 69620 6245
rect 69620 6196 69908 6236
rect 69580 6187 69620 6196
rect 69196 6102 69236 6187
rect 69388 5825 69428 6187
rect 69387 5816 69429 5825
rect 69387 5776 69388 5816
rect 69428 5776 69429 5816
rect 69387 5767 69429 5776
rect 69772 5741 69812 5826
rect 69580 5732 69620 5741
rect 69771 5732 69813 5741
rect 69292 5648 69332 5657
rect 69332 5608 69524 5648
rect 69292 5599 69332 5608
rect 68908 5440 69044 5480
rect 69100 5480 69140 5489
rect 69387 5480 69429 5489
rect 69140 5440 69236 5480
rect 68908 4976 68948 5440
rect 69100 5431 69140 5440
rect 68908 4927 68948 4936
rect 68811 4808 68853 4817
rect 68811 4768 68812 4808
rect 68852 4768 68853 4808
rect 68811 4759 68853 4768
rect 68428 4724 68468 4733
rect 68716 4724 68756 4733
rect 68331 4304 68373 4313
rect 68331 4264 68332 4304
rect 68372 4264 68373 4304
rect 68331 4255 68373 4264
rect 68332 4220 68372 4255
rect 68332 4169 68372 4180
rect 68428 4145 68468 4684
rect 68620 4684 68716 4724
rect 68523 4556 68565 4565
rect 68523 4516 68524 4556
rect 68564 4516 68565 4556
rect 68523 4507 68565 4516
rect 68524 4220 68564 4507
rect 68524 4171 68564 4180
rect 68427 4136 68469 4145
rect 68427 4096 68428 4136
rect 68468 4096 68469 4136
rect 68427 4087 68469 4096
rect 68523 4052 68565 4061
rect 68523 4012 68524 4052
rect 68564 4012 68565 4052
rect 68523 4003 68565 4012
rect 68524 3918 68564 4003
rect 68523 3716 68565 3725
rect 68620 3716 68660 4684
rect 68716 4675 68756 4684
rect 69100 4724 69140 4733
rect 69100 4640 69140 4684
rect 68812 4600 69140 4640
rect 68715 4304 68757 4313
rect 68715 4264 68716 4304
rect 68756 4264 68757 4304
rect 68715 4255 68757 4264
rect 68716 4220 68756 4255
rect 68716 4169 68756 4180
rect 68523 3676 68524 3716
rect 68564 3676 68660 3716
rect 68523 3667 68565 3676
rect 68812 3632 68852 4600
rect 69003 4388 69045 4397
rect 69003 4348 69004 4388
rect 69044 4348 69045 4388
rect 69003 4339 69045 4348
rect 68907 4304 68949 4313
rect 68907 4264 68908 4304
rect 68948 4264 68949 4304
rect 68907 4255 68949 4264
rect 68908 4220 68948 4255
rect 69004 4254 69044 4339
rect 68908 4169 68948 4180
rect 69100 4220 69140 4229
rect 69003 4136 69045 4145
rect 69003 4096 69004 4136
rect 69044 4096 69045 4136
rect 69003 4087 69045 4096
rect 68236 3592 68468 3632
rect 68236 3464 68276 3473
rect 68428 3464 68468 3592
rect 68716 3592 68852 3632
rect 68620 3464 68660 3473
rect 68428 3424 68620 3464
rect 68236 2969 68276 3424
rect 68620 3415 68660 3424
rect 68427 3212 68469 3221
rect 68427 3172 68428 3212
rect 68468 3172 68469 3212
rect 68427 3163 68469 3172
rect 68428 3078 68468 3163
rect 68235 2960 68277 2969
rect 68235 2920 68236 2960
rect 68276 2920 68277 2960
rect 68235 2911 68277 2920
rect 68716 2372 68756 3592
rect 69004 3464 69044 4087
rect 69100 4061 69140 4180
rect 69099 4052 69141 4061
rect 69099 4012 69100 4052
rect 69140 4012 69141 4052
rect 69099 4003 69141 4012
rect 69004 3415 69044 3424
rect 69196 3380 69236 5440
rect 69387 5440 69388 5480
rect 69428 5440 69429 5480
rect 69387 5431 69429 5440
rect 69291 5396 69333 5405
rect 69291 5356 69292 5396
rect 69332 5356 69333 5396
rect 69291 5347 69333 5356
rect 69292 4976 69332 5347
rect 69292 4927 69332 4936
rect 69291 4724 69333 4733
rect 69291 4684 69292 4724
rect 69332 4684 69333 4724
rect 69291 4675 69333 4684
rect 69292 4313 69332 4675
rect 69291 4304 69333 4313
rect 69291 4264 69292 4304
rect 69332 4264 69333 4304
rect 69291 4255 69333 4264
rect 69100 3340 69236 3380
rect 69292 3968 69332 3977
rect 68812 3212 68852 3221
rect 68812 2801 68852 3172
rect 68811 2792 68853 2801
rect 68811 2752 68812 2792
rect 68852 2752 68853 2792
rect 68811 2743 68853 2752
rect 68811 2624 68853 2633
rect 68811 2584 68812 2624
rect 68852 2584 68853 2624
rect 68811 2575 68853 2584
rect 67852 2332 68180 2372
rect 68428 2332 68756 2372
rect 67371 1280 67413 1289
rect 67371 1240 67372 1280
rect 67412 1240 67413 1280
rect 67371 1231 67413 1240
rect 67467 1112 67509 1121
rect 67467 1072 67468 1112
rect 67508 1072 67509 1112
rect 67467 1063 67509 1072
rect 67468 80 67508 1063
rect 67659 860 67701 869
rect 67659 820 67660 860
rect 67700 820 67701 860
rect 67659 811 67701 820
rect 67660 80 67700 811
rect 67852 80 67892 2332
rect 68235 1868 68277 1877
rect 68235 1828 68236 1868
rect 68276 1828 68277 1868
rect 68235 1819 68277 1828
rect 68043 1616 68085 1625
rect 68043 1576 68044 1616
rect 68084 1576 68085 1616
rect 68043 1567 68085 1576
rect 68044 80 68084 1567
rect 68236 80 68276 1819
rect 68428 80 68468 2332
rect 68619 1196 68661 1205
rect 68619 1156 68620 1196
rect 68660 1156 68661 1196
rect 68619 1147 68661 1156
rect 68620 80 68660 1147
rect 68812 80 68852 2575
rect 69100 2540 69140 3340
rect 69004 2500 69140 2540
rect 69196 3212 69236 3221
rect 69004 80 69044 2500
rect 69196 1373 69236 3172
rect 69195 1364 69237 1373
rect 69195 1324 69196 1364
rect 69236 1324 69237 1364
rect 69195 1315 69237 1324
rect 69195 1028 69237 1037
rect 69195 988 69196 1028
rect 69236 988 69237 1028
rect 69195 979 69237 988
rect 69196 80 69236 979
rect 69292 869 69332 3928
rect 69388 3632 69428 5431
rect 69484 4304 69524 5608
rect 69580 5573 69620 5692
rect 69676 5692 69772 5732
rect 69812 5692 69813 5732
rect 69579 5564 69621 5573
rect 69579 5524 69580 5564
rect 69620 5524 69621 5564
rect 69579 5515 69621 5524
rect 69580 5153 69620 5515
rect 69579 5144 69621 5153
rect 69579 5104 69580 5144
rect 69620 5104 69621 5144
rect 69676 5144 69716 5692
rect 69771 5683 69813 5692
rect 69772 5480 69812 5489
rect 69772 5321 69812 5440
rect 69771 5312 69813 5321
rect 69771 5272 69772 5312
rect 69812 5272 69813 5312
rect 69771 5263 69813 5272
rect 69676 5104 69812 5144
rect 69579 5095 69621 5104
rect 69675 4976 69717 4985
rect 69675 4936 69676 4976
rect 69716 4936 69717 4976
rect 69675 4927 69717 4936
rect 69580 4892 69620 4901
rect 69580 4481 69620 4852
rect 69676 4842 69716 4927
rect 69772 4901 69812 5104
rect 69771 4892 69813 4901
rect 69771 4852 69772 4892
rect 69812 4852 69813 4892
rect 69771 4843 69813 4852
rect 69868 4724 69908 6196
rect 69964 5909 70004 6280
rect 69963 5900 70005 5909
rect 69963 5860 69964 5900
rect 70004 5860 70005 5900
rect 69963 5851 70005 5860
rect 69963 5480 70005 5489
rect 69963 5440 69964 5480
rect 70004 5440 70005 5480
rect 69963 5431 70005 5440
rect 69964 5346 70004 5431
rect 70060 5405 70100 6691
rect 70156 6245 70196 6868
rect 70155 6236 70197 6245
rect 70155 6196 70156 6236
rect 70196 6196 70197 6236
rect 70155 6187 70197 6196
rect 70155 5816 70197 5825
rect 70155 5776 70156 5816
rect 70196 5776 70197 5816
rect 70540 5816 70580 7120
rect 70636 6992 70676 7001
rect 70636 6077 70676 6952
rect 71020 6572 71060 7792
rect 70828 6532 71060 6572
rect 70635 6068 70677 6077
rect 70635 6028 70636 6068
rect 70676 6028 70677 6068
rect 70635 6019 70677 6028
rect 70540 5776 70676 5816
rect 70155 5767 70197 5776
rect 70156 5661 70196 5767
rect 70540 5648 70580 5657
rect 70156 5612 70196 5621
rect 70444 5608 70540 5648
rect 70348 5480 70388 5489
rect 70252 5440 70348 5480
rect 70059 5396 70101 5405
rect 70059 5356 70060 5396
rect 70100 5356 70101 5396
rect 70059 5347 70101 5356
rect 70156 4901 70196 4986
rect 69772 4684 69908 4724
rect 69964 4892 70004 4901
rect 69579 4472 69621 4481
rect 69579 4432 69580 4472
rect 69620 4432 69621 4472
rect 69579 4423 69621 4432
rect 69484 4264 69620 4304
rect 69483 4136 69525 4145
rect 69483 4096 69484 4136
rect 69524 4096 69525 4136
rect 69483 4087 69525 4096
rect 69484 4002 69524 4087
rect 69580 4061 69620 4264
rect 69579 4052 69621 4061
rect 69579 4012 69580 4052
rect 69620 4012 69621 4052
rect 69579 4003 69621 4012
rect 69676 3968 69716 3977
rect 69388 3592 69524 3632
rect 69387 3464 69429 3473
rect 69387 3424 69388 3464
rect 69428 3424 69429 3464
rect 69387 3415 69429 3424
rect 69388 3330 69428 3415
rect 69484 2540 69524 3592
rect 69580 3212 69620 3221
rect 69580 2885 69620 3172
rect 69579 2876 69621 2885
rect 69579 2836 69580 2876
rect 69620 2836 69621 2876
rect 69579 2827 69621 2836
rect 69484 2500 69620 2540
rect 69387 1280 69429 1289
rect 69387 1240 69388 1280
rect 69428 1240 69429 1280
rect 69387 1231 69429 1240
rect 69291 860 69333 869
rect 69291 820 69292 860
rect 69332 820 69333 860
rect 69291 811 69333 820
rect 69388 80 69428 1231
rect 69580 80 69620 2500
rect 69676 1877 69716 3928
rect 69772 3464 69812 4684
rect 69964 4649 70004 4852
rect 70155 4892 70197 4901
rect 70155 4852 70156 4892
rect 70196 4852 70197 4892
rect 70155 4843 70197 4852
rect 70060 4724 70100 4733
rect 70100 4684 70196 4724
rect 70060 4675 70100 4684
rect 69963 4640 70005 4649
rect 69963 4600 69964 4640
rect 70004 4600 70005 4640
rect 69963 4591 70005 4600
rect 69867 4556 69909 4565
rect 69867 4516 69868 4556
rect 69908 4516 69909 4556
rect 69867 4507 69909 4516
rect 70059 4556 70101 4565
rect 70059 4516 70060 4556
rect 70100 4516 70101 4556
rect 70059 4507 70101 4516
rect 69868 4136 69908 4507
rect 70060 4313 70100 4507
rect 70059 4304 70101 4313
rect 70059 4264 70060 4304
rect 70100 4264 70101 4304
rect 70059 4255 70101 4264
rect 70060 4220 70100 4255
rect 70060 4169 70100 4180
rect 69868 4087 69908 4096
rect 70059 3800 70101 3809
rect 70059 3760 70060 3800
rect 70100 3760 70101 3800
rect 70059 3751 70101 3760
rect 70060 3464 70100 3751
rect 70156 3641 70196 4684
rect 70252 4388 70292 5440
rect 70348 5431 70388 5440
rect 70347 5060 70389 5069
rect 70347 5020 70348 5060
rect 70388 5020 70389 5060
rect 70347 5011 70389 5020
rect 70348 4892 70388 5011
rect 70348 4843 70388 4852
rect 70444 4817 70484 5608
rect 70540 5599 70580 5608
rect 70539 5480 70581 5489
rect 70539 5440 70540 5480
rect 70580 5440 70581 5480
rect 70539 5431 70581 5440
rect 70540 5144 70580 5431
rect 70636 5405 70676 5776
rect 70732 5480 70772 5489
rect 70635 5396 70677 5405
rect 70635 5356 70636 5396
rect 70676 5356 70677 5396
rect 70635 5347 70677 5356
rect 70540 5095 70580 5104
rect 70540 4901 70580 4986
rect 70539 4892 70581 4901
rect 70732 4892 70772 5440
rect 70828 5405 70868 6532
rect 71020 6404 71060 6415
rect 71020 6329 71060 6364
rect 71019 6320 71061 6329
rect 71019 6280 71020 6320
rect 71060 6280 71061 6320
rect 71019 6271 71061 6280
rect 71212 6068 71252 9127
rect 71404 6413 71444 9976
rect 71596 9428 71636 10228
rect 72171 9764 72213 9773
rect 72171 9724 72172 9764
rect 72212 9724 72213 9764
rect 72171 9715 72213 9724
rect 72075 9596 72117 9605
rect 72075 9556 72076 9596
rect 72116 9556 72117 9596
rect 72075 9547 72117 9556
rect 72076 9462 72116 9547
rect 71596 9353 71636 9388
rect 71787 9428 71829 9437
rect 71787 9388 71788 9428
rect 71828 9388 71829 9428
rect 71787 9379 71829 9388
rect 71980 9428 72020 9437
rect 71595 9344 71637 9353
rect 71595 9304 71596 9344
rect 71636 9304 71637 9344
rect 71595 9295 71637 9304
rect 71692 9344 71732 9353
rect 71692 8084 71732 9304
rect 71788 9294 71828 9379
rect 71980 9353 72020 9388
rect 72172 9428 72212 9715
rect 71979 9344 72021 9353
rect 71979 9304 71980 9344
rect 72020 9304 72021 9344
rect 71979 9295 72021 9304
rect 71980 8840 72020 9295
rect 72172 9017 72212 9388
rect 72171 9008 72213 9017
rect 72171 8968 72172 9008
rect 72212 8968 72213 9008
rect 72171 8959 72213 8968
rect 71980 8800 72308 8840
rect 72075 8168 72117 8177
rect 72075 8128 72076 8168
rect 72116 8128 72117 8168
rect 72075 8119 72117 8128
rect 71596 8044 71732 8084
rect 71499 7412 71541 7421
rect 71499 7372 71500 7412
rect 71540 7372 71541 7412
rect 71499 7363 71541 7372
rect 71500 6665 71540 7363
rect 71499 6656 71541 6665
rect 71499 6616 71500 6656
rect 71540 6616 71541 6656
rect 71499 6607 71541 6616
rect 71403 6404 71445 6413
rect 71403 6364 71404 6404
rect 71444 6364 71445 6404
rect 71403 6355 71445 6364
rect 71307 6320 71349 6329
rect 71307 6280 71308 6320
rect 71348 6280 71349 6320
rect 71307 6271 71349 6280
rect 71308 6186 71348 6271
rect 71500 6236 71540 6607
rect 71500 6187 71540 6196
rect 71212 6028 71444 6068
rect 71307 5732 71349 5741
rect 71307 5692 71308 5732
rect 71348 5692 71349 5732
rect 71307 5683 71349 5692
rect 70924 5648 70964 5657
rect 70924 5489 70964 5608
rect 71308 5598 71348 5683
rect 70923 5480 70965 5489
rect 70923 5440 70924 5480
rect 70964 5440 70965 5480
rect 70923 5431 70965 5440
rect 70827 5396 70869 5405
rect 70827 5356 70828 5396
rect 70868 5356 70869 5396
rect 70827 5347 70869 5356
rect 70923 4976 70965 4985
rect 70923 4936 70924 4976
rect 70964 4936 70965 4976
rect 70923 4927 70965 4936
rect 70539 4852 70540 4892
rect 70580 4852 70581 4892
rect 70539 4843 70581 4852
rect 70636 4852 70772 4892
rect 70827 4892 70869 4901
rect 70827 4852 70828 4892
rect 70868 4852 70869 4892
rect 70443 4808 70485 4817
rect 70443 4768 70444 4808
rect 70484 4768 70485 4808
rect 70443 4759 70485 4768
rect 70636 4388 70676 4852
rect 70827 4843 70869 4852
rect 70731 4724 70773 4733
rect 70731 4684 70732 4724
rect 70772 4684 70773 4724
rect 70731 4675 70773 4684
rect 70732 4590 70772 4675
rect 70252 4348 70388 4388
rect 70636 4348 70772 4388
rect 70251 4220 70293 4229
rect 70251 4180 70252 4220
rect 70292 4180 70293 4220
rect 70251 4171 70293 4180
rect 70252 4086 70292 4171
rect 70252 3968 70292 3977
rect 70155 3632 70197 3641
rect 70155 3592 70156 3632
rect 70196 3592 70197 3632
rect 70155 3583 70197 3592
rect 70252 3557 70292 3928
rect 70251 3548 70293 3557
rect 70251 3508 70252 3548
rect 70292 3508 70293 3548
rect 70251 3499 70293 3508
rect 70156 3464 70196 3473
rect 70060 3424 70156 3464
rect 69772 3415 69812 3424
rect 70156 3415 70196 3424
rect 70348 3380 70388 4348
rect 70444 4229 70484 4314
rect 70443 4220 70485 4229
rect 70443 4180 70444 4220
rect 70484 4180 70485 4220
rect 70443 4171 70485 4180
rect 70636 4220 70676 4229
rect 70636 4061 70676 4180
rect 70443 4052 70485 4061
rect 70443 4012 70444 4052
rect 70484 4012 70485 4052
rect 70443 4003 70485 4012
rect 70635 4052 70677 4061
rect 70635 4012 70636 4052
rect 70676 4012 70677 4052
rect 70635 4003 70677 4012
rect 70444 3918 70484 4003
rect 70635 3884 70677 3893
rect 70635 3844 70636 3884
rect 70676 3844 70677 3884
rect 70635 3835 70677 3844
rect 70636 3632 70676 3835
rect 70252 3340 70388 3380
rect 70444 3592 70676 3632
rect 69964 3212 70004 3221
rect 69771 2372 69813 2381
rect 69771 2332 69772 2372
rect 69812 2332 69813 2372
rect 69771 2323 69813 2332
rect 69675 1868 69717 1877
rect 69675 1828 69676 1868
rect 69716 1828 69717 1868
rect 69675 1819 69717 1828
rect 69772 80 69812 2323
rect 69964 1121 70004 3172
rect 70252 2540 70292 3340
rect 70156 2500 70292 2540
rect 70348 3212 70388 3221
rect 69963 1112 70005 1121
rect 69963 1072 69964 1112
rect 70004 1072 70005 1112
rect 69963 1063 70005 1072
rect 69963 944 70005 953
rect 69963 904 69964 944
rect 70004 904 70005 944
rect 69963 895 70005 904
rect 69964 80 70004 895
rect 70156 80 70196 2500
rect 70348 1625 70388 3172
rect 70444 2381 70484 3592
rect 70550 3451 70590 3460
rect 70550 3305 70590 3411
rect 70732 3380 70772 4348
rect 70828 4229 70868 4843
rect 70924 4842 70964 4927
rect 71115 4892 71157 4901
rect 71115 4881 71116 4892
rect 71020 4852 71116 4881
rect 71156 4852 71157 4892
rect 71020 4843 71157 4852
rect 71307 4892 71349 4901
rect 71307 4852 71308 4892
rect 71348 4852 71349 4892
rect 71307 4843 71349 4852
rect 71020 4841 71156 4843
rect 70923 4724 70965 4733
rect 70923 4684 70924 4724
rect 70964 4684 70965 4724
rect 70923 4675 70965 4684
rect 70924 4388 70964 4675
rect 71020 4397 71060 4841
rect 71116 4758 71156 4841
rect 71308 4758 71348 4843
rect 71211 4724 71253 4733
rect 71211 4684 71212 4724
rect 71252 4684 71253 4724
rect 71404 4724 71444 6028
rect 71499 5984 71541 5993
rect 71499 5944 71500 5984
rect 71540 5944 71541 5984
rect 71499 5935 71541 5944
rect 71500 5732 71540 5935
rect 71500 5683 71540 5692
rect 71499 5396 71541 5405
rect 71499 5356 71500 5396
rect 71540 5356 71541 5396
rect 71499 5347 71541 5356
rect 71500 4892 71540 5347
rect 71596 5237 71636 8044
rect 72076 8000 72116 8119
rect 71884 7960 72116 8000
rect 71691 7916 71733 7925
rect 71691 7876 71692 7916
rect 71732 7876 71733 7916
rect 71691 7867 71733 7876
rect 71884 7916 71924 7960
rect 71884 7867 71924 7876
rect 72076 7916 72116 7960
rect 72076 7867 72116 7876
rect 72268 7916 72308 8800
rect 72268 7867 72308 7876
rect 71692 7782 71732 7867
rect 71883 7412 71925 7421
rect 71883 7372 71884 7412
rect 71924 7372 71925 7412
rect 71883 7363 71925 7372
rect 71787 6656 71829 6665
rect 71787 6616 71788 6656
rect 71828 6616 71829 6656
rect 71787 6607 71829 6616
rect 71788 6413 71828 6607
rect 71787 6404 71829 6413
rect 71787 6364 71788 6404
rect 71828 6364 71829 6404
rect 71787 6355 71829 6364
rect 71788 6270 71828 6355
rect 71691 5900 71733 5909
rect 71691 5860 71692 5900
rect 71732 5860 71733 5900
rect 71691 5851 71733 5860
rect 71692 5657 71732 5851
rect 71691 5648 71733 5657
rect 71691 5608 71692 5648
rect 71732 5608 71733 5648
rect 71691 5599 71733 5608
rect 71595 5228 71637 5237
rect 71595 5188 71596 5228
rect 71636 5188 71637 5228
rect 71595 5179 71637 5188
rect 71692 5069 71732 5154
rect 71691 5060 71733 5069
rect 71691 5020 71692 5060
rect 71732 5020 71733 5060
rect 71691 5011 71733 5020
rect 71691 4892 71733 4901
rect 71540 4852 71636 4892
rect 71500 4843 71540 4852
rect 71404 4684 71540 4724
rect 71211 4675 71253 4684
rect 71212 4590 71252 4675
rect 70924 4339 70964 4348
rect 71019 4388 71061 4397
rect 71019 4348 71020 4388
rect 71060 4348 71061 4388
rect 71019 4339 71061 4348
rect 70827 4220 70869 4229
rect 70827 4180 70828 4220
rect 70868 4180 70869 4220
rect 70827 4171 70869 4180
rect 71020 4220 71060 4229
rect 70828 4086 70868 4171
rect 71020 3977 71060 4180
rect 71211 4220 71253 4229
rect 71211 4180 71212 4220
rect 71252 4180 71253 4220
rect 71211 4171 71253 4180
rect 71404 4220 71444 4229
rect 71212 4086 71252 4171
rect 71307 4136 71349 4145
rect 71307 4096 71308 4136
rect 71348 4096 71349 4136
rect 71307 4087 71349 4096
rect 71308 4002 71348 4087
rect 71404 4061 71444 4180
rect 71403 4052 71445 4061
rect 71403 4012 71404 4052
rect 71444 4012 71445 4052
rect 71403 4003 71445 4012
rect 71019 3968 71061 3977
rect 71019 3928 71020 3968
rect 71060 3928 71061 3968
rect 71019 3919 71061 3928
rect 71404 3809 71444 4003
rect 71403 3800 71445 3809
rect 71403 3760 71404 3800
rect 71444 3760 71445 3800
rect 71403 3751 71445 3760
rect 70923 3632 70965 3641
rect 70923 3592 70924 3632
rect 70964 3592 70965 3632
rect 70923 3583 70965 3592
rect 70924 3464 70964 3583
rect 70924 3415 70964 3424
rect 71308 3464 71348 3473
rect 71500 3464 71540 4684
rect 71596 4649 71636 4852
rect 71691 4852 71692 4892
rect 71732 4852 71828 4892
rect 71691 4843 71733 4852
rect 71692 4758 71732 4843
rect 71595 4640 71637 4649
rect 71595 4600 71596 4640
rect 71636 4600 71637 4640
rect 71595 4591 71637 4600
rect 71595 4472 71637 4481
rect 71595 4432 71596 4472
rect 71636 4432 71637 4472
rect 71595 4423 71637 4432
rect 71596 4220 71636 4423
rect 71788 4229 71828 4852
rect 71596 4171 71636 4180
rect 71787 4220 71829 4229
rect 71787 4180 71788 4220
rect 71828 4180 71829 4220
rect 71787 4171 71829 4180
rect 71788 4086 71828 4171
rect 71787 3968 71829 3977
rect 71787 3928 71788 3968
rect 71828 3928 71829 3968
rect 71787 3919 71829 3928
rect 71788 3834 71828 3919
rect 71787 3632 71829 3641
rect 71787 3592 71788 3632
rect 71828 3592 71829 3632
rect 71787 3583 71829 3592
rect 71692 3464 71732 3473
rect 71500 3424 71692 3464
rect 70636 3340 70772 3380
rect 70549 3296 70591 3305
rect 70549 3256 70550 3296
rect 70590 3256 70591 3296
rect 70549 3247 70591 3256
rect 70636 2540 70676 3340
rect 71308 3305 71348 3424
rect 71692 3415 71732 3424
rect 71788 3305 71828 3583
rect 71884 3389 71924 7363
rect 72364 7253 72404 10900
rect 82924 10891 82964 10900
rect 83115 10940 83157 10949
rect 83115 10900 83116 10940
rect 83156 10900 83157 10940
rect 83115 10891 83157 10900
rect 83116 10806 83156 10891
rect 80528 10604 80896 10613
rect 80568 10564 80610 10604
rect 80650 10564 80692 10604
rect 80732 10564 80774 10604
rect 80814 10564 80856 10604
rect 80528 10555 80896 10564
rect 95648 10604 96016 10613
rect 95688 10564 95730 10604
rect 95770 10564 95812 10604
rect 95852 10564 95894 10604
rect 95934 10564 95976 10604
rect 95648 10555 96016 10564
rect 73803 10520 73845 10529
rect 73803 10480 73804 10520
rect 73844 10480 73845 10520
rect 73803 10471 73845 10480
rect 73995 10520 74037 10529
rect 73995 10480 73996 10520
rect 74036 10480 74037 10520
rect 73995 10471 74037 10480
rect 77067 10520 77109 10529
rect 77067 10480 77068 10520
rect 77108 10480 77109 10520
rect 77067 10471 77109 10480
rect 78027 10520 78069 10529
rect 78027 10480 78028 10520
rect 78068 10480 78069 10520
rect 78027 10471 78069 10480
rect 82827 10520 82869 10529
rect 82827 10480 82828 10520
rect 82868 10480 82869 10520
rect 82827 10471 82869 10480
rect 84075 10520 84117 10529
rect 84075 10480 84076 10520
rect 84116 10480 84117 10520
rect 84075 10471 84117 10480
rect 88299 10520 88341 10529
rect 88299 10480 88300 10520
rect 88340 10480 88341 10520
rect 88299 10471 88341 10480
rect 92811 10520 92853 10529
rect 92811 10480 92812 10520
rect 92852 10480 92853 10520
rect 92811 10471 92853 10480
rect 73131 10352 73173 10361
rect 73131 10312 73132 10352
rect 73172 10312 73173 10352
rect 73131 10303 73173 10312
rect 72940 10268 72980 10277
rect 72940 10025 72980 10228
rect 73132 10268 73172 10303
rect 73132 10109 73172 10228
rect 73323 10268 73365 10277
rect 73323 10228 73324 10268
rect 73364 10228 73365 10268
rect 73323 10219 73365 10228
rect 73515 10268 73557 10277
rect 73515 10228 73516 10268
rect 73556 10228 73557 10268
rect 73515 10219 73557 10228
rect 73804 10268 73844 10471
rect 73996 10268 74036 10471
rect 76491 10352 76533 10361
rect 76491 10312 76492 10352
rect 76532 10312 76533 10352
rect 76491 10303 76533 10312
rect 73804 10219 73844 10228
rect 73900 10228 73996 10268
rect 73324 10134 73364 10219
rect 73516 10134 73556 10219
rect 73131 10100 73173 10109
rect 73131 10060 73132 10100
rect 73172 10060 73173 10100
rect 73131 10051 73173 10060
rect 72939 10016 72981 10025
rect 72939 9976 72940 10016
rect 72980 9976 72981 10016
rect 72939 9967 72981 9976
rect 73036 10016 73076 10025
rect 72940 9353 72980 9967
rect 73036 9521 73076 9976
rect 73227 10016 73269 10025
rect 73227 9976 73228 10016
rect 73268 9976 73269 10016
rect 73227 9967 73269 9976
rect 73228 9521 73268 9967
rect 73803 9680 73845 9689
rect 73803 9640 73804 9680
rect 73844 9640 73845 9680
rect 73803 9631 73845 9640
rect 73804 9546 73844 9631
rect 73035 9512 73077 9521
rect 73227 9512 73269 9521
rect 73035 9472 73036 9512
rect 73076 9472 73077 9512
rect 73035 9463 73077 9472
rect 73132 9472 73228 9512
rect 73268 9472 73269 9512
rect 73132 9428 73172 9472
rect 73227 9463 73269 9472
rect 73707 9512 73749 9521
rect 73707 9472 73708 9512
rect 73748 9472 73749 9512
rect 73707 9463 73749 9472
rect 72939 9344 72981 9353
rect 72939 9304 72940 9344
rect 72980 9304 72981 9344
rect 72939 9295 72981 9304
rect 72939 9008 72981 9017
rect 72939 8968 72940 9008
rect 72980 8968 72981 9008
rect 72939 8959 72981 8968
rect 72555 8168 72597 8177
rect 72555 8128 72556 8168
rect 72596 8128 72597 8168
rect 72555 8119 72597 8128
rect 72556 8034 72596 8119
rect 72747 7916 72789 7925
rect 72747 7876 72748 7916
rect 72788 7876 72789 7916
rect 72747 7867 72789 7876
rect 72748 7782 72788 7867
rect 72844 7748 72884 7757
rect 72844 7505 72884 7708
rect 72843 7496 72885 7505
rect 72843 7456 72844 7496
rect 72884 7456 72885 7496
rect 72843 7447 72885 7456
rect 72363 7244 72405 7253
rect 72363 7204 72364 7244
rect 72404 7204 72405 7244
rect 72363 7195 72405 7204
rect 71979 6656 72021 6665
rect 71979 6616 71980 6656
rect 72020 6616 72021 6656
rect 71979 6607 72021 6616
rect 71980 6572 72020 6607
rect 71980 6521 72020 6532
rect 71980 6404 72020 6413
rect 71980 6245 72020 6364
rect 72364 6245 72404 7195
rect 72844 6917 72884 7447
rect 72843 6908 72885 6917
rect 72843 6868 72844 6908
rect 72884 6868 72885 6908
rect 72843 6859 72885 6868
rect 72651 6656 72693 6665
rect 72651 6616 72652 6656
rect 72692 6616 72693 6656
rect 72651 6607 72693 6616
rect 72652 6404 72692 6607
rect 72652 6355 72692 6364
rect 72844 6404 72884 6859
rect 72844 6355 72884 6364
rect 72748 6320 72788 6329
rect 71979 6236 72021 6245
rect 71979 6196 71980 6236
rect 72020 6196 72021 6236
rect 71979 6187 72021 6196
rect 72363 6236 72405 6245
rect 72363 6196 72364 6236
rect 72404 6196 72405 6236
rect 72363 6187 72405 6196
rect 72748 5993 72788 6280
rect 72940 6245 72980 8959
rect 73035 8924 73077 8933
rect 73035 8884 73036 8924
rect 73076 8884 73077 8924
rect 73035 8875 73077 8884
rect 73036 6329 73076 8875
rect 73132 8756 73172 9388
rect 73324 9428 73364 9437
rect 73228 9344 73268 9353
rect 73228 8924 73268 9304
rect 73324 9101 73364 9388
rect 73708 9428 73748 9463
rect 73708 9377 73748 9388
rect 73900 9428 73940 10228
rect 73996 10219 74036 10228
rect 74284 10268 74324 10277
rect 74187 9680 74229 9689
rect 74187 9640 74188 9680
rect 74228 9640 74229 9680
rect 74187 9631 74229 9640
rect 73900 9379 73940 9388
rect 73323 9092 73365 9101
rect 73323 9052 73324 9092
rect 73364 9052 73365 9092
rect 73323 9043 73365 9052
rect 73420 9052 73844 9092
rect 73420 8924 73460 9052
rect 73228 8884 73460 8924
rect 73707 8924 73749 8933
rect 73707 8884 73708 8924
rect 73748 8884 73749 8924
rect 73707 8875 73749 8884
rect 73228 8756 73268 8765
rect 73132 8716 73228 8756
rect 73228 8707 73268 8716
rect 73420 8756 73460 8765
rect 73324 8504 73364 8513
rect 73324 8345 73364 8464
rect 73420 8429 73460 8716
rect 73419 8420 73461 8429
rect 73419 8380 73420 8420
rect 73460 8380 73461 8420
rect 73419 8371 73461 8380
rect 73323 8336 73365 8345
rect 73323 8296 73324 8336
rect 73364 8296 73365 8336
rect 73323 8287 73365 8296
rect 73420 7673 73460 8371
rect 73419 7664 73461 7673
rect 73419 7624 73420 7664
rect 73460 7624 73461 7664
rect 73419 7615 73461 7624
rect 73228 6404 73268 6413
rect 73035 6320 73077 6329
rect 73035 6280 73036 6320
rect 73076 6280 73077 6320
rect 73035 6271 73077 6280
rect 72939 6236 72981 6245
rect 72939 6196 72940 6236
rect 72980 6196 72981 6236
rect 72939 6187 72981 6196
rect 73228 6077 73268 6364
rect 73420 6404 73460 6413
rect 73460 6364 73652 6404
rect 73420 6355 73460 6364
rect 73515 6236 73557 6245
rect 73515 6196 73516 6236
rect 73556 6196 73557 6236
rect 73515 6187 73557 6196
rect 73227 6068 73269 6077
rect 73227 6028 73228 6068
rect 73268 6028 73269 6068
rect 73227 6019 73269 6028
rect 73516 5993 73556 6187
rect 72747 5984 72789 5993
rect 72747 5944 72748 5984
rect 72788 5944 72789 5984
rect 72747 5935 72789 5944
rect 73515 5984 73557 5993
rect 73515 5944 73516 5984
rect 73556 5944 73557 5984
rect 73515 5935 73557 5944
rect 72075 5900 72117 5909
rect 72075 5860 72076 5900
rect 72116 5860 72117 5900
rect 72075 5851 72117 5860
rect 72076 5766 72116 5851
rect 73612 5741 73652 6364
rect 71980 5732 72020 5741
rect 71980 5405 72020 5692
rect 72172 5732 72212 5741
rect 71979 5396 72021 5405
rect 71979 5356 71980 5396
rect 72020 5356 72021 5396
rect 71979 5347 72021 5356
rect 72172 5069 72212 5692
rect 72364 5732 72404 5741
rect 72364 5489 72404 5692
rect 72556 5732 72596 5741
rect 72748 5732 72788 5741
rect 72940 5732 72980 5741
rect 72596 5692 72692 5732
rect 72556 5683 72596 5692
rect 72363 5480 72405 5489
rect 72363 5440 72364 5480
rect 72404 5440 72405 5480
rect 72363 5431 72405 5440
rect 72555 5480 72597 5489
rect 72555 5440 72556 5480
rect 72596 5440 72597 5480
rect 72555 5431 72597 5440
rect 72556 5346 72596 5431
rect 72652 5405 72692 5692
rect 72748 5573 72788 5692
rect 72844 5692 72940 5732
rect 72747 5564 72789 5573
rect 72747 5524 72748 5564
rect 72788 5524 72789 5564
rect 72747 5515 72789 5524
rect 72651 5396 72693 5405
rect 72651 5356 72652 5396
rect 72692 5356 72693 5396
rect 72651 5347 72693 5356
rect 72651 5228 72693 5237
rect 72651 5188 72652 5228
rect 72692 5188 72693 5228
rect 72651 5179 72693 5188
rect 72171 5060 72213 5069
rect 72171 5020 72172 5060
rect 72212 5020 72213 5060
rect 72171 5011 72213 5020
rect 72555 5060 72597 5069
rect 72555 5020 72556 5060
rect 72596 5020 72597 5060
rect 72555 5011 72597 5020
rect 72363 4976 72405 4985
rect 72363 4936 72364 4976
rect 72404 4936 72405 4976
rect 72363 4927 72405 4936
rect 71980 4892 72020 4901
rect 71980 4481 72020 4852
rect 72172 4892 72212 4901
rect 72075 4808 72117 4817
rect 72075 4768 72076 4808
rect 72116 4768 72117 4808
rect 72075 4759 72117 4768
rect 72076 4674 72116 4759
rect 72172 4733 72212 4852
rect 72364 4892 72404 4927
rect 72171 4724 72213 4733
rect 72171 4684 72172 4724
rect 72212 4684 72213 4724
rect 72171 4675 72213 4684
rect 72075 4556 72117 4565
rect 72075 4516 72076 4556
rect 72116 4516 72117 4556
rect 72075 4507 72117 4516
rect 71979 4472 72021 4481
rect 71979 4432 71980 4472
rect 72020 4432 72021 4472
rect 71979 4423 72021 4432
rect 71980 4220 72020 4229
rect 72076 4220 72116 4507
rect 72267 4388 72309 4397
rect 72267 4348 72268 4388
rect 72308 4348 72309 4388
rect 72267 4339 72309 4348
rect 72020 4180 72116 4220
rect 72171 4220 72213 4229
rect 72171 4180 72172 4220
rect 72212 4180 72213 4220
rect 71980 4171 72020 4180
rect 72171 4171 72213 4180
rect 72172 4086 72212 4171
rect 72171 3968 72213 3977
rect 72171 3928 72172 3968
rect 72212 3928 72213 3968
rect 72171 3919 72213 3928
rect 72172 3834 72212 3919
rect 71979 3800 72021 3809
rect 71979 3760 71980 3800
rect 72020 3760 72021 3800
rect 71979 3751 72021 3760
rect 71883 3380 71925 3389
rect 71883 3340 71884 3380
rect 71924 3340 71925 3380
rect 71883 3331 71925 3340
rect 71307 3296 71349 3305
rect 71307 3256 71308 3296
rect 71348 3256 71349 3296
rect 71307 3247 71349 3256
rect 71787 3296 71829 3305
rect 71787 3256 71788 3296
rect 71828 3256 71829 3296
rect 71787 3247 71829 3256
rect 70540 2500 70676 2540
rect 70732 3212 70772 3221
rect 70443 2372 70485 2381
rect 70443 2332 70444 2372
rect 70484 2332 70485 2372
rect 70443 2323 70485 2332
rect 70347 1616 70389 1625
rect 70347 1576 70348 1616
rect 70388 1576 70389 1616
rect 70347 1567 70389 1576
rect 70347 524 70389 533
rect 70347 484 70348 524
rect 70388 484 70389 524
rect 70347 475 70389 484
rect 70348 80 70388 475
rect 70540 80 70580 2500
rect 70732 1205 70772 3172
rect 71116 3212 71156 3221
rect 71116 2633 71156 3172
rect 71211 3212 71253 3221
rect 71211 3172 71212 3212
rect 71252 3172 71253 3212
rect 71211 3163 71253 3172
rect 71500 3212 71540 3221
rect 71115 2624 71157 2633
rect 71115 2584 71116 2624
rect 71156 2584 71157 2624
rect 71115 2575 71157 2584
rect 70923 2036 70965 2045
rect 70923 1996 70924 2036
rect 70964 1996 70965 2036
rect 70923 1987 70965 1996
rect 70827 1616 70869 1625
rect 70827 1576 70828 1616
rect 70868 1576 70869 1616
rect 70827 1567 70869 1576
rect 70731 1196 70773 1205
rect 70731 1156 70732 1196
rect 70772 1156 70773 1196
rect 70731 1147 70773 1156
rect 70828 1028 70868 1567
rect 70732 988 70868 1028
rect 70732 80 70772 988
rect 70924 80 70964 1987
rect 71212 1616 71252 3163
rect 71307 1700 71349 1709
rect 71307 1660 71308 1700
rect 71348 1660 71349 1700
rect 71307 1651 71349 1660
rect 71116 1576 71252 1616
rect 71116 80 71156 1576
rect 71308 80 71348 1651
rect 71500 1037 71540 3172
rect 71884 3212 71924 3221
rect 71595 2624 71637 2633
rect 71595 2584 71596 2624
rect 71636 2584 71637 2624
rect 71595 2575 71637 2584
rect 71499 1028 71541 1037
rect 71499 988 71500 1028
rect 71540 988 71541 1028
rect 71499 979 71541 988
rect 71596 860 71636 2575
rect 71691 1532 71733 1541
rect 71691 1492 71692 1532
rect 71732 1492 71733 1532
rect 71691 1483 71733 1492
rect 71500 820 71636 860
rect 71500 80 71540 820
rect 71692 80 71732 1483
rect 71884 1289 71924 3172
rect 71883 1280 71925 1289
rect 71883 1240 71884 1280
rect 71924 1240 71925 1280
rect 71883 1231 71925 1240
rect 71980 1112 72020 3751
rect 72075 3548 72117 3557
rect 72075 3508 72076 3548
rect 72116 3508 72117 3548
rect 72075 3499 72117 3508
rect 72076 3464 72116 3499
rect 72268 3464 72308 4339
rect 72364 4229 72404 4852
rect 72556 4892 72596 5011
rect 72460 4724 72500 4733
rect 72363 4220 72405 4229
rect 72363 4180 72364 4220
rect 72404 4180 72405 4220
rect 72363 4171 72405 4180
rect 72076 3413 72116 3424
rect 72172 3424 72308 3464
rect 72364 3968 72404 3977
rect 72075 2708 72117 2717
rect 72075 2668 72076 2708
rect 72116 2668 72117 2708
rect 72075 2659 72117 2668
rect 71884 1072 72020 1112
rect 71884 80 71924 1072
rect 72076 80 72116 2659
rect 72172 776 72212 3424
rect 72268 3212 72308 3221
rect 72268 953 72308 3172
rect 72364 2540 72404 3928
rect 72460 3884 72500 4684
rect 72556 4565 72596 4852
rect 72555 4556 72597 4565
rect 72555 4516 72556 4556
rect 72596 4516 72597 4556
rect 72555 4507 72597 4516
rect 72652 4388 72692 5179
rect 72844 5069 72884 5692
rect 72940 5683 72980 5692
rect 73419 5732 73461 5741
rect 73419 5692 73420 5732
rect 73460 5692 73461 5732
rect 73419 5683 73461 5692
rect 73611 5732 73653 5741
rect 73611 5692 73612 5732
rect 73652 5692 73653 5732
rect 73611 5683 73653 5692
rect 73227 5648 73269 5657
rect 73227 5608 73228 5648
rect 73268 5608 73269 5648
rect 73227 5599 73269 5608
rect 72939 5480 72981 5489
rect 72939 5440 72940 5480
rect 72980 5440 72981 5480
rect 72939 5431 72981 5440
rect 72940 5346 72980 5431
rect 73228 5405 73268 5599
rect 73420 5598 73460 5683
rect 73515 5648 73557 5657
rect 73515 5608 73516 5648
rect 73556 5608 73557 5648
rect 73515 5599 73557 5608
rect 73516 5514 73556 5599
rect 73612 5598 73652 5683
rect 73227 5396 73269 5405
rect 73227 5356 73228 5396
rect 73268 5356 73269 5396
rect 73227 5347 73269 5356
rect 73324 5144 73364 5153
rect 73515 5144 73557 5153
rect 73364 5104 73516 5144
rect 73556 5104 73557 5144
rect 73324 5095 73364 5104
rect 73515 5095 73557 5104
rect 72843 5060 72885 5069
rect 72843 5020 72844 5060
rect 72884 5020 72885 5060
rect 72843 5011 72885 5020
rect 72940 4901 72980 4986
rect 73131 4976 73173 4985
rect 73127 4936 73132 4976
rect 73172 4936 73173 4976
rect 73127 4927 73173 4936
rect 73708 4976 73748 8875
rect 73804 6077 73844 9052
rect 74188 8084 74228 9631
rect 74284 9521 74324 10228
rect 74475 10268 74517 10277
rect 74475 10228 74476 10268
rect 74516 10228 74517 10268
rect 74475 10219 74517 10228
rect 76492 10268 76532 10303
rect 74476 10134 74516 10219
rect 76492 10217 76532 10228
rect 76684 10268 76724 10277
rect 76876 10268 76916 10277
rect 76724 10228 76876 10268
rect 74379 10100 74421 10109
rect 74379 10060 74380 10100
rect 74420 10060 74421 10100
rect 74379 10051 74421 10060
rect 74380 9966 74420 10051
rect 76588 10016 76628 10025
rect 74283 9512 74325 9521
rect 74283 9472 74284 9512
rect 74324 9472 74325 9512
rect 74283 9463 74325 9472
rect 75435 9176 75477 9185
rect 75435 9136 75436 9176
rect 75476 9136 75477 9176
rect 75435 9127 75477 9136
rect 74667 9008 74709 9017
rect 74667 8968 74668 9008
rect 74708 8968 74709 9008
rect 74667 8959 74709 8968
rect 74668 8840 74708 8959
rect 74668 8791 74708 8800
rect 75051 8840 75093 8849
rect 75051 8800 75052 8840
rect 75092 8800 75093 8840
rect 75051 8791 75093 8800
rect 74572 8756 74612 8765
rect 74572 8597 74612 8716
rect 74763 8756 74805 8765
rect 74763 8716 74764 8756
rect 74804 8716 74805 8756
rect 74763 8707 74805 8716
rect 74956 8756 74996 8765
rect 74571 8588 74613 8597
rect 74571 8548 74572 8588
rect 74612 8548 74613 8588
rect 74571 8539 74613 8548
rect 74379 8336 74421 8345
rect 74379 8296 74380 8336
rect 74420 8296 74421 8336
rect 74379 8287 74421 8296
rect 74380 8093 74420 8287
rect 74379 8084 74421 8093
rect 74764 8084 74804 8707
rect 74956 8261 74996 8716
rect 75052 8706 75092 8791
rect 75148 8765 75188 8850
rect 75436 8840 75476 9127
rect 76588 8933 76628 9976
rect 76684 9269 76724 10228
rect 76876 10219 76916 10228
rect 77068 10268 77108 10471
rect 77643 10436 77685 10445
rect 77643 10396 77644 10436
rect 77684 10396 77685 10436
rect 77643 10387 77685 10396
rect 77068 10219 77108 10228
rect 77259 10268 77301 10277
rect 77259 10228 77260 10268
rect 77300 10228 77301 10268
rect 77259 10219 77301 10228
rect 77452 10268 77492 10277
rect 77260 10134 77300 10219
rect 77452 10193 77492 10228
rect 77644 10268 77684 10387
rect 77451 10184 77493 10193
rect 77451 10144 77452 10184
rect 77492 10144 77493 10184
rect 77451 10135 77493 10144
rect 76972 10016 77012 10025
rect 76876 9976 76972 10016
rect 76683 9260 76725 9269
rect 76683 9220 76684 9260
rect 76724 9220 76725 9260
rect 76683 9211 76725 9220
rect 76587 8924 76629 8933
rect 76587 8884 76588 8924
rect 76628 8884 76629 8924
rect 76587 8875 76629 8884
rect 75436 8791 75476 8800
rect 76011 8840 76053 8849
rect 76011 8800 76012 8840
rect 76052 8800 76053 8840
rect 76011 8791 76053 8800
rect 75147 8756 75189 8765
rect 75147 8716 75148 8756
rect 75188 8716 75189 8756
rect 75147 8707 75189 8716
rect 75340 8756 75380 8767
rect 75340 8681 75380 8716
rect 75531 8756 75573 8765
rect 75531 8716 75532 8756
rect 75572 8716 75573 8756
rect 75531 8707 75573 8716
rect 75916 8756 75956 8765
rect 75339 8672 75381 8681
rect 75339 8632 75340 8672
rect 75380 8632 75381 8672
rect 75339 8623 75381 8632
rect 75147 8504 75189 8513
rect 75147 8464 75148 8504
rect 75188 8464 75189 8504
rect 75147 8455 75189 8464
rect 74955 8252 74997 8261
rect 74955 8212 74956 8252
rect 74996 8212 74997 8252
rect 74955 8203 74997 8212
rect 75051 8168 75093 8177
rect 75051 8128 75052 8168
rect 75092 8128 75093 8168
rect 75051 8119 75093 8128
rect 74188 8044 74324 8084
rect 73995 8000 74037 8009
rect 73995 7960 73996 8000
rect 74036 7960 74037 8000
rect 73995 7951 74037 7960
rect 73996 7916 74036 7951
rect 73996 7757 74036 7876
rect 74187 7916 74229 7925
rect 74187 7876 74188 7916
rect 74228 7876 74229 7916
rect 74187 7867 74229 7876
rect 74092 7832 74132 7841
rect 73995 7748 74037 7757
rect 73995 7708 73996 7748
rect 74036 7708 74037 7748
rect 73995 7699 74037 7708
rect 74092 6824 74132 7792
rect 74188 7782 74228 7867
rect 74284 7412 74324 8044
rect 74379 8044 74380 8084
rect 74420 8044 74421 8084
rect 74379 8035 74421 8044
rect 74572 8044 74804 8084
rect 74380 7916 74420 8035
rect 74572 7925 74612 8044
rect 75052 8034 75092 8119
rect 74380 7867 74420 7876
rect 74571 7916 74613 7925
rect 74571 7876 74572 7916
rect 74612 7876 74613 7916
rect 74571 7867 74613 7876
rect 74860 7916 74900 7925
rect 74900 7876 74996 7916
rect 74860 7867 74900 7876
rect 74476 7832 74516 7841
rect 74476 7421 74516 7792
rect 74572 7782 74612 7867
rect 74764 7748 74804 7757
rect 74764 7505 74804 7708
rect 74859 7580 74901 7589
rect 74859 7540 74860 7580
rect 74900 7540 74901 7580
rect 74859 7531 74901 7540
rect 74763 7496 74805 7505
rect 74763 7456 74764 7496
rect 74804 7456 74805 7496
rect 74763 7447 74805 7456
rect 74188 7372 74324 7412
rect 74475 7412 74517 7421
rect 74475 7372 74476 7412
rect 74516 7372 74517 7412
rect 74188 7001 74228 7372
rect 74475 7363 74517 7372
rect 74284 7244 74324 7253
rect 74476 7244 74516 7253
rect 74284 7085 74324 7204
rect 74380 7204 74476 7244
rect 74283 7076 74325 7085
rect 74283 7036 74284 7076
rect 74324 7036 74325 7076
rect 74283 7027 74325 7036
rect 74187 6992 74229 7001
rect 74187 6952 74188 6992
rect 74228 6952 74229 6992
rect 74187 6943 74229 6952
rect 74284 6833 74324 7027
rect 73900 6784 74132 6824
rect 74283 6824 74325 6833
rect 74283 6784 74284 6824
rect 74324 6784 74325 6824
rect 73900 6245 73940 6784
rect 74283 6775 74325 6784
rect 73995 6656 74037 6665
rect 73995 6616 73996 6656
rect 74036 6616 74037 6656
rect 73995 6607 74037 6616
rect 74187 6656 74229 6665
rect 74187 6616 74188 6656
rect 74228 6616 74229 6656
rect 74187 6607 74229 6616
rect 73996 6404 74036 6607
rect 74091 6572 74133 6581
rect 74091 6532 74092 6572
rect 74132 6532 74133 6572
rect 74091 6523 74133 6532
rect 74092 6413 74132 6523
rect 74188 6522 74228 6607
rect 74380 6488 74420 7204
rect 74476 7195 74516 7204
rect 74860 7244 74900 7531
rect 74956 7421 74996 7876
rect 75051 7580 75093 7589
rect 75051 7540 75052 7580
rect 75092 7540 75093 7580
rect 75051 7531 75093 7540
rect 74955 7412 74997 7421
rect 74955 7372 74956 7412
rect 74996 7372 74997 7412
rect 74955 7363 74997 7372
rect 74860 7195 74900 7204
rect 75052 7244 75092 7531
rect 75052 7195 75092 7204
rect 74564 7160 74606 7169
rect 74564 7120 74565 7160
rect 74605 7120 74612 7160
rect 74564 7111 74612 7120
rect 74475 6992 74517 7001
rect 74475 6952 74476 6992
rect 74516 6952 74517 6992
rect 74475 6943 74517 6952
rect 74476 6858 74516 6943
rect 74572 6656 74612 7111
rect 74956 6992 74996 7001
rect 74996 6952 75092 6992
rect 74956 6943 74996 6952
rect 74955 6824 74997 6833
rect 74955 6784 74956 6824
rect 74996 6784 74997 6824
rect 74955 6775 74997 6784
rect 74572 6616 74708 6656
rect 74373 6448 74420 6488
rect 73899 6236 73941 6245
rect 73899 6196 73900 6236
rect 73940 6196 73941 6236
rect 73899 6187 73941 6196
rect 73996 6077 74036 6364
rect 74091 6404 74133 6413
rect 74091 6364 74092 6404
rect 74132 6364 74133 6404
rect 74091 6355 74133 6364
rect 74188 6404 74228 6413
rect 74188 6320 74228 6364
rect 74373 6393 74413 6448
rect 74572 6413 74612 6498
rect 74668 6497 74708 6616
rect 74667 6488 74709 6497
rect 74667 6448 74668 6488
rect 74708 6448 74709 6488
rect 74667 6439 74709 6448
rect 74571 6404 74613 6413
rect 74571 6364 74572 6404
rect 74612 6364 74613 6404
rect 74571 6355 74613 6364
rect 74764 6404 74804 6413
rect 74373 6329 74413 6353
rect 74373 6320 74421 6329
rect 74188 6280 74380 6320
rect 74420 6280 74421 6320
rect 73803 6068 73845 6077
rect 73803 6028 73804 6068
rect 73844 6028 73845 6068
rect 73803 6019 73845 6028
rect 73995 6068 74037 6077
rect 73995 6028 73996 6068
rect 74036 6028 74037 6068
rect 73995 6019 74037 6028
rect 73899 5984 73941 5993
rect 73899 5944 73900 5984
rect 73940 5944 73941 5984
rect 73899 5935 73941 5944
rect 73900 5816 73940 5935
rect 73804 5776 73940 5816
rect 73804 5732 73844 5776
rect 73804 5683 73844 5692
rect 73995 5732 74037 5741
rect 73995 5692 73996 5732
rect 74036 5692 74132 5732
rect 73995 5683 74037 5692
rect 73996 5598 74036 5683
rect 74092 5564 74132 5692
rect 74188 5564 74228 6280
rect 74373 6271 74421 6280
rect 74667 6320 74709 6329
rect 74764 6320 74804 6364
rect 74956 6404 74996 6775
rect 74956 6355 74996 6364
rect 74667 6280 74668 6320
rect 74708 6280 74804 6320
rect 74667 6271 74709 6280
rect 74373 6163 74413 6271
rect 74476 6236 74516 6245
rect 74860 6236 74900 6245
rect 74516 6196 74612 6236
rect 74476 6187 74516 6196
rect 74283 5816 74325 5825
rect 74283 5776 74284 5816
rect 74324 5776 74325 5816
rect 74283 5767 74325 5776
rect 74284 5732 74324 5767
rect 74476 5741 74516 5826
rect 74284 5681 74324 5692
rect 74475 5732 74517 5741
rect 74475 5692 74476 5732
rect 74516 5692 74517 5732
rect 74475 5683 74517 5692
rect 74475 5564 74517 5573
rect 74092 5524 74324 5564
rect 73996 5480 74036 5489
rect 73899 5312 73941 5321
rect 73899 5272 73900 5312
rect 73940 5272 73941 5312
rect 73899 5263 73941 5272
rect 73900 4976 73940 5263
rect 73996 5153 74036 5440
rect 74187 5396 74229 5405
rect 74187 5356 74188 5396
rect 74228 5356 74229 5396
rect 74187 5347 74229 5356
rect 73995 5144 74037 5153
rect 73995 5104 73996 5144
rect 74036 5104 74037 5144
rect 73995 5095 74037 5104
rect 74188 4985 74228 5347
rect 74187 4976 74229 4985
rect 73900 4936 74036 4976
rect 73708 4927 73748 4936
rect 73127 4905 73167 4927
rect 72939 4892 72981 4901
rect 72751 4881 72791 4890
rect 72939 4852 72940 4892
rect 72980 4852 72981 4892
rect 72939 4843 72981 4852
rect 73127 4846 73167 4865
rect 73324 4892 73364 4903
rect 72751 4808 72791 4841
rect 73324 4817 73364 4852
rect 73611 4892 73653 4901
rect 73611 4852 73612 4892
rect 73652 4852 73653 4892
rect 73611 4843 73653 4852
rect 72748 4768 72791 4808
rect 73323 4808 73365 4817
rect 73323 4768 73324 4808
rect 73364 4768 73365 4808
rect 72748 4649 72788 4768
rect 73323 4759 73365 4768
rect 72843 4724 72885 4733
rect 72843 4684 72844 4724
rect 72884 4684 72885 4724
rect 72843 4675 72885 4684
rect 73516 4724 73556 4733
rect 72747 4640 72789 4649
rect 72747 4600 72748 4640
rect 72788 4600 72789 4640
rect 72747 4591 72789 4600
rect 72844 4590 72884 4675
rect 72939 4556 72981 4565
rect 72939 4516 72940 4556
rect 72980 4516 72981 4556
rect 72939 4507 72981 4516
rect 72844 4388 72884 4397
rect 72652 4348 72844 4388
rect 72844 4339 72884 4348
rect 72747 4220 72789 4229
rect 72747 4180 72748 4220
rect 72788 4180 72789 4220
rect 72747 4171 72789 4180
rect 72940 4220 72980 4507
rect 73227 4472 73269 4481
rect 73227 4432 73228 4472
rect 73268 4432 73269 4472
rect 73227 4423 73269 4432
rect 72940 4171 72980 4180
rect 73132 4220 73172 4231
rect 72555 4136 72597 4145
rect 72555 4096 72556 4136
rect 72596 4096 72597 4136
rect 72555 4087 72597 4096
rect 72556 4002 72596 4087
rect 72748 4086 72788 4171
rect 73132 4145 73172 4180
rect 73131 4136 73173 4145
rect 73131 4096 73132 4136
rect 73172 4096 73173 4136
rect 73131 4087 73173 4096
rect 72460 3844 72596 3884
rect 72460 3464 72500 3473
rect 72460 3305 72500 3424
rect 72556 3389 72596 3844
rect 73131 3632 73173 3641
rect 73131 3592 73132 3632
rect 73172 3592 73173 3632
rect 73131 3583 73173 3592
rect 72844 3464 72884 3473
rect 72555 3380 72597 3389
rect 72555 3340 72556 3380
rect 72596 3340 72597 3380
rect 72555 3331 72597 3340
rect 72844 3305 72884 3424
rect 73132 3305 73172 3583
rect 73228 3464 73268 4423
rect 73516 4397 73556 4684
rect 73515 4388 73557 4397
rect 73515 4348 73516 4388
rect 73556 4348 73557 4388
rect 73515 4339 73557 4348
rect 73324 4229 73364 4314
rect 73323 4220 73365 4229
rect 73323 4180 73324 4220
rect 73364 4180 73365 4220
rect 73323 4171 73365 4180
rect 73516 4220 73556 4229
rect 73516 4061 73556 4180
rect 73515 4052 73557 4061
rect 73515 4012 73516 4052
rect 73556 4012 73557 4052
rect 73515 4003 73557 4012
rect 73228 3415 73268 3424
rect 73324 3968 73364 3977
rect 72459 3296 72501 3305
rect 72459 3256 72460 3296
rect 72500 3256 72501 3296
rect 72459 3247 72501 3256
rect 72843 3296 72885 3305
rect 72843 3256 72844 3296
rect 72884 3256 72885 3296
rect 72843 3247 72885 3256
rect 73131 3296 73173 3305
rect 73131 3256 73132 3296
rect 73172 3256 73173 3296
rect 73131 3247 73173 3256
rect 72652 3212 72692 3221
rect 72364 2500 72596 2540
rect 72459 2120 72501 2129
rect 72459 2080 72460 2120
rect 72500 2080 72501 2120
rect 72459 2071 72501 2080
rect 72267 944 72309 953
rect 72267 904 72268 944
rect 72308 904 72309 944
rect 72267 895 72309 904
rect 72172 736 72308 776
rect 72268 80 72308 736
rect 72460 80 72500 2071
rect 72556 2045 72596 2500
rect 72555 2036 72597 2045
rect 72555 1996 72556 2036
rect 72596 1996 72597 2036
rect 72555 1987 72597 1996
rect 72652 533 72692 3172
rect 73036 3212 73076 3221
rect 72747 3128 72789 3137
rect 72747 3088 72748 3128
rect 72788 3088 72789 3128
rect 72747 3079 72789 3088
rect 72651 524 72693 533
rect 72651 484 72652 524
rect 72692 484 72693 524
rect 72651 475 72693 484
rect 72748 356 72788 3079
rect 72843 1784 72885 1793
rect 72843 1744 72844 1784
rect 72884 1744 72885 1784
rect 72843 1735 72885 1744
rect 72652 316 72788 356
rect 72652 80 72692 316
rect 72844 80 72884 1735
rect 73036 1625 73076 3172
rect 73324 1877 73364 3928
rect 73515 3632 73557 3641
rect 73515 3592 73516 3632
rect 73556 3592 73557 3632
rect 73515 3583 73557 3592
rect 73419 3212 73461 3221
rect 73419 3172 73420 3212
rect 73460 3172 73461 3212
rect 73419 3163 73461 3172
rect 73420 3078 73460 3163
rect 73516 2540 73556 3583
rect 73612 3464 73652 4843
rect 73899 4724 73941 4733
rect 73899 4684 73900 4724
rect 73940 4684 73941 4724
rect 73899 4675 73941 4684
rect 73707 4556 73749 4565
rect 73707 4516 73708 4556
rect 73748 4516 73749 4556
rect 73707 4507 73749 4516
rect 73708 4220 73748 4507
rect 73708 4171 73748 4180
rect 73900 4145 73940 4675
rect 73899 4136 73941 4145
rect 73899 4096 73900 4136
rect 73940 4096 73941 4136
rect 73899 4087 73941 4096
rect 73708 3968 73748 3977
rect 73708 3557 73748 3928
rect 73900 3968 73940 3977
rect 73900 3809 73940 3928
rect 73899 3800 73941 3809
rect 73899 3760 73900 3800
rect 73940 3760 73941 3800
rect 73899 3751 73941 3760
rect 73707 3548 73749 3557
rect 73707 3508 73708 3548
rect 73748 3508 73749 3548
rect 73707 3499 73749 3508
rect 73612 3415 73652 3424
rect 73996 3464 74036 4936
rect 74187 4936 74188 4976
rect 74228 4936 74229 4976
rect 74187 4927 74229 4936
rect 74188 4892 74228 4927
rect 74284 4892 74324 5524
rect 74475 5524 74476 5564
rect 74516 5524 74517 5564
rect 74475 5515 74517 5524
rect 74476 5430 74516 5515
rect 74475 5312 74517 5321
rect 74475 5272 74476 5312
rect 74516 5272 74517 5312
rect 74475 5263 74517 5272
rect 74380 4892 74420 4901
rect 74284 4852 74380 4892
rect 74188 4841 74228 4852
rect 74380 4843 74420 4852
rect 74284 4724 74324 4733
rect 74188 4684 74284 4724
rect 74091 4640 74133 4649
rect 74091 4600 74092 4640
rect 74132 4600 74133 4640
rect 74091 4591 74133 4600
rect 74092 4136 74132 4591
rect 74092 4087 74132 4096
rect 74188 3473 74228 4684
rect 74284 4675 74324 4684
rect 74476 4313 74516 5263
rect 74475 4304 74517 4313
rect 74475 4264 74476 4304
rect 74516 4264 74517 4304
rect 74475 4255 74517 4264
rect 74379 4136 74421 4145
rect 74379 4096 74380 4136
rect 74420 4096 74421 4136
rect 74379 4087 74421 4096
rect 74476 4136 74516 4145
rect 74572 4136 74612 6196
rect 74764 6196 74860 6236
rect 74667 5732 74709 5741
rect 74667 5692 74668 5732
rect 74708 5692 74709 5732
rect 74667 5683 74709 5692
rect 74668 4892 74708 5683
rect 74668 4843 74708 4852
rect 74667 4304 74709 4313
rect 74667 4264 74668 4304
rect 74708 4264 74709 4304
rect 74667 4255 74709 4264
rect 74668 4220 74708 4255
rect 74668 4169 74708 4180
rect 74516 4096 74612 4136
rect 74476 4087 74516 4096
rect 74284 3968 74324 3977
rect 73996 3415 74036 3424
rect 74187 3464 74229 3473
rect 74187 3424 74188 3464
rect 74228 3424 74229 3464
rect 74187 3415 74229 3424
rect 73420 2500 73556 2540
rect 73804 3212 73844 3221
rect 73323 1868 73365 1877
rect 73323 1828 73324 1868
rect 73364 1828 73365 1868
rect 73323 1819 73365 1828
rect 73035 1616 73077 1625
rect 73035 1576 73036 1616
rect 73076 1576 73077 1616
rect 73035 1567 73077 1576
rect 73227 1280 73269 1289
rect 73227 1240 73228 1280
rect 73268 1240 73269 1280
rect 73227 1231 73269 1240
rect 73035 1196 73077 1205
rect 73035 1156 73036 1196
rect 73076 1156 73077 1196
rect 73035 1147 73077 1156
rect 73036 80 73076 1147
rect 73228 80 73268 1231
rect 73420 80 73460 2500
rect 73804 1709 73844 3172
rect 74188 3212 74228 3221
rect 74188 2633 74228 3172
rect 74187 2624 74229 2633
rect 74187 2584 74188 2624
rect 74228 2584 74229 2624
rect 74187 2575 74229 2584
rect 74284 2129 74324 3928
rect 74380 3464 74420 4087
rect 74380 3415 74420 3424
rect 74764 3464 74804 6196
rect 74860 6187 74900 6196
rect 74955 6236 74997 6245
rect 74955 6196 74956 6236
rect 74996 6196 74997 6236
rect 74955 6187 74997 6196
rect 74956 6068 74996 6187
rect 74860 6028 74996 6068
rect 74860 5648 74900 6028
rect 75052 5900 75092 6952
rect 75148 6917 75188 8455
rect 75243 8168 75285 8177
rect 75243 8128 75244 8168
rect 75284 8128 75285 8168
rect 75243 8119 75285 8128
rect 75244 7916 75284 8119
rect 75244 7867 75284 7876
rect 75436 7916 75476 7925
rect 75532 7916 75572 8707
rect 75916 8177 75956 8716
rect 75915 8168 75957 8177
rect 75915 8128 75916 8168
rect 75956 8128 75957 8168
rect 75915 8119 75957 8128
rect 75724 7916 75764 7925
rect 75476 7876 75724 7916
rect 75243 7664 75285 7673
rect 75243 7624 75244 7664
rect 75284 7624 75285 7664
rect 75243 7615 75285 7624
rect 75244 7244 75284 7615
rect 75436 7589 75476 7876
rect 75724 7867 75764 7876
rect 75916 7916 75956 7927
rect 75916 7841 75956 7876
rect 75820 7832 75860 7841
rect 75820 7673 75860 7792
rect 75915 7832 75957 7841
rect 75915 7792 75916 7832
rect 75956 7792 75957 7832
rect 75915 7783 75957 7792
rect 75819 7664 75861 7673
rect 75819 7624 75820 7664
rect 75860 7624 75861 7664
rect 75819 7615 75861 7624
rect 75435 7580 75477 7589
rect 75435 7540 75436 7580
rect 75476 7540 75477 7580
rect 75435 7531 75477 7540
rect 75244 7169 75284 7204
rect 75436 7244 75476 7531
rect 76012 7496 76052 8791
rect 76108 8756 76148 8765
rect 76684 8756 76724 9211
rect 76876 8924 76916 9976
rect 76972 9967 77012 9976
rect 77355 10016 77397 10025
rect 77355 9976 77356 10016
rect 77396 9976 77397 10016
rect 77355 9967 77397 9976
rect 77356 9882 77396 9967
rect 77452 9848 77492 10135
rect 77644 10109 77684 10228
rect 77836 10268 77876 10279
rect 77836 10193 77876 10228
rect 78028 10193 78068 10471
rect 82443 10352 82485 10361
rect 82443 10312 82444 10352
rect 82484 10312 82580 10352
rect 82443 10303 82485 10312
rect 82540 10268 82580 10312
rect 82540 10219 82580 10228
rect 82732 10268 82772 10277
rect 77835 10184 77877 10193
rect 77835 10144 77836 10184
rect 77876 10144 77877 10184
rect 77835 10135 77877 10144
rect 78027 10184 78069 10193
rect 78027 10144 78028 10184
rect 78068 10144 78069 10184
rect 78027 10135 78069 10144
rect 82732 10109 82772 10228
rect 77643 10100 77685 10109
rect 77643 10060 77644 10100
rect 77684 10060 77685 10100
rect 77643 10051 77685 10060
rect 82731 10100 82773 10109
rect 82731 10060 82732 10100
rect 82772 10060 82773 10100
rect 82731 10051 82773 10060
rect 77740 10016 77780 10025
rect 77452 9808 77588 9848
rect 77451 9680 77493 9689
rect 77451 9640 77452 9680
rect 77492 9640 77493 9680
rect 77451 9631 77493 9640
rect 77452 9546 77492 9631
rect 76971 9428 77013 9437
rect 76971 9388 76972 9428
rect 77012 9388 77013 9428
rect 76971 9379 77013 9388
rect 77164 9428 77204 9437
rect 76972 9294 77012 9379
rect 77068 9344 77108 9353
rect 76876 8884 77012 8924
rect 76148 8716 76684 8756
rect 76108 8707 76148 8716
rect 76684 8707 76724 8716
rect 76876 8756 76916 8765
rect 76779 8504 76821 8513
rect 76779 8464 76780 8504
rect 76820 8464 76821 8504
rect 76779 8455 76821 8464
rect 76780 8370 76820 8455
rect 76876 8429 76916 8716
rect 76875 8420 76917 8429
rect 76875 8380 76876 8420
rect 76916 8380 76917 8420
rect 76875 8371 76917 8380
rect 76875 8168 76917 8177
rect 76875 8128 76876 8168
rect 76916 8128 76917 8168
rect 76875 8119 76917 8128
rect 76299 7832 76341 7841
rect 76299 7792 76300 7832
rect 76340 7792 76341 7832
rect 76299 7783 76341 7792
rect 75436 7195 75476 7204
rect 75724 7456 76052 7496
rect 75243 7160 75285 7169
rect 75243 7120 75244 7160
rect 75284 7120 75285 7160
rect 75243 7111 75285 7120
rect 75244 7080 75284 7111
rect 75340 6992 75380 7001
rect 75147 6908 75189 6917
rect 75147 6868 75148 6908
rect 75188 6868 75189 6908
rect 75147 6859 75189 6868
rect 75340 6749 75380 6952
rect 75627 6992 75669 7001
rect 75627 6952 75628 6992
rect 75668 6952 75669 6992
rect 75627 6943 75669 6952
rect 75339 6740 75381 6749
rect 75339 6700 75340 6740
rect 75380 6700 75381 6740
rect 75339 6691 75381 6700
rect 75339 6488 75381 6497
rect 75339 6448 75340 6488
rect 75380 6448 75381 6488
rect 75339 6439 75381 6448
rect 75148 6404 75188 6415
rect 75148 6329 75188 6364
rect 75340 6404 75380 6439
rect 75147 6320 75189 6329
rect 75147 6280 75148 6320
rect 75188 6280 75189 6320
rect 75147 6271 75189 6280
rect 75244 6236 75284 6245
rect 75052 5860 75188 5900
rect 74955 5732 74997 5741
rect 74955 5692 74956 5732
rect 74996 5692 74997 5732
rect 74955 5683 74997 5692
rect 75052 5732 75092 5741
rect 74860 5599 74900 5608
rect 74956 5598 74996 5683
rect 75052 5573 75092 5692
rect 75051 5564 75093 5573
rect 75051 5524 75052 5564
rect 75092 5524 75093 5564
rect 75051 5515 75093 5524
rect 75051 5312 75093 5321
rect 75051 5272 75052 5312
rect 75092 5272 75093 5312
rect 75051 5263 75093 5272
rect 74859 4808 74901 4817
rect 74859 4768 74860 4808
rect 74900 4768 74901 4808
rect 74859 4759 74901 4768
rect 74860 4220 74900 4759
rect 74860 4171 74900 4180
rect 75052 4145 75092 5263
rect 75148 4901 75188 5860
rect 75244 5741 75284 6196
rect 75340 6161 75380 6364
rect 75532 6236 75572 6245
rect 75436 6196 75532 6236
rect 75339 6152 75381 6161
rect 75339 6112 75340 6152
rect 75380 6112 75381 6152
rect 75339 6103 75381 6112
rect 75243 5732 75285 5741
rect 75243 5692 75244 5732
rect 75284 5692 75285 5732
rect 75243 5683 75285 5692
rect 75340 5480 75380 5489
rect 75244 5440 75340 5480
rect 75147 4892 75189 4901
rect 75147 4852 75148 4892
rect 75188 4852 75189 4892
rect 75147 4843 75189 4852
rect 75148 4724 75188 4735
rect 75148 4649 75188 4684
rect 75147 4640 75189 4649
rect 75147 4600 75148 4640
rect 75188 4600 75189 4640
rect 75147 4591 75189 4600
rect 75244 4304 75284 5440
rect 75340 5431 75380 5440
rect 75436 4388 75476 6196
rect 75532 6187 75572 6196
rect 75531 5648 75573 5657
rect 75531 5608 75532 5648
rect 75572 5608 75573 5648
rect 75531 5599 75573 5608
rect 75532 5514 75572 5599
rect 75531 4640 75573 4649
rect 75531 4600 75532 4640
rect 75572 4600 75573 4640
rect 75531 4591 75573 4600
rect 75148 4264 75284 4304
rect 75340 4348 75476 4388
rect 75051 4136 75093 4145
rect 75051 4096 75052 4136
rect 75092 4096 75093 4136
rect 75051 4087 75093 4096
rect 74859 4052 74901 4061
rect 74859 4012 74860 4052
rect 74900 4012 74901 4052
rect 74859 4003 74901 4012
rect 74860 3918 74900 4003
rect 75052 3968 75092 3977
rect 74764 3415 74804 3424
rect 74572 3212 74612 3221
rect 74379 3044 74421 3053
rect 74379 3004 74380 3044
rect 74420 3004 74421 3044
rect 74379 2995 74421 3004
rect 74283 2120 74325 2129
rect 74283 2080 74284 2120
rect 74324 2080 74325 2120
rect 74283 2071 74325 2080
rect 73803 1700 73845 1709
rect 73803 1660 73804 1700
rect 73844 1660 73845 1700
rect 73803 1651 73845 1660
rect 74187 1700 74229 1709
rect 74187 1660 74188 1700
rect 74228 1660 74229 1700
rect 74187 1651 74229 1660
rect 73803 1448 73845 1457
rect 73803 1408 73804 1448
rect 73844 1408 73845 1448
rect 73803 1399 73845 1408
rect 73611 944 73653 953
rect 73611 904 73612 944
rect 73652 904 73653 944
rect 73611 895 73653 904
rect 73612 80 73652 895
rect 73804 80 73844 1399
rect 73995 860 74037 869
rect 73995 820 73996 860
rect 74036 820 74037 860
rect 73995 811 74037 820
rect 73996 80 74036 811
rect 74188 80 74228 1651
rect 74380 80 74420 2995
rect 74572 1541 74612 3172
rect 74956 3212 74996 3221
rect 74763 2960 74805 2969
rect 74763 2920 74764 2960
rect 74804 2920 74805 2960
rect 74763 2911 74805 2920
rect 74571 1532 74613 1541
rect 74571 1492 74572 1532
rect 74612 1492 74613 1532
rect 74571 1483 74613 1492
rect 74571 1112 74613 1121
rect 74571 1072 74572 1112
rect 74612 1072 74613 1112
rect 74571 1063 74613 1072
rect 74572 80 74612 1063
rect 74764 80 74804 2911
rect 74956 2717 74996 3172
rect 74955 2708 74997 2717
rect 74955 2668 74956 2708
rect 74996 2668 74997 2708
rect 74955 2659 74997 2668
rect 74955 2540 74997 2549
rect 74955 2500 74956 2540
rect 74996 2500 74997 2540
rect 74955 2491 74997 2500
rect 74956 80 74996 2491
rect 75052 1205 75092 3928
rect 75148 3632 75188 4264
rect 75243 4136 75285 4145
rect 75243 4096 75244 4136
rect 75284 4096 75285 4136
rect 75243 4087 75285 4096
rect 75244 4002 75284 4087
rect 75148 3592 75284 3632
rect 75147 3464 75189 3473
rect 75147 3424 75148 3464
rect 75188 3424 75189 3464
rect 75147 3415 75189 3424
rect 75148 3330 75188 3415
rect 75244 3053 75284 3592
rect 75340 3380 75380 4348
rect 75532 4061 75572 4591
rect 75628 4304 75668 6943
rect 75724 6488 75764 7456
rect 75724 6439 75764 6448
rect 75724 5732 75764 5741
rect 75724 4733 75764 5692
rect 75916 5732 75956 5741
rect 75956 5692 76052 5732
rect 75916 5683 75956 5692
rect 75915 5564 75957 5573
rect 75915 5524 75916 5564
rect 75956 5524 75957 5564
rect 75915 5515 75957 5524
rect 75916 5430 75956 5515
rect 75819 5060 75861 5069
rect 75819 5020 75820 5060
rect 75860 5020 75861 5060
rect 75819 5011 75861 5020
rect 75927 5060 75969 5069
rect 75927 5020 75928 5060
rect 75968 5020 75969 5060
rect 75927 5011 75969 5020
rect 75820 4892 75860 5011
rect 75927 4985 75967 5011
rect 75916 4976 75967 4985
rect 75956 4936 75967 4976
rect 75916 4927 75956 4936
rect 75723 4724 75765 4733
rect 75723 4684 75724 4724
rect 75764 4684 75765 4724
rect 75723 4675 75765 4684
rect 75820 4397 75860 4852
rect 76012 4892 76052 5692
rect 76300 5648 76340 7783
rect 76779 7664 76821 7673
rect 76779 7624 76780 7664
rect 76820 7624 76821 7664
rect 76779 7615 76821 7624
rect 76780 6992 76820 7615
rect 76876 7169 76916 8119
rect 76875 7160 76917 7169
rect 76875 7120 76876 7160
rect 76916 7120 76917 7160
rect 76875 7111 76917 7120
rect 76780 6952 76916 6992
rect 76779 6572 76821 6581
rect 76779 6532 76780 6572
rect 76820 6532 76821 6572
rect 76779 6523 76821 6532
rect 76780 6404 76820 6523
rect 76780 6355 76820 6364
rect 76683 5900 76725 5909
rect 76683 5860 76684 5900
rect 76724 5860 76725 5900
rect 76683 5851 76725 5860
rect 76300 5599 76340 5608
rect 76684 5648 76724 5851
rect 76876 5657 76916 6952
rect 76684 5599 76724 5608
rect 76875 5648 76917 5657
rect 76875 5608 76876 5648
rect 76916 5608 76917 5648
rect 76875 5599 76917 5608
rect 76107 5480 76149 5489
rect 76107 5440 76108 5480
rect 76148 5440 76149 5480
rect 76107 5431 76149 5440
rect 76492 5480 76532 5489
rect 76108 5346 76148 5431
rect 76395 5396 76437 5405
rect 76395 5356 76396 5396
rect 76436 5356 76437 5396
rect 76395 5347 76437 5356
rect 76107 5144 76149 5153
rect 76107 5104 76108 5144
rect 76148 5104 76149 5144
rect 76107 5095 76149 5104
rect 76012 4565 76052 4852
rect 76011 4556 76053 4565
rect 76011 4516 76012 4556
rect 76052 4516 76053 4556
rect 76011 4507 76053 4516
rect 75819 4388 75861 4397
rect 75819 4348 75820 4388
rect 75860 4348 75861 4388
rect 75819 4339 75861 4348
rect 75628 4264 75764 4304
rect 75627 4136 75669 4145
rect 75627 4096 75628 4136
rect 75668 4096 75669 4136
rect 75627 4087 75669 4096
rect 75531 4052 75573 4061
rect 75531 4012 75532 4052
rect 75572 4012 75573 4052
rect 75531 4003 75573 4012
rect 75628 4002 75668 4087
rect 75436 3968 75476 3977
rect 75436 3641 75476 3928
rect 75627 3884 75669 3893
rect 75627 3844 75628 3884
rect 75668 3844 75669 3884
rect 75627 3835 75669 3844
rect 75531 3800 75573 3809
rect 75531 3760 75532 3800
rect 75572 3760 75573 3800
rect 75531 3751 75573 3760
rect 75435 3632 75477 3641
rect 75435 3592 75436 3632
rect 75476 3592 75477 3632
rect 75435 3583 75477 3592
rect 75532 3464 75572 3751
rect 75532 3415 75572 3424
rect 75340 3340 75476 3380
rect 75339 3212 75381 3221
rect 75339 3172 75340 3212
rect 75380 3172 75381 3212
rect 75339 3163 75381 3172
rect 75340 3078 75380 3163
rect 75243 3044 75285 3053
rect 75243 3004 75244 3044
rect 75284 3004 75285 3044
rect 75243 2995 75285 3004
rect 75147 2792 75189 2801
rect 75147 2752 75148 2792
rect 75188 2752 75189 2792
rect 75147 2743 75189 2752
rect 75051 1196 75093 1205
rect 75051 1156 75052 1196
rect 75092 1156 75093 1196
rect 75051 1147 75093 1156
rect 75148 80 75188 2743
rect 75436 2540 75476 3340
rect 75340 2500 75476 2540
rect 75340 80 75380 2500
rect 75531 2456 75573 2465
rect 75531 2416 75532 2456
rect 75572 2416 75573 2456
rect 75531 2407 75573 2416
rect 75532 80 75572 2407
rect 75628 2045 75668 3835
rect 75724 3548 75764 4264
rect 76012 4229 76052 4314
rect 75819 4220 75861 4229
rect 75819 4180 75820 4220
rect 75860 4180 75861 4220
rect 75819 4171 75861 4180
rect 76011 4220 76053 4229
rect 76011 4180 76012 4220
rect 76052 4180 76053 4220
rect 76011 4171 76053 4180
rect 75820 4086 75860 4171
rect 76108 4145 76148 5095
rect 76299 4976 76341 4985
rect 76299 4936 76300 4976
rect 76340 4936 76341 4976
rect 76299 4927 76341 4936
rect 76207 4881 76247 4900
rect 76300 4881 76340 4927
rect 76396 4901 76436 5347
rect 76247 4841 76340 4881
rect 76395 4892 76437 4901
rect 76395 4852 76396 4892
rect 76436 4852 76437 4892
rect 76395 4843 76437 4852
rect 76207 4817 76247 4841
rect 76203 4808 76247 4817
rect 76203 4768 76204 4808
rect 76244 4768 76247 4808
rect 76203 4759 76245 4768
rect 76299 4724 76341 4733
rect 76299 4684 76300 4724
rect 76340 4684 76341 4724
rect 76299 4675 76341 4684
rect 76300 4590 76340 4675
rect 76396 4313 76436 4843
rect 76395 4304 76437 4313
rect 76395 4264 76396 4304
rect 76436 4264 76437 4304
rect 76395 4255 76437 4264
rect 76107 4136 76149 4145
rect 76107 4096 76108 4136
rect 76148 4096 76149 4136
rect 76107 4087 76149 4096
rect 76395 4136 76437 4145
rect 76395 4096 76396 4136
rect 76436 4096 76437 4136
rect 76395 4087 76437 4096
rect 76396 4002 76436 4087
rect 76012 3968 76052 3977
rect 75724 3508 75956 3548
rect 75916 3475 75956 3508
rect 75916 3426 75956 3435
rect 76012 3296 76052 3928
rect 75916 3256 76052 3296
rect 76204 3968 76244 3977
rect 75724 3212 75764 3221
rect 75627 2036 75669 2045
rect 75627 1996 75628 2036
rect 75668 1996 75669 2036
rect 75627 1987 75669 1996
rect 75724 1793 75764 3172
rect 75916 3053 75956 3256
rect 76108 3212 76148 3221
rect 76012 3172 76108 3212
rect 75915 3044 75957 3053
rect 75915 3004 75916 3044
rect 75956 3004 75957 3044
rect 75915 2995 75957 3004
rect 75915 2288 75957 2297
rect 75915 2248 75916 2288
rect 75956 2248 75957 2288
rect 75915 2239 75957 2248
rect 75723 1784 75765 1793
rect 75723 1744 75724 1784
rect 75764 1744 75765 1784
rect 75723 1735 75765 1744
rect 75723 1028 75765 1037
rect 75723 988 75724 1028
rect 75764 988 75765 1028
rect 75723 979 75765 988
rect 75724 80 75764 979
rect 75916 80 75956 2239
rect 76012 1289 76052 3172
rect 76108 3163 76148 3172
rect 76107 2540 76149 2549
rect 76107 2500 76108 2540
rect 76148 2500 76149 2540
rect 76107 2491 76149 2500
rect 76011 1280 76053 1289
rect 76011 1240 76012 1280
rect 76052 1240 76053 1280
rect 76011 1231 76053 1240
rect 76108 80 76148 2491
rect 76204 869 76244 3928
rect 76492 3548 76532 5440
rect 76876 5480 76916 5489
rect 76876 5321 76916 5440
rect 76875 5312 76917 5321
rect 76875 5272 76876 5312
rect 76916 5272 76917 5312
rect 76875 5263 76917 5272
rect 76779 5144 76821 5153
rect 76779 5104 76780 5144
rect 76820 5104 76821 5144
rect 76779 5095 76821 5104
rect 76588 4985 76628 4987
rect 76587 4976 76629 4985
rect 76587 4936 76588 4976
rect 76628 4936 76629 4976
rect 76587 4927 76629 4936
rect 76588 4892 76628 4927
rect 76588 4843 76628 4852
rect 76780 4892 76820 5095
rect 76972 5060 77012 8884
rect 77068 7589 77108 9304
rect 77164 9269 77204 9388
rect 77356 9428 77396 9437
rect 77163 9260 77205 9269
rect 77163 9220 77164 9260
rect 77204 9220 77205 9260
rect 77163 9211 77205 9220
rect 77356 9101 77396 9388
rect 77548 9428 77588 9808
rect 77740 9605 77780 9976
rect 82636 10016 82676 10025
rect 79288 9848 79656 9857
rect 79328 9808 79370 9848
rect 79410 9808 79452 9848
rect 79492 9808 79534 9848
rect 79574 9808 79616 9848
rect 79288 9799 79656 9808
rect 77931 9764 77973 9773
rect 77931 9724 77932 9764
rect 77972 9724 77973 9764
rect 77931 9715 77973 9724
rect 80619 9764 80661 9773
rect 80619 9724 80620 9764
rect 80660 9724 80661 9764
rect 80619 9715 80661 9724
rect 77739 9596 77781 9605
rect 77739 9556 77740 9596
rect 77780 9556 77781 9596
rect 77739 9547 77781 9556
rect 77740 9428 77780 9437
rect 77588 9388 77740 9428
rect 77548 9269 77588 9388
rect 77740 9379 77780 9388
rect 77932 9428 77972 9715
rect 78316 9428 78356 9437
rect 77932 9379 77972 9388
rect 78220 9388 78316 9428
rect 77836 9344 77876 9353
rect 77547 9260 77589 9269
rect 77547 9220 77548 9260
rect 77588 9220 77589 9260
rect 77547 9211 77589 9220
rect 77355 9092 77397 9101
rect 77355 9052 77356 9092
rect 77396 9052 77397 9092
rect 77355 9043 77397 9052
rect 77836 8588 77876 9304
rect 78220 8933 78260 9388
rect 78316 9379 78356 9388
rect 78508 9428 78548 9437
rect 79276 9428 79316 9437
rect 78412 9344 78452 9353
rect 78412 9101 78452 9304
rect 78411 9092 78453 9101
rect 78411 9052 78412 9092
rect 78452 9052 78453 9092
rect 78411 9043 78453 9052
rect 78219 8924 78261 8933
rect 78508 8924 78548 9388
rect 78219 8884 78220 8924
rect 78260 8884 78261 8924
rect 78219 8875 78261 8884
rect 78316 8884 78548 8924
rect 78604 9388 79276 9428
rect 78316 8769 78356 8884
rect 77931 8756 77973 8765
rect 77931 8716 77932 8756
rect 77972 8716 77973 8756
rect 77931 8707 77973 8716
rect 78124 8756 78164 8765
rect 77932 8622 77972 8707
rect 77452 8548 77876 8588
rect 77163 8504 77205 8513
rect 77163 8464 77164 8504
rect 77204 8464 77205 8504
rect 77163 8455 77205 8464
rect 77067 7580 77109 7589
rect 77067 7540 77068 7580
rect 77108 7540 77109 7580
rect 77067 7531 77109 7540
rect 77068 7454 77108 7463
rect 77068 6581 77108 7414
rect 77067 6572 77109 6581
rect 77067 6532 77068 6572
rect 77108 6532 77109 6572
rect 77067 6523 77109 6532
rect 77067 6236 77109 6245
rect 77067 6196 77068 6236
rect 77108 6196 77109 6236
rect 77067 6187 77109 6196
rect 77068 6102 77108 6187
rect 77067 5648 77109 5657
rect 77067 5608 77068 5648
rect 77108 5608 77109 5648
rect 77067 5599 77109 5608
rect 77068 5514 77108 5599
rect 77164 5153 77204 8455
rect 77452 7673 77492 8548
rect 78028 8504 78068 8513
rect 77836 8464 78028 8504
rect 77547 8000 77589 8009
rect 77547 7960 77548 8000
rect 77588 7960 77589 8000
rect 77547 7951 77589 7960
rect 77548 7916 77588 7951
rect 77548 7865 77588 7876
rect 77739 7916 77781 7925
rect 77739 7876 77740 7916
rect 77780 7876 77781 7916
rect 77739 7867 77781 7876
rect 77644 7832 77684 7841
rect 77451 7664 77493 7673
rect 77451 7624 77452 7664
rect 77492 7624 77493 7664
rect 77451 7615 77493 7624
rect 77259 7244 77301 7253
rect 77259 7204 77260 7244
rect 77300 7204 77301 7244
rect 77259 7195 77301 7204
rect 77356 7244 77396 7253
rect 77260 6320 77300 7195
rect 77356 6917 77396 7204
rect 77547 7244 77589 7253
rect 77547 7204 77548 7244
rect 77588 7204 77589 7244
rect 77547 7195 77589 7204
rect 77548 7110 77588 7195
rect 77355 6908 77397 6917
rect 77355 6868 77356 6908
rect 77396 6868 77397 6908
rect 77355 6859 77397 6868
rect 77452 6656 77492 6665
rect 77547 6656 77589 6665
rect 77492 6616 77548 6656
rect 77588 6616 77589 6656
rect 77452 6607 77492 6616
rect 77547 6607 77589 6616
rect 77644 6581 77684 7792
rect 77740 7782 77780 7867
rect 77739 7328 77781 7337
rect 77739 7288 77740 7328
rect 77780 7288 77781 7328
rect 77739 7279 77781 7288
rect 77740 6917 77780 7279
rect 77739 6908 77781 6917
rect 77739 6868 77740 6908
rect 77780 6868 77781 6908
rect 77739 6859 77781 6868
rect 77643 6572 77685 6581
rect 77452 6497 77492 6541
rect 77643 6532 77644 6572
rect 77684 6532 77685 6572
rect 77643 6523 77685 6532
rect 77740 6497 77780 6859
rect 77451 6488 77493 6497
rect 77451 6448 77452 6488
rect 77492 6448 77493 6488
rect 77451 6446 77493 6448
rect 77451 6439 77452 6446
rect 77492 6439 77493 6446
rect 77739 6488 77781 6497
rect 77739 6448 77740 6488
rect 77780 6448 77781 6488
rect 77739 6439 77781 6448
rect 77452 6397 77492 6406
rect 77644 6404 77684 6413
rect 77644 6320 77684 6364
rect 77740 6404 77780 6439
rect 77740 6354 77780 6364
rect 77260 6280 77684 6320
rect 77260 6236 77300 6280
rect 77260 6187 77300 6196
rect 77836 5816 77876 8464
rect 78028 8455 78068 8464
rect 78124 8261 78164 8716
rect 78219 8756 78261 8765
rect 78219 8716 78220 8756
rect 78260 8729 78316 8756
rect 78508 8756 78548 8765
rect 78260 8716 78356 8729
rect 78219 8707 78261 8716
rect 78123 8252 78165 8261
rect 78123 8212 78124 8252
rect 78164 8212 78165 8252
rect 78123 8203 78165 8212
rect 77932 7916 77972 7925
rect 77932 7757 77972 7876
rect 78124 7916 78164 7925
rect 78220 7916 78260 8707
rect 78316 8634 78356 8716
rect 78507 8716 78508 8756
rect 78507 8707 78548 8716
rect 78507 8597 78547 8707
rect 78506 8588 78548 8597
rect 78506 8548 78507 8588
rect 78547 8548 78548 8588
rect 78506 8539 78548 8548
rect 78411 8504 78453 8513
rect 78411 8464 78412 8504
rect 78452 8464 78453 8504
rect 78411 8455 78453 8464
rect 78412 8370 78452 8455
rect 78411 7916 78453 7925
rect 78164 7876 78412 7916
rect 78452 7876 78453 7916
rect 78124 7867 78164 7876
rect 78027 7832 78069 7841
rect 78027 7792 78028 7832
rect 78068 7792 78069 7832
rect 78027 7783 78069 7792
rect 77931 7748 77973 7757
rect 77931 7708 77932 7748
rect 77972 7708 77973 7748
rect 77931 7699 77973 7708
rect 78028 7698 78068 7783
rect 78220 7244 78260 7876
rect 78411 7867 78453 7876
rect 78604 7916 78644 9388
rect 79276 9379 79316 9388
rect 80235 9428 80277 9437
rect 80235 9388 80236 9428
rect 80276 9388 80277 9428
rect 80235 9379 80277 9388
rect 80620 9428 80660 9715
rect 81867 9596 81909 9605
rect 81867 9556 81868 9596
rect 81908 9556 81909 9596
rect 81867 9547 81909 9556
rect 80812 9437 80852 9522
rect 81004 9437 81044 9522
rect 80620 9379 80660 9388
rect 80811 9428 80853 9437
rect 80811 9388 80812 9428
rect 80852 9388 80853 9428
rect 80811 9379 80853 9388
rect 81003 9428 81045 9437
rect 81003 9388 81004 9428
rect 81044 9388 81045 9428
rect 81003 9379 81045 9388
rect 81196 9428 81236 9439
rect 80236 9294 80276 9379
rect 81196 9353 81236 9388
rect 81868 9428 81908 9547
rect 82059 9512 82101 9521
rect 82059 9472 82060 9512
rect 82100 9472 82101 9512
rect 82059 9463 82101 9472
rect 80716 9344 80756 9353
rect 80716 9260 80756 9304
rect 81100 9344 81140 9353
rect 80716 9220 81044 9260
rect 80528 9092 80896 9101
rect 80568 9052 80610 9092
rect 80650 9052 80692 9092
rect 80732 9052 80774 9092
rect 80814 9052 80856 9092
rect 80528 9043 80896 9052
rect 81004 8924 81044 9220
rect 81100 9101 81140 9304
rect 81195 9344 81237 9353
rect 81195 9304 81196 9344
rect 81236 9304 81237 9344
rect 81195 9295 81237 9304
rect 81483 9344 81525 9353
rect 81483 9304 81484 9344
rect 81524 9304 81525 9344
rect 81483 9295 81525 9304
rect 81099 9092 81141 9101
rect 81099 9052 81100 9092
rect 81140 9052 81141 9092
rect 81099 9043 81141 9052
rect 81291 8924 81333 8933
rect 81004 8884 81140 8924
rect 78795 8840 78837 8849
rect 78795 8800 78796 8840
rect 78836 8800 78837 8840
rect 78795 8791 78837 8800
rect 78987 8840 79029 8849
rect 78987 8800 78988 8840
rect 79028 8800 79029 8840
rect 78987 8791 79029 8800
rect 80907 8840 80949 8849
rect 80907 8800 80908 8840
rect 80948 8800 80949 8840
rect 80907 8791 80949 8800
rect 78700 8756 78740 8767
rect 78700 8681 78740 8716
rect 78796 8706 78836 8791
rect 78891 8756 78933 8765
rect 78891 8716 78892 8756
rect 78932 8716 78933 8756
rect 78891 8707 78933 8716
rect 78699 8672 78741 8681
rect 78699 8632 78700 8672
rect 78740 8632 78741 8672
rect 78699 8623 78741 8632
rect 78892 8622 78932 8707
rect 78988 8345 79028 8791
rect 80811 8756 80853 8765
rect 80716 8716 80812 8756
rect 80852 8716 80853 8756
rect 78987 8336 79029 8345
rect 78987 8296 78988 8336
rect 79028 8296 79029 8336
rect 78987 8287 79029 8296
rect 79288 8336 79656 8345
rect 79328 8296 79370 8336
rect 79410 8296 79452 8336
rect 79492 8296 79534 8336
rect 79574 8296 79616 8336
rect 79288 8287 79656 8296
rect 78987 8084 79029 8093
rect 78987 8044 78988 8084
rect 79028 8044 79029 8084
rect 78987 8035 79029 8044
rect 78412 7782 78452 7867
rect 78315 7664 78357 7673
rect 78315 7624 78316 7664
rect 78356 7624 78357 7664
rect 78315 7615 78357 7624
rect 78028 7221 78068 7230
rect 78220 7195 78260 7204
rect 78028 7169 78068 7181
rect 78027 7160 78069 7169
rect 78027 7120 78028 7160
rect 78068 7120 78069 7160
rect 78027 7111 78069 7120
rect 78028 7086 78068 7111
rect 78124 6992 78164 7001
rect 77740 5776 77876 5816
rect 77932 6952 78124 6992
rect 77260 5732 77300 5741
rect 77452 5732 77492 5741
rect 77163 5144 77205 5153
rect 77163 5104 77164 5144
rect 77204 5104 77205 5144
rect 77163 5095 77205 5104
rect 76780 4843 76820 4852
rect 76876 5020 77012 5060
rect 76684 4724 76724 4733
rect 76779 4724 76821 4733
rect 76724 4684 76780 4724
rect 76820 4684 76821 4724
rect 76684 4675 76724 4684
rect 76779 4675 76821 4684
rect 76683 4556 76725 4565
rect 76683 4516 76684 4556
rect 76724 4516 76725 4556
rect 76683 4507 76725 4516
rect 76587 4388 76629 4397
rect 76587 4348 76588 4388
rect 76628 4348 76629 4388
rect 76587 4339 76629 4348
rect 76588 4220 76628 4339
rect 76588 4171 76628 4180
rect 76684 4145 76724 4507
rect 76779 4388 76821 4397
rect 76779 4348 76780 4388
rect 76820 4348 76821 4388
rect 76779 4339 76821 4348
rect 76780 4229 76820 4339
rect 76779 4220 76821 4229
rect 76779 4180 76780 4220
rect 76820 4180 76821 4220
rect 76779 4171 76821 4180
rect 76683 4136 76725 4145
rect 76683 4096 76684 4136
rect 76724 4096 76725 4136
rect 76683 4087 76725 4096
rect 76780 3968 76820 3977
rect 76683 3632 76725 3641
rect 76683 3592 76684 3632
rect 76724 3592 76725 3632
rect 76683 3583 76725 3592
rect 76492 3508 76628 3548
rect 76299 3464 76341 3473
rect 76299 3424 76300 3464
rect 76340 3424 76341 3464
rect 76299 3415 76341 3424
rect 76300 3330 76340 3415
rect 76492 3212 76532 3221
rect 76396 3172 76492 3212
rect 76299 1196 76341 1205
rect 76299 1156 76300 1196
rect 76340 1156 76341 1196
rect 76299 1147 76341 1156
rect 76203 860 76245 869
rect 76203 820 76204 860
rect 76244 820 76245 860
rect 76203 811 76245 820
rect 76300 80 76340 1147
rect 76396 953 76436 3172
rect 76492 3163 76532 3172
rect 76491 2876 76533 2885
rect 76491 2836 76492 2876
rect 76532 2836 76533 2876
rect 76491 2827 76533 2836
rect 76395 944 76437 953
rect 76395 904 76396 944
rect 76436 904 76437 944
rect 76395 895 76437 904
rect 76492 80 76532 2827
rect 76588 2465 76628 3508
rect 76684 3464 76724 3583
rect 76684 3415 76724 3424
rect 76780 2465 76820 3928
rect 76876 3464 76916 5020
rect 77260 4901 77300 5692
rect 77356 5692 77452 5732
rect 77356 5405 77396 5692
rect 77452 5683 77492 5692
rect 77451 5480 77493 5489
rect 77451 5440 77452 5480
rect 77492 5440 77493 5480
rect 77451 5431 77493 5440
rect 77355 5396 77397 5405
rect 77355 5356 77356 5396
rect 77396 5356 77397 5396
rect 77355 5347 77397 5356
rect 77452 5346 77492 5431
rect 77740 5237 77780 5776
rect 77836 5648 77876 5657
rect 77836 5489 77876 5608
rect 77835 5480 77877 5489
rect 77835 5440 77836 5480
rect 77876 5440 77877 5480
rect 77835 5431 77877 5440
rect 77547 5228 77589 5237
rect 77547 5188 77548 5228
rect 77588 5188 77589 5228
rect 77547 5179 77589 5188
rect 77739 5228 77781 5237
rect 77739 5188 77740 5228
rect 77780 5188 77781 5228
rect 77739 5179 77781 5188
rect 77451 5144 77493 5153
rect 77451 5104 77452 5144
rect 77492 5104 77493 5144
rect 77451 5095 77493 5104
rect 76971 4892 77013 4901
rect 76971 4852 76972 4892
rect 77012 4852 77013 4892
rect 76971 4843 77013 4852
rect 77164 4892 77204 4901
rect 76972 4758 77012 4843
rect 77068 4724 77108 4733
rect 77068 3893 77108 4684
rect 77164 4397 77204 4852
rect 77259 4892 77301 4901
rect 77259 4852 77260 4892
rect 77300 4852 77301 4892
rect 77259 4843 77301 4852
rect 77356 4724 77396 4733
rect 77260 4684 77356 4724
rect 77163 4388 77205 4397
rect 77163 4348 77164 4388
rect 77204 4348 77205 4388
rect 77163 4339 77205 4348
rect 77164 4220 77204 4231
rect 77164 4145 77204 4180
rect 77163 4136 77205 4145
rect 77163 4096 77164 4136
rect 77204 4096 77205 4136
rect 77163 4087 77205 4096
rect 77067 3884 77109 3893
rect 77067 3844 77068 3884
rect 77108 3844 77109 3884
rect 77067 3835 77109 3844
rect 77260 3632 77300 4684
rect 77356 4675 77396 4684
rect 77355 4220 77397 4229
rect 77355 4180 77356 4220
rect 77396 4180 77397 4220
rect 77355 4171 77397 4180
rect 77356 4086 77396 4171
rect 77164 3592 77300 3632
rect 77355 3632 77397 3641
rect 77355 3592 77356 3632
rect 77396 3592 77397 3632
rect 77068 3464 77108 3473
rect 76876 3424 77068 3464
rect 77068 3415 77108 3424
rect 76971 3296 77013 3305
rect 76971 3256 76972 3296
rect 77012 3256 77013 3296
rect 76971 3247 77013 3256
rect 76876 3212 76916 3221
rect 76587 2456 76629 2465
rect 76587 2416 76588 2456
rect 76628 2416 76629 2456
rect 76587 2407 76629 2416
rect 76779 2456 76821 2465
rect 76779 2416 76780 2456
rect 76820 2416 76821 2456
rect 76779 2407 76821 2416
rect 76683 2372 76725 2381
rect 76683 2332 76684 2372
rect 76724 2332 76725 2372
rect 76683 2323 76725 2332
rect 76684 80 76724 2323
rect 76876 1457 76916 3172
rect 76875 1448 76917 1457
rect 76875 1408 76876 1448
rect 76916 1408 76917 1448
rect 76875 1399 76917 1408
rect 76972 1280 77012 3247
rect 77164 2297 77204 3592
rect 77355 3583 77397 3592
rect 77260 3212 77300 3221
rect 77163 2288 77205 2297
rect 77163 2248 77164 2288
rect 77204 2248 77205 2288
rect 77163 2239 77205 2248
rect 77260 1709 77300 3172
rect 77259 1700 77301 1709
rect 77259 1660 77260 1700
rect 77300 1660 77301 1700
rect 77259 1651 77301 1660
rect 77356 1532 77396 3583
rect 77452 3464 77492 5095
rect 77548 4976 77588 5179
rect 77548 4927 77588 4936
rect 77835 4892 77877 4901
rect 77835 4852 77836 4892
rect 77876 4852 77877 4892
rect 77835 4843 77877 4852
rect 77836 4758 77876 4843
rect 77643 4304 77685 4313
rect 77643 4264 77644 4304
rect 77684 4264 77685 4304
rect 77643 4255 77685 4264
rect 77644 4170 77684 4255
rect 77739 3800 77781 3809
rect 77739 3760 77740 3800
rect 77780 3760 77781 3800
rect 77739 3751 77781 3760
rect 77452 3415 77492 3424
rect 76876 1240 77012 1280
rect 77260 1492 77396 1532
rect 77644 3212 77684 3221
rect 76876 80 76916 1240
rect 77067 1028 77109 1037
rect 77067 988 77068 1028
rect 77108 988 77109 1028
rect 77067 979 77109 988
rect 77068 80 77108 979
rect 77260 80 77300 1492
rect 77451 1280 77493 1289
rect 77451 1240 77452 1280
rect 77492 1240 77493 1280
rect 77451 1231 77493 1240
rect 77452 80 77492 1231
rect 77644 1121 77684 3172
rect 77740 3137 77780 3751
rect 77836 3464 77876 3473
rect 77932 3464 77972 6952
rect 78124 6943 78164 6952
rect 78219 6572 78261 6581
rect 78219 6532 78220 6572
rect 78260 6532 78261 6572
rect 78219 6523 78261 6532
rect 78027 6488 78069 6497
rect 78027 6448 78028 6488
rect 78068 6448 78069 6488
rect 78027 6439 78069 6448
rect 78028 5732 78068 6439
rect 78028 5683 78068 5692
rect 78027 5480 78069 5489
rect 78027 5440 78028 5480
rect 78068 5440 78069 5480
rect 78027 5431 78069 5440
rect 78028 5346 78068 5431
rect 78027 5144 78069 5153
rect 78027 5104 78028 5144
rect 78068 5104 78069 5144
rect 78027 5095 78069 5104
rect 78028 4892 78068 5095
rect 78028 4843 78068 4852
rect 78027 3884 78069 3893
rect 78027 3844 78028 3884
rect 78068 3844 78069 3884
rect 78027 3835 78069 3844
rect 77876 3424 77972 3464
rect 77836 3415 77876 3424
rect 78028 3380 78068 3835
rect 78220 3809 78260 6523
rect 78316 5657 78356 7615
rect 78412 7412 78452 7421
rect 78412 6329 78452 7372
rect 78508 7337 78548 7339
rect 78507 7328 78549 7337
rect 78507 7288 78508 7328
rect 78548 7288 78549 7328
rect 78507 7279 78549 7288
rect 78508 7244 78548 7279
rect 78604 7253 78644 7876
rect 78795 7916 78837 7925
rect 78795 7876 78796 7916
rect 78836 7876 78837 7916
rect 78795 7867 78837 7876
rect 78988 7916 79028 8035
rect 80716 7925 80756 8716
rect 80811 8707 80853 8716
rect 80812 8622 80852 8707
rect 80908 8706 80948 8791
rect 81004 8756 81044 8765
rect 80907 8504 80949 8513
rect 80907 8464 80908 8504
rect 80948 8464 80949 8504
rect 80907 8455 80949 8464
rect 80908 8177 80948 8455
rect 81004 8429 81044 8716
rect 81003 8420 81045 8429
rect 81003 8380 81004 8420
rect 81044 8380 81045 8420
rect 81003 8371 81045 8380
rect 81004 8261 81044 8371
rect 81003 8252 81045 8261
rect 81003 8212 81004 8252
rect 81044 8212 81045 8252
rect 81003 8203 81045 8212
rect 80907 8168 80949 8177
rect 80907 8128 80908 8168
rect 80948 8128 80949 8168
rect 80907 8119 80949 8128
rect 78988 7867 79028 7876
rect 80715 7916 80757 7925
rect 80715 7876 80716 7916
rect 80756 7876 80757 7916
rect 80715 7867 80757 7876
rect 80908 7916 80948 8119
rect 81100 8084 81140 8884
rect 81291 8884 81292 8924
rect 81332 8884 81333 8924
rect 81291 8875 81333 8884
rect 81195 8756 81237 8765
rect 81195 8716 81196 8756
rect 81236 8716 81237 8756
rect 81195 8707 81237 8716
rect 81292 8756 81332 8875
rect 81484 8849 81524 9295
rect 81675 9260 81717 9269
rect 81675 9220 81676 9260
rect 81716 9220 81717 9260
rect 81675 9211 81717 9220
rect 81483 8840 81525 8849
rect 81483 8800 81484 8840
rect 81524 8800 81525 8840
rect 81483 8791 81525 8800
rect 81676 8840 81716 9211
rect 81868 9185 81908 9388
rect 82060 9428 82100 9463
rect 82060 9377 82100 9388
rect 81964 9344 82004 9353
rect 81964 9260 82004 9304
rect 81964 9220 82292 9260
rect 81867 9176 81909 9185
rect 81867 9136 81868 9176
rect 81908 9136 81909 9176
rect 81867 9127 81909 9136
rect 82059 9008 82101 9017
rect 82059 8968 82060 9008
rect 82100 8968 82101 9008
rect 82059 8959 82101 8968
rect 81676 8791 81716 8800
rect 82060 8840 82100 8959
rect 82060 8791 82100 8800
rect 81292 8707 81332 8716
rect 81388 8756 81428 8767
rect 81196 8622 81236 8707
rect 81388 8681 81428 8716
rect 81579 8756 81621 8765
rect 81579 8716 81580 8756
rect 81620 8716 81621 8756
rect 81579 8707 81621 8716
rect 81772 8756 81812 8765
rect 81387 8672 81429 8681
rect 81387 8632 81388 8672
rect 81428 8632 81429 8672
rect 81387 8623 81429 8632
rect 81580 8622 81620 8707
rect 81772 8597 81812 8716
rect 81963 8756 82005 8765
rect 81963 8716 81964 8756
rect 82004 8716 82005 8756
rect 81963 8707 82005 8716
rect 82155 8756 82197 8765
rect 82155 8716 82156 8756
rect 82196 8716 82197 8756
rect 82155 8707 82197 8716
rect 81964 8622 82004 8707
rect 82156 8622 82196 8707
rect 81771 8588 81813 8597
rect 81771 8548 81772 8588
rect 81812 8548 81813 8588
rect 81771 8539 81813 8548
rect 81579 8336 81621 8345
rect 81579 8296 81580 8336
rect 81620 8296 81621 8336
rect 81579 8287 81621 8296
rect 81580 8168 81620 8287
rect 81772 8177 81812 8539
rect 81580 8119 81620 8128
rect 81771 8168 81813 8177
rect 81771 8128 81772 8168
rect 81812 8128 81813 8168
rect 81771 8119 81813 8128
rect 80908 7867 80948 7876
rect 81004 8044 81140 8084
rect 81675 8084 81717 8093
rect 81675 8044 81676 8084
rect 81716 8044 81717 8084
rect 78796 7782 78836 7867
rect 78892 7832 78932 7841
rect 78892 7580 78932 7792
rect 80716 7782 80756 7867
rect 80811 7832 80853 7841
rect 80811 7792 80812 7832
rect 80852 7792 80853 7832
rect 80811 7783 80853 7792
rect 80812 7698 80852 7783
rect 80528 7580 80896 7589
rect 78892 7540 79124 7580
rect 78891 7412 78933 7421
rect 78891 7372 78892 7412
rect 78932 7372 78933 7412
rect 78891 7363 78933 7372
rect 78699 7328 78741 7337
rect 78699 7288 78700 7328
rect 78740 7288 78741 7328
rect 78699 7279 78741 7288
rect 78508 7195 78548 7204
rect 78603 7244 78645 7253
rect 78603 7204 78604 7244
rect 78644 7204 78645 7244
rect 78603 7195 78645 7204
rect 78700 7194 78740 7279
rect 78892 7278 78932 7363
rect 78988 7244 79028 7253
rect 78507 7076 78549 7085
rect 78507 7036 78508 7076
rect 78548 7036 78549 7076
rect 78507 7027 78549 7036
rect 78411 6320 78453 6329
rect 78411 6280 78412 6320
rect 78452 6280 78453 6320
rect 78411 6271 78453 6280
rect 78508 6161 78548 7027
rect 78988 7001 79028 7204
rect 78987 6992 79029 7001
rect 78987 6952 78988 6992
rect 79028 6952 79029 6992
rect 78987 6943 79029 6952
rect 78699 6908 78741 6917
rect 78699 6868 78700 6908
rect 78740 6868 78741 6908
rect 78699 6859 78741 6868
rect 78603 6656 78645 6665
rect 78603 6616 78604 6656
rect 78644 6616 78645 6656
rect 78603 6607 78645 6616
rect 78507 6152 78549 6161
rect 78507 6112 78508 6152
rect 78548 6112 78549 6152
rect 78507 6103 78549 6112
rect 78411 6068 78453 6077
rect 78411 6028 78412 6068
rect 78452 6028 78453 6068
rect 78411 6019 78453 6028
rect 78412 5741 78452 6019
rect 78507 5984 78549 5993
rect 78507 5944 78508 5984
rect 78548 5944 78549 5984
rect 78507 5935 78549 5944
rect 78411 5732 78453 5741
rect 78411 5692 78412 5732
rect 78452 5692 78453 5732
rect 78411 5683 78453 5692
rect 78508 5732 78548 5935
rect 78508 5683 78548 5692
rect 78315 5648 78357 5657
rect 78315 5608 78316 5648
rect 78356 5608 78357 5648
rect 78315 5599 78357 5608
rect 78411 5480 78453 5489
rect 78411 5440 78412 5480
rect 78452 5440 78453 5480
rect 78411 5431 78453 5440
rect 78316 4724 78356 4733
rect 78219 3800 78261 3809
rect 78219 3760 78220 3800
rect 78260 3760 78261 3800
rect 78219 3751 78261 3760
rect 78219 3548 78261 3557
rect 78219 3508 78220 3548
rect 78260 3508 78261 3548
rect 78219 3499 78261 3508
rect 78220 3464 78260 3499
rect 78220 3413 78260 3424
rect 77932 3340 78068 3380
rect 77739 3128 77781 3137
rect 77739 3088 77740 3128
rect 77780 3088 77781 3128
rect 77739 3079 77781 3088
rect 77932 2036 77972 3340
rect 78028 3212 78068 3221
rect 78028 2969 78068 3172
rect 78027 2960 78069 2969
rect 78027 2920 78028 2960
rect 78068 2920 78069 2960
rect 78027 2911 78069 2920
rect 78316 2540 78356 4684
rect 78412 4229 78452 5431
rect 78507 5060 78549 5069
rect 78507 5020 78508 5060
rect 78548 5020 78549 5060
rect 78507 5011 78549 5020
rect 78508 4976 78548 5011
rect 78508 4925 78548 4936
rect 78604 4881 78644 6607
rect 78700 6413 78740 6859
rect 79084 6572 79124 7540
rect 80568 7540 80610 7580
rect 80650 7540 80692 7580
rect 80732 7540 80774 7580
rect 80814 7540 80856 7580
rect 80528 7531 80896 7540
rect 80427 7496 80469 7505
rect 80427 7456 80428 7496
rect 80468 7456 80469 7496
rect 80427 7447 80469 7456
rect 79179 7412 79221 7421
rect 79179 7372 79180 7412
rect 79220 7372 79221 7412
rect 79179 7363 79221 7372
rect 79180 7278 79220 7363
rect 79179 6992 79221 7001
rect 79179 6952 79180 6992
rect 79220 6952 79221 6992
rect 79179 6943 79221 6952
rect 79180 6833 79220 6943
rect 79179 6824 79221 6833
rect 79179 6784 79180 6824
rect 79220 6784 79221 6824
rect 79179 6775 79221 6784
rect 79288 6824 79656 6833
rect 79328 6784 79370 6824
rect 79410 6784 79452 6824
rect 79492 6784 79534 6824
rect 79574 6784 79616 6824
rect 79288 6775 79656 6784
rect 78988 6532 79124 6572
rect 78795 6488 78837 6497
rect 78795 6448 78796 6488
rect 78836 6448 78837 6488
rect 78795 6439 78837 6448
rect 78699 6404 78741 6413
rect 78699 6364 78700 6404
rect 78740 6364 78741 6404
rect 78699 6355 78741 6364
rect 78700 6270 78740 6355
rect 78796 6354 78836 6439
rect 78892 6404 78932 6413
rect 78795 6152 78837 6161
rect 78795 6112 78796 6152
rect 78836 6112 78837 6152
rect 78795 6103 78837 6112
rect 78796 5900 78836 6103
rect 78892 6077 78932 6364
rect 78891 6068 78933 6077
rect 78891 6028 78892 6068
rect 78932 6028 78933 6068
rect 78891 6019 78933 6028
rect 78891 5900 78933 5909
rect 78796 5860 78892 5900
rect 78932 5860 78933 5900
rect 78891 5851 78933 5860
rect 78700 5732 78740 5741
rect 78795 5732 78837 5741
rect 78740 5692 78796 5732
rect 78836 5692 78837 5732
rect 78700 5683 78740 5692
rect 78795 5683 78837 5692
rect 78892 5732 78932 5851
rect 78892 5683 78932 5692
rect 78699 5480 78741 5489
rect 78699 5440 78700 5480
rect 78740 5440 78741 5480
rect 78699 5431 78741 5440
rect 78700 5346 78740 5431
rect 78796 5153 78836 5683
rect 78795 5144 78837 5153
rect 78795 5104 78796 5144
rect 78836 5104 78837 5144
rect 78795 5095 78837 5104
rect 78892 4976 78932 4985
rect 78988 4976 79028 6532
rect 79180 6488 79220 6775
rect 79276 6581 79316 6666
rect 79467 6656 79509 6665
rect 79467 6616 79468 6656
rect 79508 6616 79509 6656
rect 79467 6607 79509 6616
rect 79275 6572 79317 6581
rect 79275 6532 79276 6572
rect 79316 6532 79317 6572
rect 79275 6523 79317 6532
rect 79468 6522 79508 6607
rect 79851 6572 79893 6581
rect 79851 6532 79852 6572
rect 79892 6532 79893 6572
rect 79851 6523 79893 6532
rect 80236 6572 80276 6581
rect 79660 6488 79700 6497
rect 79084 6448 79220 6488
rect 79564 6448 79660 6488
rect 79084 6404 79124 6448
rect 79084 6355 79124 6364
rect 79276 6404 79316 6413
rect 79276 6320 79316 6364
rect 79564 6320 79604 6448
rect 79660 6439 79700 6448
rect 79852 6438 79892 6523
rect 80044 6488 80084 6497
rect 79180 6280 79316 6320
rect 79372 6280 79604 6320
rect 79083 6068 79125 6077
rect 79180 6068 79220 6280
rect 79372 6236 79412 6280
rect 79083 6028 79084 6068
rect 79124 6028 79220 6068
rect 79276 6196 79412 6236
rect 79659 6236 79701 6245
rect 79659 6196 79660 6236
rect 79700 6196 79701 6236
rect 79083 6019 79125 6028
rect 79084 5741 79124 6019
rect 79276 5984 79316 6196
rect 79659 6187 79701 6196
rect 79371 6068 79413 6077
rect 79371 6028 79372 6068
rect 79412 6028 79413 6068
rect 79371 6019 79413 6028
rect 79180 5944 79316 5984
rect 79083 5732 79125 5741
rect 79083 5692 79084 5732
rect 79124 5692 79125 5732
rect 79083 5683 79125 5692
rect 79084 5564 79124 5573
rect 79180 5564 79220 5944
rect 79372 5900 79412 6019
rect 79372 5851 79412 5860
rect 79276 5732 79316 5743
rect 79276 5657 79316 5692
rect 79467 5732 79509 5741
rect 79467 5692 79468 5732
rect 79508 5692 79509 5732
rect 79467 5683 79509 5692
rect 79660 5732 79700 6187
rect 80044 6077 80084 6448
rect 80139 6488 80181 6497
rect 80139 6448 80140 6488
rect 80180 6448 80181 6488
rect 80139 6439 80181 6448
rect 80043 6068 80085 6077
rect 80043 6028 80044 6068
rect 80084 6028 80085 6068
rect 80043 6019 80085 6028
rect 79660 5683 79700 5692
rect 79851 5732 79893 5741
rect 79851 5692 79852 5732
rect 79892 5692 79893 5732
rect 79851 5683 79893 5692
rect 80043 5732 80085 5741
rect 80043 5692 80044 5732
rect 80084 5692 80085 5732
rect 80043 5683 80085 5692
rect 79275 5648 79317 5657
rect 79275 5608 79276 5648
rect 79316 5608 79317 5648
rect 79275 5599 79317 5608
rect 79468 5598 79508 5683
rect 79852 5598 79892 5683
rect 80044 5598 80084 5683
rect 79124 5524 79220 5564
rect 79084 5515 79124 5524
rect 79755 5480 79797 5489
rect 79755 5440 79756 5480
rect 79796 5440 79797 5480
rect 79755 5431 79797 5440
rect 79852 5480 79892 5489
rect 79083 5312 79125 5321
rect 79083 5272 79084 5312
rect 79124 5272 79125 5312
rect 79083 5263 79125 5272
rect 79288 5312 79656 5321
rect 79328 5272 79370 5312
rect 79410 5272 79452 5312
rect 79492 5272 79534 5312
rect 79574 5272 79616 5312
rect 79288 5263 79656 5272
rect 78932 4936 79028 4976
rect 78892 4927 78932 4936
rect 78604 4841 78932 4881
rect 78700 4724 78740 4733
rect 78411 4220 78453 4229
rect 78411 4180 78412 4220
rect 78452 4180 78453 4220
rect 78411 4171 78453 4180
rect 78412 4086 78452 4171
rect 78700 3641 78740 4684
rect 78796 4220 78836 4229
rect 78796 4145 78836 4180
rect 78794 4136 78836 4145
rect 78794 4096 78795 4136
rect 78835 4096 78836 4136
rect 78794 4087 78836 4096
rect 78796 3968 78836 3977
rect 78699 3632 78741 3641
rect 78699 3592 78700 3632
rect 78740 3592 78741 3632
rect 78699 3583 78741 3592
rect 78796 3473 78836 3928
rect 78603 3464 78645 3473
rect 78603 3424 78604 3464
rect 78644 3424 78645 3464
rect 78603 3415 78645 3424
rect 78795 3464 78837 3473
rect 78795 3424 78796 3464
rect 78836 3424 78837 3464
rect 78795 3415 78837 3424
rect 78604 3330 78644 3415
rect 78892 3296 78932 4841
rect 78987 4472 79029 4481
rect 78987 4432 78988 4472
rect 79028 4432 79029 4472
rect 78987 4423 79029 4432
rect 78988 4220 79028 4423
rect 79084 4313 79124 5263
rect 79371 5144 79413 5153
rect 79371 5104 79372 5144
rect 79412 5104 79413 5144
rect 79371 5095 79413 5104
rect 79276 4985 79316 5016
rect 79275 4976 79317 4985
rect 79275 4936 79276 4976
rect 79316 4936 79317 4976
rect 79275 4927 79317 4936
rect 79276 4892 79316 4927
rect 79372 4892 79412 5095
rect 79468 5069 79508 5154
rect 79563 5144 79605 5153
rect 79563 5104 79564 5144
rect 79604 5104 79605 5144
rect 79563 5095 79605 5104
rect 79467 5060 79509 5069
rect 79467 5020 79468 5060
rect 79508 5020 79509 5060
rect 79467 5011 79509 5020
rect 79468 4892 79508 4901
rect 79372 4852 79468 4892
rect 79276 4481 79316 4852
rect 79468 4843 79508 4852
rect 79564 4724 79604 5095
rect 79372 4684 79604 4724
rect 79660 4724 79700 4733
rect 79275 4472 79317 4481
rect 79275 4432 79276 4472
rect 79316 4432 79317 4472
rect 79275 4423 79317 4432
rect 79083 4304 79125 4313
rect 79083 4264 79084 4304
rect 79124 4264 79125 4304
rect 79083 4255 79125 4264
rect 78988 4145 79028 4180
rect 78987 4136 79029 4145
rect 78987 4096 78988 4136
rect 79028 4096 79029 4136
rect 78987 4087 79029 4096
rect 79372 4136 79412 4684
rect 79372 4087 79412 4096
rect 78988 4056 79028 4087
rect 79564 3977 79604 4062
rect 79180 3968 79220 3977
rect 78987 3800 79029 3809
rect 78987 3760 78988 3800
rect 79028 3760 79029 3800
rect 78987 3751 79029 3760
rect 78988 3464 79028 3751
rect 78988 3415 79028 3424
rect 79180 3389 79220 3928
rect 79563 3968 79605 3977
rect 79563 3928 79564 3968
rect 79604 3928 79605 3968
rect 79660 3968 79700 4684
rect 79756 4136 79796 5431
rect 79852 5237 79892 5440
rect 80044 5480 80084 5489
rect 79851 5228 79893 5237
rect 79851 5188 79852 5228
rect 79892 5188 79893 5228
rect 79851 5179 79893 5188
rect 80044 5069 80084 5440
rect 79851 5060 79893 5069
rect 79851 5020 79852 5060
rect 79892 5020 79893 5060
rect 79851 5011 79893 5020
rect 80043 5060 80085 5069
rect 80043 5020 80044 5060
rect 80084 5020 80085 5060
rect 80043 5011 80085 5020
rect 79852 4976 79892 5011
rect 79852 4925 79892 4936
rect 80044 4724 80084 4733
rect 80044 4145 80084 4684
rect 79756 4087 79796 4096
rect 80043 4136 80085 4145
rect 80043 4096 80044 4136
rect 80084 4096 80085 4136
rect 80043 4087 80085 4096
rect 80140 4136 80180 6439
rect 80236 6329 80276 6532
rect 80331 6488 80373 6497
rect 80331 6448 80332 6488
rect 80372 6448 80373 6488
rect 80331 6439 80373 6448
rect 80428 6488 80468 7447
rect 81004 7412 81044 8044
rect 81675 8035 81717 8044
rect 82155 8084 82197 8093
rect 82155 8044 82156 8084
rect 82196 8044 82197 8084
rect 82155 8035 82197 8044
rect 81098 7916 81140 7925
rect 81098 7876 81099 7916
rect 81098 7867 81140 7876
rect 81099 7782 81140 7867
rect 81292 7916 81332 7925
rect 80908 7372 81044 7412
rect 80811 7328 80853 7337
rect 80811 7288 80812 7328
rect 80852 7288 80853 7328
rect 80811 7279 80853 7288
rect 80812 7244 80852 7279
rect 80812 7193 80852 7204
rect 80428 6439 80468 6448
rect 80235 6320 80277 6329
rect 80235 6280 80236 6320
rect 80276 6280 80277 6320
rect 80235 6271 80277 6280
rect 80235 5816 80277 5825
rect 80235 5776 80236 5816
rect 80276 5776 80277 5816
rect 80235 5767 80277 5776
rect 80236 5732 80276 5767
rect 80236 5681 80276 5692
rect 80236 4976 80276 4985
rect 80332 4976 80372 6439
rect 80427 6320 80469 6329
rect 80427 6280 80428 6320
rect 80468 6280 80469 6320
rect 80908 6320 80948 7372
rect 81004 7244 81044 7253
rect 81100 7244 81140 7782
rect 81196 7832 81236 7841
rect 81196 7496 81236 7792
rect 81292 7757 81332 7876
rect 81483 7916 81525 7925
rect 81483 7876 81484 7916
rect 81524 7876 81525 7916
rect 81483 7867 81525 7876
rect 81676 7916 81716 8035
rect 82059 8000 82101 8009
rect 82059 7960 82060 8000
rect 82100 7960 82101 8000
rect 82059 7951 82101 7960
rect 81676 7867 81716 7876
rect 81867 7916 81909 7925
rect 81867 7876 81868 7916
rect 81908 7876 81909 7916
rect 81867 7867 81909 7876
rect 82060 7916 82100 7951
rect 81387 7832 81429 7841
rect 81387 7792 81388 7832
rect 81428 7792 81429 7832
rect 81387 7783 81429 7792
rect 81291 7748 81333 7757
rect 81291 7708 81292 7748
rect 81332 7708 81333 7748
rect 81291 7699 81333 7708
rect 81196 7456 81332 7496
rect 81044 7204 81140 7244
rect 81004 7195 81044 7204
rect 81292 6749 81332 7456
rect 81291 6740 81333 6749
rect 81291 6700 81292 6740
rect 81332 6700 81333 6740
rect 81291 6691 81333 6700
rect 80908 6280 81236 6320
rect 80427 6271 80469 6280
rect 80428 5900 80468 6271
rect 80528 6068 80896 6077
rect 80568 6028 80610 6068
rect 80650 6028 80692 6068
rect 80732 6028 80774 6068
rect 80814 6028 80856 6068
rect 80528 6019 80896 6028
rect 81099 6068 81141 6077
rect 81099 6028 81100 6068
rect 81140 6028 81141 6068
rect 81099 6019 81141 6028
rect 80907 5900 80949 5909
rect 80428 5860 80564 5900
rect 80427 5732 80469 5741
rect 80427 5692 80428 5732
rect 80468 5692 80469 5732
rect 80427 5683 80469 5692
rect 80428 5598 80468 5683
rect 80276 4936 80372 4976
rect 80524 4976 80564 5860
rect 80907 5860 80908 5900
rect 80948 5860 80949 5900
rect 80907 5851 80949 5860
rect 80811 5816 80853 5825
rect 80811 5776 80812 5816
rect 80852 5776 80853 5816
rect 80811 5767 80853 5776
rect 80620 5732 80660 5743
rect 80620 5657 80660 5692
rect 80619 5648 80661 5657
rect 80619 5608 80620 5648
rect 80660 5608 80661 5648
rect 80619 5599 80661 5608
rect 80619 5480 80661 5489
rect 80619 5440 80620 5480
rect 80660 5440 80661 5480
rect 80619 5431 80661 5440
rect 80620 5346 80660 5431
rect 80812 5153 80852 5767
rect 80908 5741 80948 5851
rect 80907 5732 80949 5741
rect 81100 5732 81140 6019
rect 80907 5692 80908 5732
rect 80948 5692 80949 5732
rect 80907 5683 80949 5692
rect 81004 5692 81100 5732
rect 80908 5598 80948 5683
rect 80811 5144 80853 5153
rect 80811 5104 80812 5144
rect 80852 5104 80853 5144
rect 80811 5095 80853 5104
rect 80620 4976 80660 4985
rect 80524 4936 80620 4976
rect 80236 4927 80276 4936
rect 80620 4927 80660 4936
rect 80812 4892 80852 5095
rect 80907 4976 80949 4985
rect 80907 4936 80908 4976
rect 80948 4936 80949 4976
rect 80907 4927 80949 4936
rect 80812 4843 80852 4852
rect 80908 4842 80948 4927
rect 81004 4892 81044 5692
rect 81100 5683 81140 5692
rect 81100 5480 81140 5489
rect 81100 5321 81140 5440
rect 81099 5312 81141 5321
rect 81099 5272 81100 5312
rect 81140 5272 81141 5312
rect 81099 5263 81141 5272
rect 81196 5060 81236 6280
rect 81388 5909 81428 7783
rect 81484 7782 81524 7867
rect 81868 7782 81908 7867
rect 82060 7865 82100 7876
rect 81964 7832 82004 7841
rect 81964 6740 82004 7792
rect 82156 7076 82196 8035
rect 81868 6700 82004 6740
rect 82060 7036 82196 7076
rect 81772 6236 81812 6245
rect 81868 6236 81908 6700
rect 81963 6488 82005 6497
rect 81963 6448 81964 6488
rect 82004 6448 82005 6488
rect 81963 6439 82005 6448
rect 81964 6354 82004 6439
rect 81970 6236 82012 6245
rect 81868 6196 81971 6236
rect 82011 6196 82012 6236
rect 81387 5900 81429 5909
rect 81387 5860 81388 5900
rect 81428 5860 81429 5900
rect 81387 5851 81429 5860
rect 81292 5741 81332 5826
rect 81291 5732 81333 5741
rect 81291 5692 81292 5732
rect 81332 5692 81333 5732
rect 81291 5683 81333 5692
rect 81483 5732 81525 5741
rect 81483 5692 81484 5732
rect 81524 5692 81525 5732
rect 81483 5683 81525 5692
rect 81676 5732 81716 5741
rect 81387 5648 81429 5657
rect 81387 5608 81388 5648
rect 81428 5608 81429 5648
rect 81387 5599 81429 5608
rect 80428 4724 80468 4733
rect 80140 4087 80180 4096
rect 80236 4684 80428 4724
rect 79851 3968 79893 3977
rect 79660 3928 79796 3968
rect 79563 3919 79605 3928
rect 79288 3800 79656 3809
rect 79328 3760 79370 3800
rect 79410 3760 79452 3800
rect 79492 3760 79534 3800
rect 79574 3760 79616 3800
rect 79288 3751 79656 3760
rect 79756 3632 79796 3928
rect 79851 3928 79852 3968
rect 79892 3928 79893 3968
rect 79851 3919 79893 3928
rect 79948 3968 79988 3977
rect 79988 3928 80084 3968
rect 79948 3919 79988 3928
rect 79660 3592 79796 3632
rect 79275 3548 79317 3557
rect 79275 3508 79276 3548
rect 79316 3508 79317 3548
rect 79275 3499 79317 3508
rect 79179 3380 79221 3389
rect 79179 3340 79180 3380
rect 79220 3340 79221 3380
rect 79179 3331 79221 3340
rect 78892 3256 79028 3296
rect 78412 3212 78452 3221
rect 78412 2801 78452 3172
rect 78796 3212 78836 3221
rect 78411 2792 78453 2801
rect 78411 2752 78412 2792
rect 78452 2752 78453 2792
rect 78411 2743 78453 2752
rect 78124 2500 78356 2540
rect 78027 2372 78069 2381
rect 78124 2372 78164 2500
rect 78027 2332 78028 2372
rect 78068 2332 78164 2372
rect 78219 2372 78261 2381
rect 78219 2332 78220 2372
rect 78260 2332 78261 2372
rect 78027 2323 78069 2332
rect 78219 2323 78261 2332
rect 77932 1996 78068 2036
rect 77643 1112 77685 1121
rect 77643 1072 77644 1112
rect 77684 1072 77685 1112
rect 77643 1063 77685 1072
rect 77643 944 77685 953
rect 77643 904 77644 944
rect 77684 904 77685 944
rect 77643 895 77685 904
rect 77644 80 77684 895
rect 77835 776 77877 785
rect 77835 736 77836 776
rect 77876 736 77877 776
rect 77835 727 77877 736
rect 77836 80 77876 727
rect 78028 80 78068 1996
rect 78220 80 78260 2323
rect 78411 2288 78453 2297
rect 78411 2248 78412 2288
rect 78452 2248 78453 2288
rect 78411 2239 78453 2248
rect 78412 80 78452 2239
rect 78603 2204 78645 2213
rect 78603 2164 78604 2204
rect 78644 2164 78645 2204
rect 78603 2155 78645 2164
rect 78604 80 78644 2155
rect 78796 869 78836 3172
rect 78891 2792 78933 2801
rect 78891 2752 78892 2792
rect 78932 2752 78933 2792
rect 78891 2743 78933 2752
rect 78795 860 78837 869
rect 78795 820 78796 860
rect 78836 820 78837 860
rect 78795 811 78837 820
rect 78892 692 78932 2743
rect 78796 652 78932 692
rect 78796 80 78836 652
rect 78988 80 79028 3256
rect 79180 3212 79220 3221
rect 79180 1205 79220 3172
rect 79179 1196 79221 1205
rect 79179 1156 79180 1196
rect 79220 1156 79221 1196
rect 79179 1147 79221 1156
rect 79276 1028 79316 3499
rect 79371 3464 79413 3473
rect 79371 3424 79372 3464
rect 79412 3424 79413 3464
rect 79371 3415 79413 3424
rect 79372 3330 79412 3415
rect 79564 3212 79604 3221
rect 79564 2885 79604 3172
rect 79563 2876 79605 2885
rect 79563 2836 79564 2876
rect 79604 2836 79605 2876
rect 79563 2827 79605 2836
rect 79660 2381 79700 3592
rect 79756 3464 79796 3475
rect 79756 3389 79796 3424
rect 79755 3380 79797 3389
rect 79755 3340 79756 3380
rect 79796 3340 79797 3380
rect 79755 3331 79797 3340
rect 79852 3212 79892 3919
rect 79756 3172 79892 3212
rect 79948 3212 79988 3221
rect 79659 2372 79701 2381
rect 79659 2332 79660 2372
rect 79700 2332 79701 2372
rect 79659 2323 79701 2332
rect 79756 1289 79796 3172
rect 79948 2540 79988 3172
rect 79852 2500 79988 2540
rect 79755 1280 79797 1289
rect 79755 1240 79756 1280
rect 79796 1240 79797 1280
rect 79755 1231 79797 1240
rect 79563 1112 79605 1121
rect 79563 1072 79564 1112
rect 79604 1072 79605 1112
rect 79563 1063 79605 1072
rect 79180 988 79316 1028
rect 79180 80 79220 988
rect 79371 188 79413 197
rect 79371 148 79372 188
rect 79412 148 79413 188
rect 79371 139 79413 148
rect 79372 80 79412 139
rect 79564 80 79604 1063
rect 79852 1037 79892 2500
rect 79947 1280 79989 1289
rect 79947 1240 79948 1280
rect 79988 1240 79989 1280
rect 79947 1231 79989 1240
rect 79851 1028 79893 1037
rect 79851 988 79852 1028
rect 79892 988 79893 1028
rect 79851 979 79893 988
rect 79755 692 79797 701
rect 79755 652 79756 692
rect 79796 652 79797 692
rect 79755 643 79797 652
rect 79756 80 79796 643
rect 79948 80 79988 1231
rect 80044 785 80084 3928
rect 80139 3464 80181 3473
rect 80139 3424 80140 3464
rect 80180 3424 80181 3464
rect 80139 3415 80181 3424
rect 80140 3330 80180 3415
rect 80236 2213 80276 4684
rect 80428 4675 80468 4684
rect 80427 4556 80469 4565
rect 80427 4516 80428 4556
rect 80468 4516 80469 4556
rect 80427 4507 80469 4516
rect 80528 4556 80896 4565
rect 80568 4516 80610 4556
rect 80650 4516 80692 4556
rect 80732 4516 80774 4556
rect 80814 4516 80856 4556
rect 80528 4507 80896 4516
rect 80428 4388 80468 4507
rect 80907 4388 80949 4397
rect 80428 4348 80564 4388
rect 80427 4136 80469 4145
rect 80427 4096 80428 4136
rect 80468 4096 80469 4136
rect 80427 4087 80469 4096
rect 80524 4136 80564 4348
rect 80907 4348 80908 4388
rect 80948 4348 80949 4388
rect 80907 4339 80949 4348
rect 80619 4304 80661 4313
rect 80619 4264 80620 4304
rect 80660 4264 80661 4304
rect 80619 4255 80661 4264
rect 80524 4087 80564 4096
rect 80331 3968 80373 3977
rect 80331 3928 80332 3968
rect 80372 3928 80373 3968
rect 80331 3919 80373 3928
rect 80332 3834 80372 3919
rect 80332 3212 80372 3221
rect 80235 2204 80277 2213
rect 80235 2164 80236 2204
rect 80276 2164 80277 2204
rect 80235 2155 80277 2164
rect 80139 1196 80181 1205
rect 80139 1156 80140 1196
rect 80180 1156 80181 1196
rect 80139 1147 80181 1156
rect 80043 776 80085 785
rect 80043 736 80044 776
rect 80084 736 80085 776
rect 80043 727 80085 736
rect 80140 80 80180 1147
rect 80332 953 80372 3172
rect 80428 2297 80468 4087
rect 80620 3893 80660 4255
rect 80716 4220 80756 4229
rect 80619 3884 80661 3893
rect 80619 3844 80620 3884
rect 80660 3844 80661 3884
rect 80619 3835 80661 3844
rect 80716 3809 80756 4180
rect 80908 4220 80948 4339
rect 81004 4313 81044 4852
rect 81100 5020 81236 5060
rect 81003 4304 81045 4313
rect 81003 4264 81004 4304
rect 81044 4264 81045 4304
rect 81003 4255 81045 4264
rect 80908 4145 80948 4180
rect 80907 4136 80949 4145
rect 80907 4096 80908 4136
rect 80948 4096 80949 4136
rect 80907 4087 80949 4096
rect 80908 3968 80948 3977
rect 80948 3928 81044 3968
rect 80908 3919 80948 3928
rect 80715 3800 80757 3809
rect 80715 3760 80716 3800
rect 80756 3760 80757 3800
rect 80715 3751 80757 3760
rect 80523 3464 80565 3473
rect 80523 3424 80524 3464
rect 80564 3424 80565 3464
rect 80523 3415 80565 3424
rect 80524 3330 80564 3415
rect 80528 3044 80896 3053
rect 80568 3004 80610 3044
rect 80650 3004 80692 3044
rect 80732 3004 80774 3044
rect 80814 3004 80856 3044
rect 80528 2995 80896 3004
rect 80427 2288 80469 2297
rect 80427 2248 80428 2288
rect 80468 2248 80469 2288
rect 80427 2239 80469 2248
rect 81004 2129 81044 3928
rect 81100 3473 81140 5020
rect 81388 4905 81428 5599
rect 81484 5598 81524 5683
rect 81676 5489 81716 5692
rect 81484 5480 81524 5489
rect 81675 5480 81717 5489
rect 81524 5440 81620 5480
rect 81484 5431 81524 5440
rect 81483 5312 81525 5321
rect 81483 5272 81484 5312
rect 81524 5272 81525 5312
rect 81580 5312 81620 5440
rect 81675 5440 81676 5480
rect 81716 5440 81717 5480
rect 81675 5431 81717 5440
rect 81675 5312 81717 5321
rect 81580 5272 81676 5312
rect 81716 5272 81717 5312
rect 81483 5263 81525 5272
rect 81675 5263 81717 5272
rect 81196 4892 81236 4901
rect 81388 4856 81428 4865
rect 81196 3809 81236 4852
rect 81291 4724 81333 4733
rect 81291 4684 81292 4724
rect 81332 4684 81333 4724
rect 81291 4675 81333 4684
rect 81292 4590 81332 4675
rect 81484 4481 81524 5263
rect 81579 5144 81621 5153
rect 81579 5104 81580 5144
rect 81620 5104 81621 5144
rect 81579 5095 81621 5104
rect 81580 4892 81620 5095
rect 81772 5060 81812 6196
rect 81970 6187 82012 6196
rect 81963 6068 82005 6077
rect 81963 6028 81964 6068
rect 82004 6028 82005 6068
rect 81963 6019 82005 6028
rect 81868 5732 81908 5743
rect 81868 5657 81908 5692
rect 81867 5648 81909 5657
rect 81867 5608 81868 5648
rect 81908 5608 81909 5648
rect 81867 5599 81909 5608
rect 81867 5480 81909 5489
rect 81867 5440 81868 5480
rect 81908 5440 81909 5480
rect 81867 5431 81909 5440
rect 81868 5346 81908 5431
rect 81964 5153 82004 6019
rect 81963 5144 82005 5153
rect 81963 5104 81964 5144
rect 82004 5104 82005 5144
rect 81963 5095 82005 5104
rect 81772 5020 81908 5060
rect 81580 4843 81620 4852
rect 81771 4892 81813 4901
rect 81771 4852 81772 4892
rect 81812 4852 81813 4892
rect 81771 4843 81813 4852
rect 81772 4758 81812 4843
rect 81676 4724 81716 4733
rect 81483 4472 81525 4481
rect 81483 4432 81484 4472
rect 81524 4432 81525 4472
rect 81483 4423 81525 4432
rect 81579 4304 81621 4313
rect 81579 4264 81580 4304
rect 81620 4264 81621 4304
rect 81579 4255 81621 4264
rect 81291 4220 81333 4229
rect 81291 4180 81292 4220
rect 81332 4180 81333 4220
rect 81291 4171 81333 4180
rect 81292 4086 81332 4171
rect 81580 4052 81620 4255
rect 81580 4003 81620 4012
rect 81195 3800 81237 3809
rect 81195 3760 81196 3800
rect 81236 3760 81237 3800
rect 81195 3751 81237 3760
rect 81099 3464 81141 3473
rect 81099 3424 81100 3464
rect 81140 3424 81141 3464
rect 81099 3415 81141 3424
rect 81196 3380 81236 3389
rect 81099 3212 81141 3221
rect 81099 3172 81100 3212
rect 81140 3172 81141 3212
rect 81099 3163 81141 3172
rect 81003 2120 81045 2129
rect 81003 2080 81004 2120
rect 81044 2080 81045 2120
rect 81003 2071 81045 2080
rect 80907 1448 80949 1457
rect 80907 1408 80908 1448
rect 80948 1408 80949 1448
rect 80907 1399 80949 1408
rect 80523 1280 80565 1289
rect 80523 1240 80524 1280
rect 80564 1240 80565 1280
rect 80523 1231 80565 1240
rect 80331 944 80373 953
rect 80331 904 80332 944
rect 80372 904 80373 944
rect 80331 895 80373 904
rect 80331 776 80373 785
rect 80331 736 80332 776
rect 80372 736 80373 776
rect 80331 727 80373 736
rect 80332 80 80372 727
rect 80524 80 80564 1231
rect 80715 440 80757 449
rect 80715 400 80716 440
rect 80756 400 80757 440
rect 80715 391 80757 400
rect 80716 80 80756 391
rect 80908 80 80948 1399
rect 81100 80 81140 3163
rect 81196 2045 81236 3340
rect 81676 3305 81716 4684
rect 81771 4388 81813 4397
rect 81771 4348 81772 4388
rect 81812 4348 81813 4388
rect 81771 4339 81813 4348
rect 81772 3632 81812 4339
rect 81772 3583 81812 3592
rect 81675 3296 81717 3305
rect 81675 3256 81676 3296
rect 81716 3256 81717 3296
rect 81675 3247 81717 3256
rect 81868 2540 81908 5020
rect 81676 2500 81908 2540
rect 81964 4724 82004 4733
rect 81195 2036 81237 2045
rect 81195 1996 81196 2036
rect 81236 1996 81237 2036
rect 81195 1987 81237 1996
rect 81291 1952 81333 1961
rect 81291 1912 81292 1952
rect 81332 1912 81333 1952
rect 81291 1903 81333 1912
rect 81292 1373 81332 1903
rect 81483 1532 81525 1541
rect 81483 1492 81484 1532
rect 81524 1492 81525 1532
rect 81483 1483 81525 1492
rect 81291 1364 81333 1373
rect 81291 1324 81292 1364
rect 81332 1324 81333 1364
rect 81291 1315 81333 1324
rect 81291 1028 81333 1037
rect 81291 988 81292 1028
rect 81332 988 81333 1028
rect 81291 979 81333 988
rect 81292 80 81332 979
rect 81484 80 81524 1483
rect 81676 80 81716 2500
rect 81867 1700 81909 1709
rect 81867 1660 81868 1700
rect 81908 1660 81909 1700
rect 81867 1651 81909 1660
rect 81868 80 81908 1651
rect 81964 785 82004 4684
rect 82060 3473 82100 7036
rect 82155 6908 82197 6917
rect 82155 6868 82156 6908
rect 82196 6868 82197 6908
rect 82155 6859 82197 6868
rect 82156 6404 82196 6859
rect 82252 6665 82292 9220
rect 82347 8840 82389 8849
rect 82347 8800 82348 8840
rect 82388 8800 82389 8840
rect 82347 8791 82389 8800
rect 82348 6824 82388 8791
rect 82443 8588 82485 8597
rect 82443 8548 82444 8588
rect 82484 8548 82485 8588
rect 82443 8539 82485 8548
rect 82444 7939 82484 8539
rect 82636 8084 82676 9976
rect 82732 9521 82772 10051
rect 82731 9512 82773 9521
rect 82731 9472 82732 9512
rect 82772 9472 82773 9512
rect 82731 9463 82773 9472
rect 82828 8093 82868 10471
rect 83211 10352 83253 10361
rect 83211 10312 83212 10352
rect 83252 10312 83253 10352
rect 83211 10303 83253 10312
rect 84076 10352 84116 10471
rect 87147 10436 87189 10445
rect 87147 10396 87148 10436
rect 87188 10396 87189 10436
rect 87147 10387 87189 10396
rect 84076 10303 84116 10312
rect 83212 10268 83252 10303
rect 83212 10217 83252 10228
rect 83404 10268 83444 10277
rect 83404 10109 83444 10228
rect 83595 10268 83637 10277
rect 83595 10228 83596 10268
rect 83636 10228 83637 10268
rect 83595 10219 83637 10228
rect 83788 10268 83828 10277
rect 83596 10134 83636 10219
rect 83788 10109 83828 10228
rect 83980 10268 84020 10279
rect 83980 10193 84020 10228
rect 84172 10268 84212 10277
rect 83979 10184 84021 10193
rect 83979 10144 83980 10184
rect 84020 10144 84021 10184
rect 83979 10135 84021 10144
rect 83403 10100 83445 10109
rect 83403 10060 83404 10100
rect 83444 10060 83445 10100
rect 83403 10051 83445 10060
rect 83787 10100 83829 10109
rect 83787 10060 83788 10100
rect 83828 10060 83829 10100
rect 83787 10051 83829 10060
rect 83307 10016 83349 10025
rect 83307 9976 83308 10016
rect 83348 9976 83349 10016
rect 83307 9967 83349 9976
rect 83692 10016 83732 10025
rect 83308 9882 83348 9967
rect 83211 9680 83253 9689
rect 83211 9640 83212 9680
rect 83252 9640 83253 9680
rect 83211 9631 83253 9640
rect 83212 8840 83252 9631
rect 83595 9092 83637 9101
rect 83595 9052 83596 9092
rect 83636 9052 83637 9092
rect 83595 9043 83637 9052
rect 83212 8791 83252 8800
rect 83596 8840 83636 9043
rect 83692 8924 83732 9976
rect 83883 10016 83925 10025
rect 83883 9976 83884 10016
rect 83924 9976 83925 10016
rect 83883 9967 83925 9976
rect 83692 8884 83828 8924
rect 83596 8791 83636 8800
rect 83020 8756 83159 8769
rect 83020 8729 83116 8756
rect 83020 8681 83060 8729
rect 83156 8716 83159 8756
rect 83308 8756 83348 8765
rect 83116 8707 83156 8716
rect 83019 8672 83061 8681
rect 83019 8632 83020 8672
rect 83060 8632 83061 8672
rect 83019 8623 83061 8632
rect 83020 8093 83060 8623
rect 83308 8168 83348 8716
rect 83500 8756 83540 8767
rect 83500 8681 83540 8716
rect 83691 8756 83733 8765
rect 83691 8716 83692 8756
rect 83732 8716 83733 8756
rect 83691 8707 83733 8716
rect 83499 8672 83541 8681
rect 83499 8632 83500 8672
rect 83540 8632 83541 8672
rect 83499 8623 83541 8632
rect 83692 8622 83732 8707
rect 83403 8420 83445 8429
rect 83403 8380 83404 8420
rect 83444 8380 83445 8420
rect 83403 8371 83445 8380
rect 83116 8128 83348 8168
rect 82827 8084 82869 8093
rect 82636 8044 82772 8084
rect 82443 7876 82444 7925
rect 82484 7876 82485 7925
rect 82443 7867 82485 7876
rect 82636 7916 82676 7927
rect 82444 7775 82484 7867
rect 82636 7841 82676 7876
rect 82540 7832 82580 7841
rect 82348 6784 82484 6824
rect 82251 6656 82293 6665
rect 82251 6616 82252 6656
rect 82292 6616 82293 6656
rect 82251 6607 82293 6616
rect 82348 6581 82388 6666
rect 82347 6572 82389 6581
rect 82347 6532 82348 6572
rect 82388 6532 82389 6572
rect 82347 6523 82389 6532
rect 82251 6488 82293 6497
rect 82251 6448 82252 6488
rect 82292 6448 82293 6488
rect 82251 6439 82293 6448
rect 82156 5909 82196 6364
rect 82155 5900 82197 5909
rect 82155 5860 82156 5900
rect 82196 5860 82197 5900
rect 82155 5851 82197 5860
rect 82156 5732 82196 5741
rect 82156 5573 82196 5692
rect 82155 5564 82197 5573
rect 82155 5524 82156 5564
rect 82196 5524 82197 5564
rect 82155 5515 82197 5524
rect 82156 4976 82196 4985
rect 82156 4733 82196 4936
rect 82155 4724 82197 4733
rect 82155 4684 82156 4724
rect 82196 4684 82197 4724
rect 82155 4675 82197 4684
rect 82155 3968 82197 3977
rect 82155 3928 82156 3968
rect 82196 3928 82197 3968
rect 82155 3919 82197 3928
rect 82059 3464 82101 3473
rect 82059 3424 82060 3464
rect 82100 3424 82101 3464
rect 82059 3415 82101 3424
rect 82059 2372 82101 2381
rect 82059 2332 82060 2372
rect 82100 2332 82101 2372
rect 82059 2323 82101 2332
rect 82060 1709 82100 2323
rect 82059 1700 82101 1709
rect 82059 1660 82060 1700
rect 82100 1660 82101 1700
rect 82059 1651 82101 1660
rect 81963 776 82005 785
rect 81963 736 81964 776
rect 82004 736 82005 776
rect 81963 727 82005 736
rect 82156 701 82196 3919
rect 82252 3725 82292 6439
rect 82347 6404 82389 6413
rect 82347 6364 82348 6404
rect 82388 6364 82389 6404
rect 82347 6355 82389 6364
rect 82348 6270 82388 6355
rect 82347 5816 82389 5825
rect 82347 5776 82348 5816
rect 82388 5776 82389 5816
rect 82347 5767 82389 5776
rect 82348 5732 82388 5767
rect 82348 5681 82388 5692
rect 82347 5480 82389 5489
rect 82347 5440 82348 5480
rect 82388 5440 82389 5480
rect 82347 5431 82389 5440
rect 82348 5346 82388 5431
rect 82444 4733 82484 6784
rect 82540 5993 82580 7792
rect 82635 7832 82677 7841
rect 82635 7792 82636 7832
rect 82676 7792 82677 7832
rect 82635 7783 82677 7792
rect 82635 7244 82677 7253
rect 82635 7204 82636 7244
rect 82676 7204 82677 7244
rect 82635 7195 82677 7204
rect 82636 7110 82676 7195
rect 82732 6572 82772 8044
rect 82827 8044 82828 8084
rect 82868 8044 82869 8084
rect 82827 8035 82869 8044
rect 83019 8084 83061 8093
rect 83019 8044 83020 8084
rect 83060 8044 83061 8084
rect 83019 8035 83061 8044
rect 83116 8009 83156 8128
rect 83115 8000 83157 8009
rect 83115 7960 83116 8000
rect 83156 7960 83157 8000
rect 82827 7916 82869 7925
rect 82827 7876 82828 7916
rect 82868 7876 82869 7916
rect 82827 7867 82869 7876
rect 83020 7916 83060 7956
rect 83115 7951 83157 7960
rect 82828 7782 82868 7867
rect 83020 7841 83060 7876
rect 82924 7832 82964 7841
rect 82924 7589 82964 7792
rect 83019 7832 83061 7841
rect 83019 7792 83020 7832
rect 83060 7792 83061 7832
rect 83019 7783 83061 7792
rect 82923 7580 82965 7589
rect 82923 7540 82924 7580
rect 82964 7540 82965 7580
rect 82923 7531 82965 7540
rect 82828 7244 82868 7255
rect 83020 7253 83060 7783
rect 83116 7748 83156 7951
rect 83212 7925 83252 8010
rect 83404 7925 83444 8371
rect 83788 8336 83828 8884
rect 83500 8296 83828 8336
rect 83211 7916 83253 7925
rect 83211 7876 83212 7916
rect 83252 7876 83253 7916
rect 83211 7867 83253 7876
rect 83403 7916 83445 7925
rect 83403 7876 83404 7916
rect 83444 7876 83445 7916
rect 83403 7867 83445 7876
rect 83308 7832 83348 7841
rect 83116 7708 83252 7748
rect 82828 7169 82868 7204
rect 83019 7244 83061 7253
rect 83019 7204 83020 7244
rect 83060 7204 83061 7244
rect 83019 7195 83061 7204
rect 83212 7244 83252 7708
rect 83308 7673 83348 7792
rect 83404 7782 83444 7867
rect 83307 7664 83349 7673
rect 83307 7624 83308 7664
rect 83348 7624 83349 7664
rect 83307 7615 83349 7624
rect 83500 7412 83540 8296
rect 83595 8168 83637 8177
rect 83595 8128 83596 8168
rect 83636 8128 83637 8168
rect 83595 8119 83637 8128
rect 83692 8168 83732 8177
rect 83787 8168 83829 8177
rect 83732 8128 83788 8168
rect 83828 8128 83829 8168
rect 83692 8119 83732 8128
rect 83787 8119 83829 8128
rect 83212 7195 83252 7204
rect 83308 7372 83540 7412
rect 83596 7916 83636 8119
rect 83788 8009 83828 8040
rect 83787 8000 83829 8009
rect 83787 7960 83788 8000
rect 83828 7960 83829 8000
rect 83787 7951 83829 7960
rect 82827 7160 82869 7169
rect 82827 7120 82828 7160
rect 82868 7120 82869 7160
rect 82827 7111 82869 7120
rect 83020 7110 83060 7195
rect 82828 6992 82868 7001
rect 82923 6992 82965 7001
rect 82868 6952 82924 6992
rect 82964 6952 82965 6992
rect 82828 6943 82868 6952
rect 82923 6943 82965 6952
rect 83116 6992 83156 7001
rect 83116 6833 83156 6952
rect 82827 6824 82869 6833
rect 82827 6784 82828 6824
rect 82868 6784 82869 6824
rect 82827 6775 82869 6784
rect 83115 6824 83157 6833
rect 83308 6824 83348 7372
rect 83403 7244 83445 7253
rect 83403 7204 83404 7244
rect 83444 7204 83445 7244
rect 83403 7195 83445 7204
rect 83596 7244 83636 7876
rect 83788 7916 83828 7951
rect 83788 7589 83828 7876
rect 83787 7580 83829 7589
rect 83787 7540 83788 7580
rect 83828 7540 83829 7580
rect 83787 7531 83829 7540
rect 83596 7195 83636 7204
rect 83788 7244 83828 7531
rect 83884 7505 83924 9967
rect 83980 9521 84020 10135
rect 84172 10109 84212 10228
rect 84171 10100 84213 10109
rect 84171 10060 84172 10100
rect 84212 10060 84213 10100
rect 84171 10051 84213 10060
rect 83979 9512 84021 9521
rect 83979 9472 83980 9512
rect 84020 9472 84021 9512
rect 83979 9463 84021 9472
rect 83979 8840 84021 8849
rect 83979 8800 83980 8840
rect 84020 8800 84021 8840
rect 83979 8791 84021 8800
rect 83980 8588 84020 8791
rect 84076 8756 84116 8765
rect 84172 8756 84212 10051
rect 86859 9428 86901 9437
rect 86859 9388 86860 9428
rect 86900 9388 86901 9428
rect 86859 9379 86901 9388
rect 87148 9428 87188 10387
rect 88300 10352 88340 10471
rect 89643 10436 89685 10445
rect 89643 10396 89644 10436
rect 89684 10396 89685 10436
rect 89643 10387 89685 10396
rect 89931 10436 89973 10445
rect 89931 10396 89932 10436
rect 89972 10396 89973 10436
rect 89931 10387 89973 10396
rect 88300 10303 88340 10312
rect 89163 10352 89205 10361
rect 89163 10312 89164 10352
rect 89204 10312 89205 10352
rect 89163 10303 89205 10312
rect 87820 10268 87860 10277
rect 87724 10228 87820 10268
rect 87531 9596 87573 9605
rect 87531 9556 87532 9596
rect 87572 9556 87573 9596
rect 87531 9547 87573 9556
rect 87148 9379 87188 9388
rect 87340 9428 87380 9437
rect 87380 9388 87476 9428
rect 87340 9379 87380 9388
rect 86763 9344 86805 9353
rect 86763 9304 86764 9344
rect 86804 9304 86805 9344
rect 86763 9295 86805 9304
rect 85995 9260 86037 9269
rect 85995 9220 85996 9260
rect 86036 9220 86037 9260
rect 85995 9211 86037 9220
rect 85035 8924 85077 8933
rect 85035 8884 85036 8924
rect 85076 8884 85077 8924
rect 85035 8875 85077 8884
rect 84116 8716 84212 8756
rect 84268 8756 84308 8767
rect 84076 8707 84116 8716
rect 84268 8681 84308 8716
rect 84363 8756 84405 8765
rect 84363 8716 84364 8756
rect 84404 8716 84405 8756
rect 84363 8707 84405 8716
rect 84267 8672 84309 8681
rect 84267 8632 84268 8672
rect 84308 8632 84309 8672
rect 84267 8623 84309 8632
rect 84172 8588 84212 8597
rect 83980 8548 84172 8588
rect 84172 8539 84212 8548
rect 84267 8504 84309 8513
rect 84267 8464 84268 8504
rect 84308 8464 84309 8504
rect 84267 8455 84309 8464
rect 83979 7916 84021 7925
rect 83979 7876 83980 7916
rect 84020 7876 84021 7916
rect 83979 7867 84021 7876
rect 84171 7916 84213 7925
rect 84171 7876 84172 7916
rect 84212 7876 84213 7916
rect 84171 7867 84213 7876
rect 83980 7782 84020 7867
rect 84076 7832 84116 7841
rect 83979 7664 84021 7673
rect 83979 7624 83980 7664
rect 84020 7624 84021 7664
rect 83979 7615 84021 7624
rect 83883 7496 83925 7505
rect 83883 7456 83884 7496
rect 83924 7456 83925 7496
rect 83883 7447 83925 7456
rect 83788 7195 83828 7204
rect 83980 7244 84020 7615
rect 84076 7589 84116 7792
rect 84172 7782 84212 7867
rect 84171 7664 84213 7673
rect 84171 7624 84172 7664
rect 84212 7624 84213 7664
rect 84171 7615 84213 7624
rect 84075 7580 84117 7589
rect 84075 7540 84076 7580
rect 84116 7540 84117 7580
rect 84075 7531 84117 7540
rect 84172 7505 84212 7615
rect 84171 7496 84213 7505
rect 84171 7456 84172 7496
rect 84212 7456 84213 7496
rect 84171 7447 84213 7456
rect 83980 7195 84020 7204
rect 84172 7244 84212 7447
rect 84268 7244 84308 8455
rect 84364 7916 84404 8707
rect 84843 8000 84885 8009
rect 84843 7960 84844 8000
rect 84884 7960 84885 8000
rect 84843 7951 84885 7960
rect 84364 7867 84404 7876
rect 84555 7916 84597 7925
rect 84555 7876 84556 7916
rect 84596 7876 84597 7916
rect 84555 7867 84597 7876
rect 84748 7916 84788 7925
rect 84459 7832 84501 7841
rect 84459 7792 84460 7832
rect 84500 7792 84501 7832
rect 84459 7783 84501 7792
rect 84460 7698 84500 7783
rect 84556 7782 84596 7867
rect 84748 7757 84788 7876
rect 84844 7866 84884 7951
rect 84939 7916 84981 7925
rect 84939 7876 84940 7916
rect 84980 7876 84981 7916
rect 84939 7867 84981 7876
rect 84940 7757 84980 7867
rect 84747 7748 84789 7757
rect 84747 7708 84748 7748
rect 84788 7708 84789 7748
rect 84747 7699 84789 7708
rect 84939 7748 84981 7757
rect 84939 7708 84940 7748
rect 84980 7708 84981 7748
rect 84939 7699 84981 7708
rect 84364 7244 84404 7253
rect 84268 7204 84364 7244
rect 84172 7195 84212 7204
rect 84364 7195 84404 7204
rect 83404 7110 83444 7195
rect 84075 7160 84117 7169
rect 84075 7120 84076 7160
rect 84116 7120 84117 7160
rect 84075 7111 84117 7120
rect 83499 6992 83541 7001
rect 83499 6952 83500 6992
rect 83540 6952 83541 6992
rect 83499 6943 83541 6952
rect 83884 6992 83924 7001
rect 83500 6858 83540 6943
rect 83115 6784 83116 6824
rect 83156 6784 83157 6824
rect 83115 6775 83157 6784
rect 83212 6784 83348 6824
rect 83787 6824 83829 6833
rect 83787 6784 83788 6824
rect 83828 6784 83829 6824
rect 82636 6532 82772 6572
rect 82828 6572 82868 6775
rect 82828 6532 83060 6572
rect 82636 6329 82676 6532
rect 82828 6488 82868 6532
rect 82732 6448 82868 6488
rect 83020 6488 83060 6532
rect 83115 6488 83157 6497
rect 83020 6448 83116 6488
rect 83156 6448 83157 6488
rect 82732 6404 82772 6448
rect 83115 6439 83157 6448
rect 82732 6355 82772 6364
rect 82923 6404 82965 6413
rect 82923 6364 82924 6404
rect 82964 6364 82965 6404
rect 82923 6355 82965 6364
rect 83116 6404 83156 6439
rect 82635 6320 82677 6329
rect 82635 6280 82636 6320
rect 82676 6280 82677 6320
rect 82635 6271 82677 6280
rect 82827 6320 82869 6329
rect 82827 6280 82828 6320
rect 82868 6280 82869 6320
rect 82827 6271 82869 6280
rect 82828 6186 82868 6271
rect 82924 6270 82964 6355
rect 83116 6354 83156 6364
rect 83019 6320 83061 6329
rect 83019 6280 83020 6320
rect 83060 6280 83061 6320
rect 83019 6271 83061 6280
rect 83020 6068 83060 6271
rect 82732 6028 83060 6068
rect 82539 5984 82581 5993
rect 82539 5944 82540 5984
rect 82580 5944 82581 5984
rect 82539 5935 82581 5944
rect 82540 5732 82580 5741
rect 82540 5573 82580 5692
rect 82732 5732 82772 6028
rect 83115 5984 83157 5993
rect 83115 5944 83116 5984
rect 83156 5944 83157 5984
rect 83115 5935 83157 5944
rect 82923 5900 82965 5909
rect 82923 5860 82924 5900
rect 82964 5860 82965 5900
rect 82923 5851 82965 5860
rect 82827 5816 82869 5825
rect 82827 5776 82828 5816
rect 82868 5776 82869 5816
rect 82827 5767 82869 5776
rect 82635 5648 82677 5657
rect 82635 5608 82636 5648
rect 82676 5608 82677 5648
rect 82635 5599 82677 5608
rect 82539 5564 82581 5573
rect 82539 5524 82540 5564
rect 82580 5524 82581 5564
rect 82539 5515 82581 5524
rect 82636 5514 82676 5599
rect 82635 5228 82677 5237
rect 82635 5188 82636 5228
rect 82676 5188 82677 5228
rect 82635 5179 82677 5188
rect 82540 4976 82580 4985
rect 82348 4724 82388 4733
rect 82251 3716 82293 3725
rect 82251 3676 82252 3716
rect 82292 3676 82293 3716
rect 82251 3667 82293 3676
rect 82252 3212 82292 3221
rect 82252 2717 82292 3172
rect 82251 2708 82293 2717
rect 82251 2668 82252 2708
rect 82292 2668 82293 2708
rect 82251 2659 82293 2668
rect 82348 1457 82388 4684
rect 82443 4724 82485 4733
rect 82443 4684 82444 4724
rect 82484 4684 82485 4724
rect 82443 4675 82485 4684
rect 82540 4145 82580 4936
rect 82539 4136 82581 4145
rect 82539 4096 82540 4136
rect 82580 4096 82581 4136
rect 82539 4087 82581 4096
rect 82636 4136 82676 5179
rect 82732 5153 82772 5692
rect 82828 5564 82868 5767
rect 82924 5732 82964 5851
rect 83116 5732 83156 5935
rect 82924 5683 82964 5692
rect 83020 5692 83116 5732
rect 83020 5564 83060 5692
rect 83116 5683 83156 5692
rect 82828 5524 83060 5564
rect 82731 5144 82773 5153
rect 82731 5104 82732 5144
rect 82772 5104 82773 5144
rect 82731 5095 82773 5104
rect 82924 4901 82964 5524
rect 83116 5480 83156 5489
rect 83116 5237 83156 5440
rect 83115 5228 83157 5237
rect 83115 5188 83116 5228
rect 83156 5188 83157 5228
rect 83115 5179 83157 5188
rect 83019 5060 83061 5069
rect 83019 5020 83020 5060
rect 83060 5020 83061 5060
rect 83019 5011 83061 5020
rect 82732 4892 82772 4901
rect 82732 4565 82772 4852
rect 82923 4892 82965 4901
rect 82923 4852 82924 4892
rect 82964 4852 82965 4892
rect 82923 4843 82965 4852
rect 82828 4724 82868 4733
rect 82868 4684 82964 4724
rect 82828 4675 82868 4684
rect 82731 4556 82773 4565
rect 82731 4516 82732 4556
rect 82772 4516 82773 4556
rect 82731 4507 82773 4516
rect 82732 4145 82772 4507
rect 82636 4087 82676 4096
rect 82731 4136 82773 4145
rect 82731 4096 82732 4136
rect 82772 4096 82773 4136
rect 82731 4087 82773 4096
rect 82443 3968 82485 3977
rect 82828 3968 82868 3977
rect 82443 3928 82444 3968
rect 82484 3928 82485 3968
rect 82443 3919 82485 3928
rect 82732 3928 82828 3968
rect 82444 3834 82484 3919
rect 82443 3716 82485 3725
rect 82443 3676 82444 3716
rect 82484 3676 82485 3716
rect 82443 3667 82485 3676
rect 82444 3464 82484 3667
rect 82635 3548 82677 3557
rect 82635 3508 82636 3548
rect 82676 3508 82677 3548
rect 82635 3499 82677 3508
rect 82444 3415 82484 3424
rect 82636 3414 82676 3499
rect 82347 1448 82389 1457
rect 82347 1408 82348 1448
rect 82388 1408 82389 1448
rect 82347 1399 82389 1408
rect 82635 1448 82677 1457
rect 82635 1408 82636 1448
rect 82676 1408 82677 1448
rect 82635 1399 82677 1408
rect 82251 1364 82293 1373
rect 82251 1324 82252 1364
rect 82292 1324 82293 1364
rect 82251 1315 82293 1324
rect 82155 692 82197 701
rect 82155 652 82156 692
rect 82196 652 82197 692
rect 82155 643 82197 652
rect 82059 608 82101 617
rect 82059 568 82060 608
rect 82100 568 82101 608
rect 82059 559 82101 568
rect 82060 80 82100 559
rect 82252 80 82292 1315
rect 82443 860 82485 869
rect 82443 820 82444 860
rect 82484 820 82485 860
rect 82443 811 82485 820
rect 82444 80 82484 811
rect 82636 80 82676 1399
rect 82732 1289 82772 3928
rect 82828 3919 82868 3928
rect 82924 3557 82964 4684
rect 83020 4136 83060 5011
rect 83212 4388 83252 6784
rect 83787 6775 83829 6784
rect 83308 6581 83348 6666
rect 83307 6572 83349 6581
rect 83307 6532 83308 6572
rect 83348 6532 83349 6572
rect 83307 6523 83349 6532
rect 83403 6488 83445 6497
rect 83403 6448 83404 6488
rect 83444 6448 83445 6488
rect 83403 6439 83445 6448
rect 83595 6488 83637 6497
rect 83595 6448 83596 6488
rect 83636 6448 83637 6488
rect 83595 6439 83637 6448
rect 83308 6404 83348 6415
rect 83308 6329 83348 6364
rect 83307 6320 83349 6329
rect 83307 6280 83308 6320
rect 83348 6280 83349 6320
rect 83307 6271 83349 6280
rect 83307 6152 83349 6161
rect 83307 6112 83308 6152
rect 83348 6112 83349 6152
rect 83307 6103 83349 6112
rect 83308 5732 83348 6103
rect 83308 5683 83348 5692
rect 83308 4892 83348 4901
rect 83404 4892 83444 6439
rect 83500 6404 83540 6413
rect 83500 6161 83540 6364
rect 83596 6354 83636 6439
rect 83692 6404 83732 6415
rect 83692 6329 83732 6364
rect 83691 6320 83733 6329
rect 83691 6280 83692 6320
rect 83732 6280 83733 6320
rect 83691 6271 83733 6280
rect 83499 6152 83541 6161
rect 83499 6112 83500 6152
rect 83540 6112 83541 6152
rect 83499 6103 83541 6112
rect 83788 5984 83828 6775
rect 83884 6749 83924 6952
rect 83883 6740 83925 6749
rect 83883 6700 83884 6740
rect 83924 6700 83925 6740
rect 83883 6691 83925 6700
rect 83884 6404 83924 6413
rect 83884 6161 83924 6364
rect 84076 6404 84116 7111
rect 84651 7076 84693 7085
rect 84651 7036 84652 7076
rect 84692 7036 84693 7076
rect 84651 7027 84693 7036
rect 83979 6320 84021 6329
rect 83979 6280 83980 6320
rect 84020 6280 84021 6320
rect 83979 6271 84021 6280
rect 83980 6186 84020 6271
rect 83883 6152 83925 6161
rect 83883 6112 83884 6152
rect 83924 6112 83925 6152
rect 83883 6103 83925 6112
rect 84076 5993 84116 6364
rect 84268 6992 84308 7001
rect 84171 6068 84213 6077
rect 84171 6028 84172 6068
rect 84212 6028 84213 6068
rect 84171 6019 84213 6028
rect 84075 5984 84117 5993
rect 83788 5944 84020 5984
rect 83691 5900 83733 5909
rect 83691 5860 83692 5900
rect 83732 5860 83733 5900
rect 83691 5851 83733 5860
rect 83500 5732 83540 5741
rect 83692 5732 83732 5851
rect 83883 5816 83925 5825
rect 83883 5776 83884 5816
rect 83924 5776 83925 5816
rect 83883 5767 83925 5776
rect 83540 5692 83636 5732
rect 83500 5683 83540 5692
rect 83499 5480 83541 5489
rect 83499 5440 83500 5480
rect 83540 5440 83541 5480
rect 83499 5431 83541 5440
rect 83500 5346 83540 5431
rect 83348 4852 83444 4892
rect 83499 4892 83541 4901
rect 83499 4852 83500 4892
rect 83540 4852 83541 4892
rect 83596 4892 83636 5692
rect 83692 5683 83732 5692
rect 83787 5732 83829 5741
rect 83787 5692 83788 5732
rect 83828 5692 83829 5732
rect 83787 5683 83829 5692
rect 83884 5732 83924 5767
rect 83692 4892 83732 4901
rect 83596 4852 83692 4892
rect 83788 4892 83828 5683
rect 83884 5681 83924 5692
rect 83883 5564 83925 5573
rect 83883 5524 83884 5564
rect 83924 5524 83925 5564
rect 83883 5515 83925 5524
rect 83884 5430 83924 5515
rect 83980 5321 84020 5944
rect 84075 5944 84076 5984
rect 84116 5944 84117 5984
rect 84075 5935 84117 5944
rect 83979 5312 84021 5321
rect 83979 5272 83980 5312
rect 84020 5272 84021 5312
rect 83979 5263 84021 5272
rect 84075 5060 84117 5069
rect 84075 5020 84076 5060
rect 84116 5020 84117 5060
rect 84075 5011 84117 5020
rect 83884 4892 83924 4901
rect 83788 4852 83884 4892
rect 83924 4852 84020 4892
rect 83308 4843 83348 4852
rect 83499 4843 83541 4852
rect 83500 4758 83540 4843
rect 83403 4724 83445 4733
rect 83403 4684 83404 4724
rect 83444 4684 83445 4724
rect 83403 4675 83445 4684
rect 83404 4590 83444 4675
rect 83692 4397 83732 4852
rect 83884 4843 83924 4852
rect 83788 4724 83828 4733
rect 83788 4565 83828 4684
rect 83883 4724 83925 4733
rect 83883 4684 83884 4724
rect 83924 4684 83925 4724
rect 83883 4675 83925 4684
rect 83787 4556 83829 4565
rect 83787 4516 83788 4556
rect 83828 4516 83829 4556
rect 83787 4507 83829 4516
rect 83403 4388 83445 4397
rect 83212 4348 83348 4388
rect 83212 4220 83252 4229
rect 83212 4145 83252 4180
rect 83020 4087 83060 4096
rect 83211 4136 83253 4145
rect 83211 4096 83212 4136
rect 83252 4096 83253 4136
rect 83211 4087 83253 4096
rect 83212 3641 83252 4087
rect 83211 3632 83253 3641
rect 83211 3592 83212 3632
rect 83252 3592 83253 3632
rect 83211 3583 83253 3592
rect 82923 3548 82965 3557
rect 82923 3508 82924 3548
rect 82964 3508 82965 3548
rect 82923 3499 82965 3508
rect 82827 3464 82869 3473
rect 82827 3424 82828 3464
rect 82868 3424 82869 3464
rect 82827 3415 82869 3424
rect 83212 3464 83252 3473
rect 83308 3464 83348 4348
rect 83403 4348 83404 4388
rect 83444 4348 83445 4388
rect 83403 4339 83445 4348
rect 83691 4388 83733 4397
rect 83691 4348 83692 4388
rect 83732 4348 83733 4388
rect 83691 4339 83733 4348
rect 83404 4220 83444 4339
rect 83404 4171 83444 4180
rect 83788 4136 83828 4145
rect 83692 4096 83788 4136
rect 83404 3968 83444 3977
rect 83596 3968 83636 3977
rect 83404 3725 83444 3928
rect 83500 3928 83596 3968
rect 83403 3716 83445 3725
rect 83403 3676 83404 3716
rect 83444 3676 83445 3716
rect 83403 3667 83445 3676
rect 83252 3424 83348 3464
rect 83212 3415 83252 3424
rect 82828 3330 82868 3415
rect 83020 3212 83060 3221
rect 83020 2540 83060 3172
rect 82924 2500 83060 2540
rect 83404 3212 83444 3221
rect 82731 1280 82773 1289
rect 82731 1240 82732 1280
rect 82772 1240 82773 1280
rect 82731 1231 82773 1240
rect 82924 1121 82964 2500
rect 83307 2036 83349 2045
rect 83307 1996 83308 2036
rect 83348 1996 83349 2036
rect 83307 1987 83349 1996
rect 83019 1616 83061 1625
rect 83019 1576 83020 1616
rect 83060 1576 83061 1616
rect 83019 1567 83061 1576
rect 82923 1112 82965 1121
rect 82923 1072 82924 1112
rect 82964 1072 82965 1112
rect 82923 1063 82965 1072
rect 82827 272 82869 281
rect 82827 232 82828 272
rect 82868 232 82869 272
rect 82827 223 82869 232
rect 82828 80 82868 223
rect 83020 80 83060 1567
rect 83211 1112 83253 1121
rect 83211 1072 83212 1112
rect 83252 1072 83253 1112
rect 83211 1063 83253 1072
rect 83212 80 83252 1063
rect 83308 1028 83348 1987
rect 83404 1205 83444 3172
rect 83403 1196 83445 1205
rect 83403 1156 83404 1196
rect 83444 1156 83445 1196
rect 83403 1147 83445 1156
rect 83500 1037 83540 3928
rect 83596 3919 83636 3928
rect 83595 3800 83637 3809
rect 83595 3760 83596 3800
rect 83636 3760 83637 3800
rect 83595 3751 83637 3760
rect 83596 3464 83636 3751
rect 83596 3415 83636 3424
rect 83692 2213 83732 4096
rect 83788 4087 83828 4096
rect 83884 3473 83924 4675
rect 83980 4313 84020 4852
rect 84076 4565 84116 5011
rect 84075 4556 84117 4565
rect 84075 4516 84076 4556
rect 84116 4516 84117 4556
rect 84075 4507 84117 4516
rect 83979 4304 84021 4313
rect 83979 4264 83980 4304
rect 84020 4264 84021 4304
rect 83979 4255 84021 4264
rect 83883 3464 83925 3473
rect 83883 3424 83884 3464
rect 83924 3424 83925 3464
rect 83883 3415 83925 3424
rect 83980 3464 84020 3473
rect 84172 3464 84212 6019
rect 84268 5153 84308 6952
rect 84652 6404 84692 7027
rect 84556 6236 84596 6245
rect 84460 6196 84556 6236
rect 84363 5732 84405 5741
rect 84460 5732 84500 6196
rect 84556 6187 84596 6196
rect 84363 5692 84364 5732
rect 84404 5692 84500 5732
rect 84556 5732 84596 5741
rect 84652 5732 84692 6364
rect 84843 6320 84885 6329
rect 84843 6280 84844 6320
rect 84884 6280 84885 6320
rect 84843 6271 84885 6280
rect 84844 6186 84884 6271
rect 85036 6068 85076 8875
rect 85131 8504 85173 8513
rect 85131 8464 85132 8504
rect 85172 8464 85173 8504
rect 85131 8455 85173 8464
rect 85132 7916 85172 8455
rect 85899 8336 85941 8345
rect 85899 8296 85900 8336
rect 85940 8296 85941 8336
rect 85899 8287 85941 8296
rect 85227 8084 85269 8093
rect 85227 8044 85228 8084
rect 85268 8044 85269 8084
rect 85227 8035 85269 8044
rect 85228 7950 85268 8035
rect 85132 7867 85172 7876
rect 85324 7916 85364 7925
rect 85324 7757 85364 7876
rect 85323 7748 85365 7757
rect 85323 7708 85324 7748
rect 85364 7708 85365 7748
rect 85323 7699 85365 7708
rect 85515 7412 85557 7421
rect 85707 7412 85749 7421
rect 85515 7372 85516 7412
rect 85556 7372 85652 7412
rect 85515 7363 85557 7372
rect 85612 7253 85652 7372
rect 85707 7372 85708 7412
rect 85748 7372 85749 7412
rect 85707 7363 85749 7372
rect 85708 7328 85748 7363
rect 85708 7277 85748 7288
rect 85611 7244 85653 7253
rect 85611 7204 85612 7244
rect 85652 7204 85653 7244
rect 85611 7195 85653 7204
rect 85804 7244 85844 7253
rect 85612 7110 85652 7195
rect 85707 7160 85749 7169
rect 85707 7120 85708 7160
rect 85748 7120 85749 7160
rect 85707 7111 85749 7120
rect 85419 6572 85461 6581
rect 85419 6532 85420 6572
rect 85460 6532 85461 6572
rect 85419 6523 85461 6532
rect 85323 6488 85365 6497
rect 85323 6448 85324 6488
rect 85364 6448 85365 6488
rect 85323 6439 85365 6448
rect 84596 5692 84692 5732
rect 84748 6028 85076 6068
rect 84363 5683 84405 5692
rect 84556 5683 84596 5692
rect 84364 5648 84404 5683
rect 84364 5597 84404 5608
rect 84556 5480 84596 5489
rect 84363 5312 84405 5321
rect 84363 5272 84364 5312
rect 84404 5272 84405 5312
rect 84363 5263 84405 5272
rect 84267 5144 84309 5153
rect 84267 5104 84268 5144
rect 84308 5104 84309 5144
rect 84267 5095 84309 5104
rect 84267 4892 84309 4901
rect 84267 4852 84268 4892
rect 84308 4852 84309 4892
rect 84267 4843 84309 4852
rect 84268 4733 84308 4843
rect 84267 4724 84309 4733
rect 84267 4684 84268 4724
rect 84308 4684 84309 4724
rect 84267 4675 84309 4684
rect 84267 4556 84309 4565
rect 84267 4516 84268 4556
rect 84308 4516 84309 4556
rect 84267 4507 84309 4516
rect 84268 4220 84308 4507
rect 84268 4171 84308 4180
rect 84364 4145 84404 5263
rect 84556 4892 84596 5440
rect 84556 4565 84596 4852
rect 84651 4892 84693 4901
rect 84651 4852 84652 4892
rect 84692 4852 84693 4892
rect 84651 4843 84693 4852
rect 84555 4556 84597 4565
rect 84555 4516 84556 4556
rect 84596 4516 84597 4556
rect 84555 4507 84597 4516
rect 84459 4220 84501 4229
rect 84459 4180 84460 4220
rect 84500 4180 84501 4220
rect 84459 4171 84501 4180
rect 84363 4136 84405 4145
rect 84363 4096 84364 4136
rect 84404 4096 84405 4136
rect 84363 4087 84405 4096
rect 84460 4052 84500 4171
rect 84460 4003 84500 4012
rect 84363 3968 84405 3977
rect 84363 3928 84364 3968
rect 84404 3928 84405 3968
rect 84363 3919 84405 3928
rect 84020 3424 84212 3464
rect 84364 3464 84404 3919
rect 84459 3800 84501 3809
rect 84459 3760 84460 3800
rect 84500 3760 84501 3800
rect 84459 3751 84501 3760
rect 83980 3415 84020 3424
rect 84364 3415 84404 3424
rect 83788 3212 83828 3221
rect 83691 2204 83733 2213
rect 83691 2164 83692 2204
rect 83732 2164 83733 2204
rect 83691 2155 83733 2164
rect 83499 1028 83541 1037
rect 83308 988 83444 1028
rect 83404 80 83444 988
rect 83499 988 83500 1028
rect 83540 988 83541 1028
rect 83499 979 83541 988
rect 83595 776 83637 785
rect 83595 736 83596 776
rect 83636 736 83637 776
rect 83595 727 83637 736
rect 83596 80 83636 727
rect 83788 692 83828 3172
rect 84171 3212 84213 3221
rect 84171 3172 84172 3212
rect 84212 3172 84213 3212
rect 84171 3163 84213 3172
rect 84172 3078 84212 3163
rect 83979 1280 84021 1289
rect 84460 1280 84500 3751
rect 84556 3212 84596 3221
rect 84556 1541 84596 3172
rect 84652 2540 84692 4843
rect 84748 3464 84788 6028
rect 85131 5900 85173 5909
rect 85131 5860 85132 5900
rect 85172 5860 85173 5900
rect 85131 5851 85173 5860
rect 85036 5648 85076 5657
rect 84748 3415 84788 3424
rect 84844 5480 84884 5489
rect 84652 2500 84788 2540
rect 84555 1532 84597 1541
rect 84555 1492 84556 1532
rect 84596 1492 84597 1532
rect 84555 1483 84597 1492
rect 83979 1240 83980 1280
rect 84020 1240 84021 1280
rect 83979 1231 84021 1240
rect 84364 1240 84500 1280
rect 83692 652 83828 692
rect 83692 449 83732 652
rect 83787 524 83829 533
rect 83787 484 83788 524
rect 83828 484 83829 524
rect 83787 475 83829 484
rect 83691 440 83733 449
rect 83691 400 83692 440
rect 83732 400 83733 440
rect 83691 391 83733 400
rect 83788 80 83828 475
rect 83980 80 84020 1231
rect 84171 1196 84213 1205
rect 84171 1156 84172 1196
rect 84212 1156 84213 1196
rect 84171 1147 84213 1156
rect 84172 80 84212 1147
rect 84364 80 84404 1240
rect 84555 692 84597 701
rect 84555 652 84556 692
rect 84596 652 84597 692
rect 84555 643 84597 652
rect 84556 80 84596 643
rect 84748 80 84788 2500
rect 84844 1121 84884 5440
rect 85036 4817 85076 5608
rect 85035 4808 85077 4817
rect 85035 4768 85036 4808
rect 85076 4768 85077 4808
rect 85035 4759 85077 4768
rect 84939 4724 84981 4733
rect 84939 4684 84940 4724
rect 84980 4684 84981 4724
rect 84939 4675 84981 4684
rect 84940 4590 84980 4675
rect 85132 4061 85172 5851
rect 85228 5480 85268 5489
rect 85131 4052 85173 4061
rect 85131 4012 85132 4052
rect 85172 4012 85173 4052
rect 85131 4003 85173 4012
rect 85035 3968 85077 3977
rect 85035 3928 85036 3968
rect 85076 3928 85077 3968
rect 85035 3919 85077 3928
rect 84939 3632 84981 3641
rect 84939 3592 84940 3632
rect 84980 3592 84981 3632
rect 84939 3583 84981 3592
rect 84940 3380 84980 3583
rect 84940 3331 84980 3340
rect 85036 2540 85076 3919
rect 85131 3632 85173 3641
rect 85131 3592 85132 3632
rect 85172 3592 85173 3632
rect 85131 3583 85173 3592
rect 85132 3498 85172 3583
rect 85131 3380 85173 3389
rect 85131 3340 85132 3380
rect 85172 3340 85173 3380
rect 85131 3331 85173 3340
rect 85132 3246 85172 3331
rect 85036 2500 85172 2540
rect 84939 2456 84981 2465
rect 84939 2416 84940 2456
rect 84980 2416 84981 2456
rect 84939 2407 84981 2416
rect 84843 1112 84885 1121
rect 84843 1072 84844 1112
rect 84884 1072 84885 1112
rect 84843 1063 84885 1072
rect 84940 80 84980 2407
rect 85132 80 85172 2500
rect 85228 1289 85268 5440
rect 85324 5069 85364 6439
rect 85420 5648 85460 6523
rect 85515 5816 85557 5825
rect 85515 5776 85516 5816
rect 85556 5776 85557 5816
rect 85515 5767 85557 5776
rect 85420 5599 85460 5608
rect 85323 5060 85365 5069
rect 85323 5020 85324 5060
rect 85364 5020 85365 5060
rect 85323 5011 85365 5020
rect 85419 4556 85461 4565
rect 85419 4516 85420 4556
rect 85460 4516 85461 4556
rect 85419 4507 85461 4516
rect 85420 4388 85460 4507
rect 85420 4339 85460 4348
rect 85323 4304 85365 4313
rect 85323 4264 85324 4304
rect 85364 4264 85365 4304
rect 85323 4255 85365 4264
rect 85324 4220 85364 4255
rect 85516 4220 85556 5767
rect 85612 5480 85652 5489
rect 85612 4901 85652 5440
rect 85611 4892 85653 4901
rect 85611 4852 85612 4892
rect 85652 4852 85653 4892
rect 85611 4843 85653 4852
rect 85324 4169 85364 4180
rect 85420 4180 85516 4220
rect 85420 3389 85460 4180
rect 85516 4171 85556 4180
rect 85612 4724 85652 4733
rect 85515 4052 85557 4061
rect 85515 4012 85516 4052
rect 85556 4012 85557 4052
rect 85515 4003 85557 4012
rect 85516 3464 85556 4003
rect 85516 3415 85556 3424
rect 85419 3380 85461 3389
rect 85419 3340 85420 3380
rect 85460 3340 85461 3380
rect 85419 3331 85461 3340
rect 85324 3212 85364 3221
rect 85324 2381 85364 3172
rect 85612 2540 85652 4684
rect 85708 4313 85748 7111
rect 85804 7085 85844 7204
rect 85803 7076 85845 7085
rect 85803 7036 85804 7076
rect 85844 7036 85845 7076
rect 85803 7027 85845 7036
rect 85804 5648 85844 5659
rect 85804 5573 85844 5608
rect 85803 5564 85845 5573
rect 85803 5524 85804 5564
rect 85844 5524 85845 5564
rect 85803 5515 85845 5524
rect 85804 4976 85844 4985
rect 85900 4976 85940 8287
rect 85996 7169 86036 9211
rect 86091 9008 86133 9017
rect 86091 8968 86092 9008
rect 86132 8968 86133 9008
rect 86091 8959 86133 8968
rect 85995 7160 86037 7169
rect 85995 7120 85996 7160
rect 86036 7120 86037 7160
rect 85995 7111 86037 7120
rect 85844 4936 85940 4976
rect 85996 5480 86036 5489
rect 85804 4927 85844 4936
rect 85996 4901 86036 5440
rect 85995 4892 86037 4901
rect 85995 4852 85996 4892
rect 86036 4852 86037 4892
rect 85995 4843 86037 4852
rect 85803 4724 85845 4733
rect 85803 4684 85804 4724
rect 85844 4684 85845 4724
rect 85803 4675 85845 4684
rect 85996 4724 86036 4733
rect 85707 4304 85749 4313
rect 85707 4264 85708 4304
rect 85748 4264 85749 4304
rect 85707 4255 85749 4264
rect 85708 3968 85748 3977
rect 85708 3389 85748 3928
rect 85707 3380 85749 3389
rect 85707 3340 85708 3380
rect 85748 3340 85749 3380
rect 85707 3331 85749 3340
rect 85516 2500 85652 2540
rect 85708 3212 85748 3221
rect 85323 2372 85365 2381
rect 85323 2332 85324 2372
rect 85364 2332 85365 2372
rect 85323 2323 85365 2332
rect 85516 2045 85556 2500
rect 85515 2036 85557 2045
rect 85515 1996 85516 2036
rect 85556 1996 85557 2036
rect 85515 1987 85557 1996
rect 85708 1364 85748 3172
rect 85612 1324 85748 1364
rect 85227 1280 85269 1289
rect 85227 1240 85228 1280
rect 85268 1240 85269 1280
rect 85227 1231 85269 1240
rect 85515 1280 85557 1289
rect 85515 1240 85516 1280
rect 85556 1240 85557 1280
rect 85515 1231 85557 1240
rect 85323 1028 85365 1037
rect 85323 988 85324 1028
rect 85364 988 85365 1028
rect 85323 979 85365 988
rect 85324 80 85364 979
rect 85516 80 85556 1231
rect 85612 617 85652 1324
rect 85804 1112 85844 4675
rect 85900 4136 85940 4145
rect 85900 3893 85940 4096
rect 85899 3884 85941 3893
rect 85899 3844 85900 3884
rect 85940 3844 85941 3884
rect 85899 3835 85941 3844
rect 85900 3464 85940 3473
rect 85900 2549 85940 3424
rect 85996 2633 86036 4684
rect 86092 4220 86132 8959
rect 86764 8504 86804 9295
rect 86860 8765 86900 9379
rect 87051 9344 87093 9353
rect 87051 9304 87052 9344
rect 87092 9304 87093 9344
rect 87051 9295 87093 9304
rect 87244 9344 87284 9353
rect 86955 8924 86997 8933
rect 86955 8884 86956 8924
rect 86996 8884 86997 8924
rect 86955 8875 86997 8884
rect 86956 8840 86996 8875
rect 86956 8789 86996 8800
rect 86859 8756 86901 8765
rect 86859 8716 86860 8756
rect 86900 8716 86901 8756
rect 86859 8707 86901 8716
rect 87052 8756 87092 9295
rect 87244 8924 87284 9304
rect 86860 8622 86900 8707
rect 86764 8464 86900 8504
rect 86860 8000 86900 8464
rect 86956 8168 86996 8177
rect 87052 8168 87092 8716
rect 86996 8128 87092 8168
rect 87148 8884 87284 8924
rect 86956 8119 86996 8128
rect 86860 7960 87092 8000
rect 86764 7916 86804 7925
rect 86804 7876 86900 7916
rect 86764 7867 86804 7876
rect 86860 7757 86900 7876
rect 86859 7748 86901 7757
rect 86859 7708 86860 7748
rect 86900 7708 86901 7748
rect 86859 7699 86901 7708
rect 86860 7412 86900 7699
rect 86860 7363 86900 7372
rect 86379 7244 86421 7253
rect 86379 7204 86380 7244
rect 86420 7204 86421 7244
rect 86379 7195 86421 7204
rect 86283 7160 86325 7169
rect 86283 7120 86284 7160
rect 86324 7120 86325 7160
rect 86283 7111 86325 7120
rect 86187 5648 86229 5657
rect 86187 5608 86188 5648
rect 86228 5608 86229 5648
rect 86187 5599 86229 5608
rect 86188 5514 86228 5599
rect 86188 4976 86228 4985
rect 86284 4976 86324 7111
rect 86380 7110 86420 7195
rect 86859 7076 86901 7085
rect 86859 7036 86860 7076
rect 86900 7036 86901 7076
rect 86859 7027 86901 7036
rect 86571 6992 86613 7001
rect 86571 6952 86572 6992
rect 86612 6952 86613 6992
rect 86571 6943 86613 6952
rect 86475 6572 86517 6581
rect 86475 6532 86476 6572
rect 86516 6532 86517 6572
rect 86475 6523 86517 6532
rect 86476 5564 86516 6523
rect 86572 5825 86612 6943
rect 86668 6404 86708 6415
rect 86668 6329 86708 6364
rect 86860 6404 86900 7027
rect 86860 6355 86900 6364
rect 86667 6320 86709 6329
rect 86667 6280 86668 6320
rect 86708 6280 86709 6320
rect 86667 6271 86709 6280
rect 86764 6320 86804 6329
rect 86571 5816 86613 5825
rect 86571 5776 86572 5816
rect 86612 5776 86613 5816
rect 86571 5767 86613 5776
rect 86590 5661 86630 5670
rect 86630 5621 86708 5648
rect 86590 5608 86708 5621
rect 86476 5524 86612 5564
rect 86380 5480 86420 5489
rect 86420 5440 86516 5480
rect 86380 5431 86420 5440
rect 86228 4936 86324 4976
rect 86188 4927 86228 4936
rect 86380 4724 86420 4733
rect 86380 4397 86420 4684
rect 86379 4388 86421 4397
rect 86379 4348 86380 4388
rect 86420 4348 86421 4388
rect 86379 4339 86421 4348
rect 86092 4180 86228 4220
rect 86188 4136 86228 4180
rect 86283 4136 86325 4145
rect 86476 4136 86516 5440
rect 86572 4976 86612 5524
rect 86572 4927 86612 4936
rect 86571 4640 86613 4649
rect 86571 4600 86572 4640
rect 86612 4600 86613 4640
rect 86571 4591 86613 4600
rect 86188 4096 86238 4136
rect 86092 4052 86132 4061
rect 86092 3389 86132 4012
rect 86198 3968 86238 4096
rect 86283 4096 86284 4136
rect 86324 4096 86325 4136
rect 86283 4087 86325 4096
rect 86380 4096 86516 4136
rect 86572 4136 86612 4591
rect 86668 4565 86708 5608
rect 86764 4892 86804 6280
rect 86955 5060 86997 5069
rect 86955 5020 86956 5060
rect 86996 5020 86997 5060
rect 86955 5011 86997 5020
rect 86956 4976 86996 5011
rect 87052 4985 87092 7960
rect 87148 7916 87188 8884
rect 87436 8849 87476 9388
rect 87435 8840 87477 8849
rect 87435 8800 87436 8840
rect 87476 8800 87477 8840
rect 87435 8791 87477 8800
rect 87244 8756 87284 8767
rect 87244 8681 87284 8716
rect 87436 8756 87476 8791
rect 87436 8705 87476 8716
rect 87532 8681 87572 9547
rect 87724 9428 87764 10228
rect 87820 10219 87860 10228
rect 88011 10268 88053 10277
rect 88011 10228 88012 10268
rect 88052 10228 88053 10268
rect 88011 10219 88053 10228
rect 88204 10268 88244 10279
rect 88012 10134 88052 10219
rect 88204 10193 88244 10228
rect 88395 10268 88437 10277
rect 88588 10268 88628 10277
rect 88395 10228 88396 10268
rect 88436 10228 88532 10268
rect 88395 10219 88437 10228
rect 88203 10184 88245 10193
rect 88203 10144 88204 10184
rect 88244 10144 88245 10184
rect 88203 10135 88245 10144
rect 88396 10134 88436 10219
rect 87915 10100 87957 10109
rect 87915 10060 87916 10100
rect 87956 10060 87957 10100
rect 87915 10051 87957 10060
rect 87916 9966 87956 10051
rect 88107 9764 88149 9773
rect 88107 9724 88108 9764
rect 88148 9724 88149 9764
rect 88107 9715 88149 9724
rect 87915 9512 87957 9521
rect 87915 9472 87916 9512
rect 87956 9472 87957 9512
rect 87915 9463 87957 9472
rect 87724 9353 87764 9388
rect 87819 9428 87861 9437
rect 87819 9388 87820 9428
rect 87860 9388 87861 9428
rect 87819 9379 87861 9388
rect 87916 9428 87956 9463
rect 87723 9344 87765 9353
rect 87723 9304 87724 9344
rect 87764 9304 87765 9344
rect 87723 9295 87765 9304
rect 87820 9294 87860 9379
rect 87916 9377 87956 9388
rect 87723 9008 87765 9017
rect 87723 8968 87724 9008
rect 87764 8968 87765 9008
rect 87723 8959 87765 8968
rect 87724 8840 87764 8959
rect 87724 8791 87764 8800
rect 87915 8840 87957 8849
rect 87915 8800 87916 8840
rect 87956 8800 87957 8840
rect 87915 8791 87957 8800
rect 87627 8756 87669 8765
rect 87627 8716 87628 8756
rect 87668 8716 87669 8756
rect 87627 8707 87669 8716
rect 87820 8756 87860 8765
rect 87243 8672 87285 8681
rect 87243 8632 87244 8672
rect 87284 8632 87285 8672
rect 87243 8623 87285 8632
rect 87531 8672 87573 8681
rect 87531 8632 87532 8672
rect 87572 8632 87573 8672
rect 87531 8623 87573 8632
rect 87628 8622 87668 8707
rect 87820 8672 87860 8716
rect 87724 8632 87860 8672
rect 87340 8504 87380 8513
rect 87148 7876 87284 7916
rect 86956 4925 86996 4936
rect 87051 4976 87093 4985
rect 87051 4936 87052 4976
rect 87092 4936 87093 4976
rect 87051 4927 87093 4936
rect 86764 4852 86900 4892
rect 86763 4724 86805 4733
rect 86763 4684 86764 4724
rect 86804 4684 86805 4724
rect 86763 4675 86805 4684
rect 86764 4590 86804 4675
rect 86860 4565 86900 4852
rect 87148 4724 87188 4733
rect 86956 4684 87148 4724
rect 86667 4556 86709 4565
rect 86667 4516 86668 4556
rect 86708 4516 86709 4556
rect 86667 4507 86709 4516
rect 86859 4556 86901 4565
rect 86859 4516 86860 4556
rect 86900 4516 86901 4556
rect 86859 4507 86901 4516
rect 86763 4304 86805 4313
rect 86763 4264 86764 4304
rect 86804 4264 86805 4304
rect 86763 4255 86805 4264
rect 86668 4136 86708 4145
rect 86572 4096 86668 4136
rect 86284 4002 86324 4087
rect 86188 3928 86238 3968
rect 86188 3464 86228 3928
rect 86284 3464 86324 3473
rect 86188 3424 86284 3464
rect 86284 3415 86324 3424
rect 86091 3380 86133 3389
rect 86091 3340 86092 3380
rect 86132 3340 86133 3380
rect 86091 3331 86133 3340
rect 86092 3212 86132 3221
rect 85995 2624 86037 2633
rect 85995 2584 85996 2624
rect 86036 2584 86037 2624
rect 85995 2575 86037 2584
rect 85899 2540 85941 2549
rect 85899 2500 85900 2540
rect 85940 2500 85941 2540
rect 86092 2540 86132 3172
rect 86380 2540 86420 4096
rect 86668 4087 86708 4096
rect 86476 3968 86516 3977
rect 86516 3928 86612 3968
rect 86476 3919 86516 3928
rect 86092 2500 86228 2540
rect 85899 2491 85941 2500
rect 85899 2372 85941 2381
rect 85899 2332 85900 2372
rect 85940 2332 85941 2372
rect 85899 2323 85941 2332
rect 85708 1072 85844 1112
rect 85611 608 85653 617
rect 85611 568 85612 608
rect 85652 568 85653 608
rect 85611 559 85653 568
rect 85708 80 85748 1072
rect 85900 80 85940 2323
rect 86091 1532 86133 1541
rect 86091 1492 86092 1532
rect 86132 1492 86133 1532
rect 86091 1483 86133 1492
rect 86092 80 86132 1483
rect 86188 1373 86228 2500
rect 86284 2500 86420 2540
rect 86476 3212 86516 3221
rect 86572 3212 86612 3928
rect 86668 3464 86708 3473
rect 86764 3464 86804 4255
rect 86860 3968 86900 3977
rect 86860 3809 86900 3928
rect 86859 3800 86901 3809
rect 86859 3760 86860 3800
rect 86900 3760 86901 3800
rect 86859 3751 86901 3760
rect 86859 3548 86901 3557
rect 86859 3508 86860 3548
rect 86900 3508 86901 3548
rect 86859 3499 86901 3508
rect 86708 3424 86804 3464
rect 86668 3415 86708 3424
rect 86860 3389 86900 3499
rect 86859 3380 86901 3389
rect 86859 3340 86860 3380
rect 86900 3340 86901 3380
rect 86859 3331 86901 3340
rect 86860 3212 86900 3221
rect 86572 3172 86804 3212
rect 86187 1364 86229 1373
rect 86187 1324 86188 1364
rect 86228 1324 86229 1364
rect 86187 1315 86229 1324
rect 86284 80 86324 2500
rect 86476 1457 86516 3172
rect 86667 2960 86709 2969
rect 86667 2920 86668 2960
rect 86708 2920 86709 2960
rect 86667 2911 86709 2920
rect 86668 2633 86708 2911
rect 86667 2624 86709 2633
rect 86667 2584 86668 2624
rect 86708 2584 86709 2624
rect 86667 2575 86709 2584
rect 86571 2540 86613 2549
rect 86571 2500 86572 2540
rect 86612 2500 86613 2540
rect 86571 2491 86613 2500
rect 86475 1448 86517 1457
rect 86475 1408 86476 1448
rect 86516 1408 86517 1448
rect 86475 1399 86517 1408
rect 86572 1280 86612 2491
rect 86667 1364 86709 1373
rect 86667 1324 86668 1364
rect 86708 1324 86709 1364
rect 86667 1315 86709 1324
rect 86476 1240 86612 1280
rect 86476 80 86516 1240
rect 86668 80 86708 1315
rect 86764 785 86804 3172
rect 86860 1625 86900 3172
rect 86956 2549 86996 4684
rect 87148 4675 87188 4684
rect 87052 4136 87092 4145
rect 87244 4136 87284 7876
rect 87340 7169 87380 8464
rect 87435 8504 87477 8513
rect 87435 8464 87436 8504
rect 87476 8464 87477 8504
rect 87435 8455 87477 8464
rect 87339 7160 87381 7169
rect 87339 7120 87340 7160
rect 87380 7120 87381 7160
rect 87339 7111 87381 7120
rect 87339 6992 87381 7001
rect 87339 6952 87340 6992
rect 87380 6952 87381 6992
rect 87339 6943 87381 6952
rect 87340 4976 87380 6943
rect 87436 6581 87476 8455
rect 87531 8168 87573 8177
rect 87531 8128 87532 8168
rect 87572 8128 87573 8168
rect 87531 8119 87573 8128
rect 87532 8000 87572 8119
rect 87532 7951 87572 7960
rect 87627 7832 87669 7841
rect 87627 7792 87628 7832
rect 87668 7792 87669 7832
rect 87627 7783 87669 7792
rect 87531 7244 87573 7253
rect 87531 7204 87532 7244
rect 87572 7204 87573 7244
rect 87531 7195 87573 7204
rect 87532 7110 87572 7195
rect 87628 7169 87668 7783
rect 87724 7748 87764 8632
rect 87819 8336 87861 8345
rect 87819 8296 87820 8336
rect 87860 8296 87861 8336
rect 87819 8287 87861 8296
rect 87820 7916 87860 8287
rect 87916 8000 87956 8791
rect 88011 8756 88053 8765
rect 88011 8716 88012 8756
rect 88052 8716 88053 8756
rect 88011 8707 88053 8716
rect 88012 8622 88052 8707
rect 88108 8672 88148 9715
rect 88203 9512 88245 9521
rect 88203 9472 88204 9512
rect 88244 9472 88245 9512
rect 88203 9463 88245 9472
rect 88204 9428 88244 9463
rect 88204 9377 88244 9388
rect 88396 9428 88436 9437
rect 88492 9428 88532 10228
rect 88588 9605 88628 10228
rect 88683 10268 88725 10277
rect 88683 10228 88684 10268
rect 88724 10228 88725 10268
rect 88683 10219 88725 10228
rect 88780 10268 88820 10277
rect 89164 10268 89204 10303
rect 88820 10228 88821 10268
rect 88780 10219 88821 10228
rect 88684 10134 88724 10219
rect 88781 10184 88821 10219
rect 88963 10253 89003 10262
rect 88963 10193 89003 10213
rect 88963 10184 89013 10193
rect 88781 10144 88972 10184
rect 89012 10144 89013 10184
rect 88587 9596 88629 9605
rect 88587 9556 88588 9596
rect 88628 9556 88629 9596
rect 88587 9547 88629 9556
rect 88588 9428 88628 9437
rect 88492 9388 88588 9428
rect 88300 9344 88340 9353
rect 88203 9260 88245 9269
rect 88203 9220 88204 9260
rect 88244 9220 88245 9260
rect 88203 9211 88245 9220
rect 88204 8769 88244 9211
rect 88204 8720 88244 8729
rect 88108 8632 88244 8672
rect 88107 8504 88149 8513
rect 88107 8464 88108 8504
rect 88148 8464 88149 8504
rect 88107 8455 88149 8464
rect 88108 8370 88148 8455
rect 88204 8345 88244 8632
rect 88203 8336 88245 8345
rect 88203 8296 88204 8336
rect 88244 8296 88245 8336
rect 88203 8287 88245 8296
rect 88203 8168 88245 8177
rect 88203 8128 88204 8168
rect 88244 8128 88245 8168
rect 88203 8119 88245 8128
rect 87916 7960 88052 8000
rect 87820 7867 87860 7876
rect 88012 7916 88052 7960
rect 87916 7832 87956 7841
rect 87819 7748 87861 7757
rect 87724 7708 87820 7748
rect 87860 7708 87861 7748
rect 87819 7699 87861 7708
rect 87723 7328 87765 7337
rect 87723 7288 87724 7328
rect 87764 7288 87765 7328
rect 87723 7279 87765 7288
rect 87724 7244 87764 7279
rect 87724 7193 87764 7204
rect 87627 7160 87669 7169
rect 87627 7120 87628 7160
rect 87668 7120 87669 7160
rect 87627 7111 87669 7120
rect 87724 6656 87764 6665
rect 87820 6656 87860 7699
rect 87764 6616 87860 6656
rect 87724 6607 87764 6616
rect 87435 6572 87477 6581
rect 87435 6532 87436 6572
rect 87476 6532 87477 6572
rect 87435 6523 87477 6532
rect 87436 6404 87476 6415
rect 87916 6404 87956 7792
rect 88012 7412 88052 7876
rect 88204 7916 88244 8119
rect 88300 8084 88340 9304
rect 88396 9269 88436 9388
rect 88588 9379 88628 9388
rect 88780 9428 88820 9437
rect 88684 9344 88724 9353
rect 88395 9260 88437 9269
rect 88395 9220 88396 9260
rect 88436 9220 88437 9260
rect 88395 9211 88437 9220
rect 88396 8765 88436 9211
rect 88395 8756 88437 8765
rect 88395 8716 88396 8756
rect 88436 8716 88437 8756
rect 88395 8707 88437 8716
rect 88684 8177 88724 9304
rect 88780 9269 88820 9388
rect 88779 9260 88821 9269
rect 88779 9220 88780 9260
rect 88820 9220 88821 9260
rect 88779 9211 88821 9220
rect 88876 8849 88916 10144
rect 88963 10135 89013 10144
rect 88963 10029 89003 10135
rect 89067 10100 89109 10109
rect 89067 10060 89068 10100
rect 89108 10060 89109 10100
rect 89067 10051 89109 10060
rect 89068 9966 89108 10051
rect 88972 9428 89012 9437
rect 88972 9185 89012 9388
rect 89164 9428 89204 10228
rect 89452 10268 89492 10279
rect 89452 10193 89492 10228
rect 89644 10268 89684 10387
rect 89644 10219 89684 10228
rect 89451 10184 89493 10193
rect 89451 10144 89452 10184
rect 89492 10144 89493 10184
rect 89451 10135 89493 10144
rect 89548 10016 89588 10025
rect 89588 9976 89684 10016
rect 89548 9967 89588 9976
rect 89356 9428 89396 9437
rect 89204 9388 89356 9428
rect 89164 9379 89204 9388
rect 89356 9379 89396 9388
rect 89548 9428 89588 9437
rect 89067 9344 89109 9353
rect 89067 9304 89068 9344
rect 89108 9304 89109 9344
rect 89067 9295 89109 9304
rect 89452 9344 89492 9353
rect 89068 9210 89108 9295
rect 89452 9260 89492 9304
rect 89548 9269 89588 9388
rect 89260 9220 89492 9260
rect 89547 9260 89589 9269
rect 89547 9220 89548 9260
rect 89588 9220 89589 9260
rect 88971 9176 89013 9185
rect 88971 9136 88972 9176
rect 89012 9136 89013 9176
rect 88971 9127 89013 9136
rect 88875 8840 88917 8849
rect 88875 8800 88876 8840
rect 88916 8800 88917 8840
rect 88875 8791 88917 8800
rect 88972 8756 89012 9127
rect 89067 8840 89109 8849
rect 89067 8800 89068 8840
rect 89108 8800 89109 8840
rect 89067 8791 89109 8800
rect 88683 8168 88725 8177
rect 88683 8128 88684 8168
rect 88724 8128 88725 8168
rect 88683 8119 88725 8128
rect 88300 8044 88532 8084
rect 88204 7867 88244 7876
rect 88395 7916 88437 7925
rect 88395 7876 88396 7916
rect 88436 7876 88437 7916
rect 88395 7867 88437 7876
rect 88299 7832 88341 7841
rect 88299 7792 88300 7832
rect 88340 7792 88341 7832
rect 88299 7783 88341 7792
rect 88300 7698 88340 7783
rect 88396 7782 88436 7867
rect 88203 7496 88245 7505
rect 88180 7456 88204 7496
rect 88244 7456 88245 7496
rect 88180 7447 88245 7456
rect 88180 7412 88220 7447
rect 88012 7372 88220 7412
rect 88012 7244 88052 7253
rect 88012 7085 88052 7204
rect 88204 7244 88244 7253
rect 88204 7085 88244 7204
rect 88011 7076 88053 7085
rect 88011 7036 88012 7076
rect 88052 7036 88053 7076
rect 88011 7027 88053 7036
rect 88203 7076 88245 7085
rect 88203 7036 88204 7076
rect 88244 7036 88245 7076
rect 88203 7027 88245 7036
rect 88107 6992 88149 7001
rect 88107 6952 88108 6992
rect 88148 6952 88149 6992
rect 88107 6943 88149 6952
rect 88108 6858 88148 6943
rect 87436 6329 87476 6364
rect 87628 6364 87956 6404
rect 87435 6320 87477 6329
rect 87435 6280 87436 6320
rect 87476 6280 87477 6320
rect 87435 6271 87477 6280
rect 87340 4927 87380 4936
rect 87532 4724 87572 4733
rect 87052 3641 87092 4096
rect 87148 4096 87284 4136
rect 87340 4684 87532 4724
rect 87051 3632 87093 3641
rect 87051 3592 87052 3632
rect 87092 3592 87093 3632
rect 87051 3583 87093 3592
rect 87148 3557 87188 4096
rect 87243 3968 87285 3977
rect 87243 3928 87244 3968
rect 87284 3928 87285 3968
rect 87243 3919 87285 3928
rect 87244 3834 87284 3919
rect 87147 3548 87189 3557
rect 87147 3508 87148 3548
rect 87188 3508 87189 3548
rect 87147 3499 87189 3508
rect 87052 3464 87092 3473
rect 87052 3221 87092 3424
rect 87340 3380 87380 4684
rect 87532 4675 87572 4684
rect 87435 4472 87477 4481
rect 87435 4432 87436 4472
rect 87476 4432 87477 4472
rect 87435 4423 87477 4432
rect 87436 4136 87476 4423
rect 87628 4136 87668 6364
rect 87819 6236 87861 6245
rect 87819 6196 87820 6236
rect 87860 6196 87861 6236
rect 87819 6187 87861 6196
rect 87723 4976 87765 4985
rect 87723 4936 87724 4976
rect 87764 4936 87765 4976
rect 87723 4927 87765 4936
rect 87724 4842 87764 4927
rect 87436 4087 87476 4096
rect 87532 4096 87668 4136
rect 87820 4136 87860 6187
rect 88492 5144 88532 8044
rect 88587 7916 88629 7925
rect 88587 7876 88588 7916
rect 88628 7876 88629 7916
rect 88587 7867 88629 7876
rect 88684 7916 88724 7925
rect 88972 7916 89012 8716
rect 89068 8706 89108 8791
rect 89164 8756 89204 8767
rect 89164 8681 89204 8716
rect 89163 8672 89205 8681
rect 89163 8632 89164 8672
rect 89204 8632 89205 8672
rect 89163 8623 89205 8632
rect 89260 8177 89300 9220
rect 89547 9211 89589 9220
rect 89355 8756 89397 8765
rect 89355 8716 89356 8756
rect 89396 8716 89397 8756
rect 89355 8707 89397 8716
rect 89548 8756 89588 8767
rect 89356 8622 89396 8707
rect 89548 8681 89588 8716
rect 89547 8672 89589 8681
rect 89547 8632 89548 8672
rect 89588 8632 89589 8672
rect 89547 8623 89589 8632
rect 89644 8588 89684 9976
rect 89740 9428 89780 9437
rect 89740 9269 89780 9388
rect 89932 9428 89972 10387
rect 92427 10268 92469 10277
rect 92427 10228 92428 10268
rect 92468 10228 92469 10268
rect 92427 10219 92469 10228
rect 90027 9680 90069 9689
rect 90027 9640 90028 9680
rect 90068 9640 90069 9680
rect 90027 9631 90069 9640
rect 89932 9379 89972 9388
rect 89836 9344 89876 9353
rect 89739 9260 89781 9269
rect 89739 9220 89740 9260
rect 89780 9220 89781 9260
rect 89739 9211 89781 9220
rect 89836 9185 89876 9304
rect 89835 9176 89877 9185
rect 89835 9136 89836 9176
rect 89876 9136 89877 9176
rect 89835 9127 89877 9136
rect 89644 8548 89876 8588
rect 89452 8504 89492 8513
rect 89492 8464 89780 8504
rect 89452 8455 89492 8464
rect 89451 8336 89493 8345
rect 89451 8296 89452 8336
rect 89492 8296 89493 8336
rect 89451 8287 89493 8296
rect 89259 8168 89301 8177
rect 89259 8128 89260 8168
rect 89300 8128 89301 8168
rect 89259 8119 89301 8128
rect 89452 8000 89492 8287
rect 89263 7960 89684 8000
rect 89263 7939 89303 7960
rect 89068 7916 89108 7925
rect 88588 7782 88628 7867
rect 88587 7580 88629 7589
rect 88587 7540 88588 7580
rect 88628 7540 88629 7580
rect 88587 7531 88629 7540
rect 88588 6908 88628 7531
rect 88684 7085 88724 7876
rect 88789 7903 88829 7912
rect 88972 7876 89068 7916
rect 89644 7916 89684 7960
rect 89263 7890 89303 7899
rect 89452 7903 89492 7912
rect 89068 7867 89108 7876
rect 88789 7832 88829 7863
rect 89644 7867 89684 7876
rect 89164 7832 89204 7841
rect 88789 7792 89012 7832
rect 88972 7673 89012 7792
rect 89164 7673 89204 7792
rect 89452 7757 89492 7863
rect 89548 7832 89588 7841
rect 89451 7748 89493 7757
rect 89451 7708 89452 7748
rect 89492 7708 89493 7748
rect 89451 7699 89493 7708
rect 88971 7664 89013 7673
rect 88971 7624 88972 7664
rect 89012 7624 89013 7664
rect 88971 7615 89013 7624
rect 89163 7664 89205 7673
rect 89163 7624 89164 7664
rect 89204 7624 89205 7664
rect 89163 7615 89205 7624
rect 88779 7496 88821 7505
rect 88779 7456 88780 7496
rect 88820 7456 88821 7496
rect 88779 7447 88821 7456
rect 88683 7076 88725 7085
rect 88683 7036 88684 7076
rect 88724 7036 88725 7076
rect 88683 7027 88725 7036
rect 88588 6868 88724 6908
rect 88587 6740 88629 6749
rect 88587 6700 88588 6740
rect 88628 6700 88629 6740
rect 88587 6691 88629 6700
rect 88396 5104 88532 5144
rect 88107 4976 88149 4985
rect 88107 4936 88108 4976
rect 88148 4936 88149 4976
rect 88107 4927 88149 4936
rect 88108 4842 88148 4927
rect 88203 4892 88245 4901
rect 88203 4852 88204 4892
rect 88244 4852 88245 4892
rect 88203 4843 88245 4852
rect 87916 4724 87956 4733
rect 87956 4684 88148 4724
rect 87916 4675 87956 4684
rect 87436 3464 87476 3473
rect 87532 3464 87572 4096
rect 87820 4087 87860 4096
rect 87628 3968 87668 3977
rect 88012 3968 88052 3977
rect 87668 3928 87764 3968
rect 87628 3919 87668 3928
rect 87476 3424 87572 3464
rect 87436 3415 87476 3424
rect 87148 3340 87380 3380
rect 87051 3212 87093 3221
rect 87051 3172 87052 3212
rect 87092 3172 87093 3212
rect 87051 3163 87093 3172
rect 86955 2540 86997 2549
rect 87148 2540 87188 3340
rect 86955 2500 86956 2540
rect 86996 2500 86997 2540
rect 86955 2491 86997 2500
rect 87052 2500 87188 2540
rect 87244 3212 87284 3221
rect 87244 2540 87284 3172
rect 87435 3212 87477 3221
rect 87628 3212 87668 3221
rect 87435 3172 87436 3212
rect 87476 3172 87477 3212
rect 87435 3163 87477 3172
rect 87532 3172 87628 3212
rect 87244 2500 87380 2540
rect 86859 1616 86901 1625
rect 86859 1576 86860 1616
rect 86900 1576 86901 1616
rect 86859 1567 86901 1576
rect 86859 1112 86901 1121
rect 86859 1072 86860 1112
rect 86900 1072 86901 1112
rect 86859 1063 86901 1072
rect 86763 776 86805 785
rect 86763 736 86764 776
rect 86804 736 86805 776
rect 86763 727 86805 736
rect 86860 80 86900 1063
rect 87052 80 87092 2500
rect 87243 1448 87285 1457
rect 87243 1408 87244 1448
rect 87284 1408 87285 1448
rect 87243 1399 87285 1408
rect 87244 80 87284 1399
rect 87340 533 87380 2500
rect 87339 524 87381 533
rect 87339 484 87340 524
rect 87380 484 87381 524
rect 87339 475 87381 484
rect 87436 80 87476 3163
rect 87532 701 87572 3172
rect 87628 3163 87668 3172
rect 87724 3044 87764 3928
rect 87916 3928 88012 3968
rect 87819 3548 87861 3557
rect 87819 3508 87820 3548
rect 87860 3508 87861 3548
rect 87819 3499 87861 3508
rect 87820 3464 87860 3499
rect 87820 3413 87860 3424
rect 87628 3004 87764 3044
rect 87628 2549 87668 3004
rect 87723 2708 87765 2717
rect 87723 2668 87724 2708
rect 87764 2668 87765 2708
rect 87723 2659 87765 2668
rect 87627 2540 87669 2549
rect 87627 2500 87628 2540
rect 87668 2500 87669 2540
rect 87627 2491 87669 2500
rect 87724 1280 87764 2659
rect 87916 1373 87956 3928
rect 88012 3919 88052 3928
rect 88012 3212 88052 3221
rect 88012 2540 88052 3172
rect 88108 2717 88148 4684
rect 88204 4136 88244 4843
rect 88204 4087 88244 4096
rect 88300 4724 88340 4733
rect 88203 3968 88245 3977
rect 88203 3928 88204 3968
rect 88244 3928 88245 3968
rect 88203 3919 88245 3928
rect 88204 3464 88244 3919
rect 88204 3415 88244 3424
rect 88107 2708 88149 2717
rect 88107 2668 88108 2708
rect 88148 2668 88149 2708
rect 88107 2659 88149 2668
rect 88300 2540 88340 4684
rect 88396 4145 88436 5104
rect 88491 4976 88533 4985
rect 88491 4936 88492 4976
rect 88532 4936 88533 4976
rect 88491 4927 88533 4936
rect 88492 4842 88532 4927
rect 88395 4136 88437 4145
rect 88395 4096 88396 4136
rect 88436 4096 88437 4136
rect 88395 4087 88437 4096
rect 88588 4136 88628 6691
rect 88684 4901 88724 6868
rect 88780 5069 88820 7447
rect 88972 7412 89012 7615
rect 89355 7580 89397 7589
rect 89355 7540 89356 7580
rect 89396 7540 89397 7580
rect 89355 7531 89397 7540
rect 89068 7412 89108 7421
rect 88972 7372 89068 7412
rect 89068 7363 89108 7372
rect 89067 5144 89109 5153
rect 89067 5104 89068 5144
rect 89108 5104 89109 5144
rect 89067 5095 89109 5104
rect 88779 5060 88821 5069
rect 88779 5020 88780 5060
rect 88820 5020 88821 5060
rect 88779 5011 88821 5020
rect 88683 4892 88725 4901
rect 88683 4852 88684 4892
rect 88724 4852 88725 4892
rect 88683 4843 88725 4852
rect 88971 4724 89013 4733
rect 88971 4684 88972 4724
rect 89012 4684 89013 4724
rect 88971 4675 89013 4684
rect 88972 4149 89012 4675
rect 88972 4100 89012 4109
rect 88588 4087 88628 4096
rect 89068 4052 89108 5095
rect 89356 4136 89396 7531
rect 89452 7244 89492 7699
rect 89452 7195 89492 7204
rect 89548 6329 89588 7792
rect 89643 6908 89685 6917
rect 89643 6868 89644 6908
rect 89684 6868 89685 6908
rect 89643 6859 89685 6868
rect 89547 6320 89589 6329
rect 89547 6280 89548 6320
rect 89588 6280 89589 6320
rect 89547 6271 89589 6280
rect 89644 4817 89684 6859
rect 89740 5069 89780 8464
rect 89739 5060 89781 5069
rect 89739 5020 89740 5060
rect 89780 5020 89781 5060
rect 89739 5011 89781 5020
rect 89643 4808 89685 4817
rect 89643 4768 89644 4808
rect 89684 4768 89685 4808
rect 89643 4759 89685 4768
rect 89739 4304 89781 4313
rect 89739 4264 89740 4304
rect 89780 4264 89781 4304
rect 89739 4255 89781 4264
rect 89356 4087 89396 4096
rect 89740 4136 89780 4255
rect 89836 4145 89876 8548
rect 89931 8252 89973 8261
rect 89931 8212 89932 8252
rect 89972 8212 89973 8252
rect 89931 8203 89973 8212
rect 89932 4313 89972 8203
rect 89931 4304 89973 4313
rect 89931 4264 89932 4304
rect 89972 4264 89973 4304
rect 89931 4255 89973 4264
rect 89740 4087 89780 4096
rect 89835 4136 89877 4145
rect 89835 4096 89836 4136
rect 89876 4096 89877 4136
rect 89835 4087 89877 4096
rect 88972 4012 89108 4052
rect 88396 3968 88436 3977
rect 88780 3968 88820 3977
rect 88436 3928 88532 3968
rect 88396 3919 88436 3928
rect 88012 2500 88148 2540
rect 88011 1616 88053 1625
rect 88011 1576 88012 1616
rect 88052 1576 88053 1616
rect 88011 1567 88053 1576
rect 87915 1364 87957 1373
rect 87915 1324 87916 1364
rect 87956 1324 87957 1364
rect 87915 1315 87957 1324
rect 87628 1240 87764 1280
rect 87819 1280 87861 1289
rect 87819 1240 87820 1280
rect 87860 1240 87861 1280
rect 87531 692 87573 701
rect 87531 652 87532 692
rect 87572 652 87573 692
rect 87531 643 87573 652
rect 87628 80 87668 1240
rect 87819 1231 87861 1240
rect 87820 80 87860 1231
rect 88012 80 88052 1567
rect 88108 1037 88148 2500
rect 88204 2500 88340 2540
rect 88396 3212 88436 3221
rect 88107 1028 88149 1037
rect 88107 988 88108 1028
rect 88148 988 88149 1028
rect 88107 979 88149 988
rect 88204 80 88244 2500
rect 88396 1541 88436 3172
rect 88395 1532 88437 1541
rect 88395 1492 88396 1532
rect 88436 1492 88437 1532
rect 88395 1483 88437 1492
rect 88492 1457 88532 3928
rect 88684 3928 88780 3968
rect 88587 3464 88629 3473
rect 88587 3424 88588 3464
rect 88628 3424 88629 3464
rect 88587 3415 88629 3424
rect 88588 3330 88628 3415
rect 88587 3044 88629 3053
rect 88587 3004 88588 3044
rect 88628 3004 88629 3044
rect 88587 2995 88629 3004
rect 88588 2717 88628 2995
rect 88587 2708 88629 2717
rect 88587 2668 88588 2708
rect 88628 2668 88629 2708
rect 88587 2659 88629 2668
rect 88587 1952 88629 1961
rect 88587 1912 88588 1952
rect 88628 1912 88629 1952
rect 88587 1903 88629 1912
rect 88491 1448 88533 1457
rect 88491 1408 88492 1448
rect 88532 1408 88533 1448
rect 88491 1399 88533 1408
rect 88395 1364 88437 1373
rect 88395 1324 88396 1364
rect 88436 1324 88437 1364
rect 88395 1315 88437 1324
rect 88396 80 88436 1315
rect 88588 80 88628 1903
rect 88684 1289 88724 3928
rect 88780 3919 88820 3928
rect 88972 3464 89012 4012
rect 89164 3968 89204 3977
rect 89548 3968 89588 3977
rect 89932 3968 89972 3977
rect 88972 3415 89012 3424
rect 89068 3928 89164 3968
rect 88780 3212 88820 3221
rect 88683 1280 88725 1289
rect 88683 1240 88684 1280
rect 88724 1240 88725 1280
rect 88683 1231 88725 1240
rect 88780 1121 88820 3172
rect 88875 2456 88917 2465
rect 88875 2416 88876 2456
rect 88916 2416 88917 2456
rect 88875 2407 88917 2416
rect 88876 1709 88916 2407
rect 88875 1700 88917 1709
rect 88875 1660 88876 1700
rect 88916 1660 88917 1700
rect 88875 1651 88917 1660
rect 88971 1532 89013 1541
rect 88971 1492 88972 1532
rect 89012 1492 89013 1532
rect 88971 1483 89013 1492
rect 88779 1112 88821 1121
rect 88779 1072 88780 1112
rect 88820 1072 88821 1112
rect 88779 1063 88821 1072
rect 88779 104 88821 113
rect 88779 80 88780 104
rect 38132 64 38152 80
rect 38072 0 38152 64
rect 38264 0 38344 80
rect 38456 0 38536 80
rect 38648 0 38728 80
rect 38840 0 38920 80
rect 39032 0 39112 80
rect 39224 0 39304 80
rect 39416 0 39496 80
rect 39608 0 39688 80
rect 39800 0 39880 80
rect 39992 0 40072 80
rect 40184 0 40264 80
rect 40376 0 40456 80
rect 40568 0 40648 80
rect 40760 0 40840 80
rect 40952 0 41032 80
rect 41144 0 41224 80
rect 41336 0 41416 80
rect 41528 0 41608 80
rect 41720 0 41800 80
rect 41912 0 41992 80
rect 42104 0 42184 80
rect 42231 64 42376 80
rect 42296 0 42376 64
rect 42488 0 42568 80
rect 42680 0 42760 80
rect 42872 0 42952 80
rect 43064 0 43144 80
rect 43256 0 43336 80
rect 43448 0 43528 80
rect 43640 0 43720 80
rect 43832 0 43912 80
rect 44024 0 44104 80
rect 44216 0 44296 80
rect 44408 0 44488 80
rect 44600 0 44680 80
rect 44792 0 44872 80
rect 44984 0 45064 80
rect 45176 0 45256 80
rect 45368 0 45448 80
rect 45560 0 45640 80
rect 45752 0 45832 80
rect 45944 0 46024 80
rect 46136 0 46216 80
rect 46328 0 46408 80
rect 46520 0 46600 80
rect 46712 0 46792 80
rect 46904 0 46984 80
rect 47096 0 47176 80
rect 47288 0 47368 80
rect 47480 0 47560 80
rect 47672 0 47752 80
rect 47864 0 47944 80
rect 48056 0 48136 80
rect 48248 0 48328 80
rect 48440 0 48520 80
rect 48632 0 48712 80
rect 48824 0 48904 80
rect 49016 0 49096 80
rect 49208 0 49288 80
rect 49400 0 49480 80
rect 49592 0 49672 80
rect 49784 0 49864 80
rect 49976 0 50056 80
rect 50168 0 50248 80
rect 50360 0 50440 80
rect 50552 0 50632 80
rect 50744 0 50824 80
rect 50936 0 51016 80
rect 51128 0 51208 80
rect 51320 0 51400 80
rect 51512 0 51592 80
rect 51704 0 51784 80
rect 51896 0 51976 80
rect 52088 0 52168 80
rect 52280 0 52360 80
rect 52472 0 52552 80
rect 52664 0 52744 80
rect 52856 0 52936 80
rect 53048 0 53128 80
rect 53240 0 53320 80
rect 53432 0 53512 80
rect 53624 0 53704 80
rect 53816 0 53896 80
rect 54008 0 54088 80
rect 54200 0 54280 80
rect 54392 0 54472 80
rect 54584 0 54664 80
rect 54776 0 54856 80
rect 54968 0 55048 80
rect 55160 0 55240 80
rect 55352 0 55432 80
rect 55544 0 55624 80
rect 55736 0 55816 80
rect 55928 0 56008 80
rect 56120 0 56200 80
rect 56312 0 56392 80
rect 56504 0 56584 80
rect 56696 0 56776 80
rect 56888 0 56968 80
rect 57080 0 57160 80
rect 57272 0 57352 80
rect 57464 0 57544 80
rect 57656 0 57736 80
rect 57848 0 57928 80
rect 58040 0 58120 80
rect 58232 0 58312 80
rect 58424 0 58504 80
rect 58616 0 58696 80
rect 58808 0 58888 80
rect 59000 0 59080 80
rect 59192 0 59272 80
rect 59384 0 59464 80
rect 59576 0 59656 80
rect 59768 0 59848 80
rect 59960 0 60040 80
rect 60152 0 60232 80
rect 60344 0 60424 80
rect 60536 0 60616 80
rect 60728 0 60808 80
rect 60920 0 61000 80
rect 61112 0 61192 80
rect 61304 0 61384 80
rect 61496 0 61576 80
rect 61688 0 61768 80
rect 61880 0 61960 80
rect 62072 0 62152 80
rect 62264 0 62344 80
rect 62456 0 62536 80
rect 62648 0 62728 80
rect 62840 0 62920 80
rect 63032 0 63112 80
rect 63224 0 63304 80
rect 63416 0 63496 80
rect 63608 0 63688 80
rect 63800 0 63880 80
rect 63992 0 64072 80
rect 64184 0 64264 80
rect 64376 0 64456 80
rect 64568 0 64648 80
rect 64760 0 64840 80
rect 64952 0 65032 80
rect 65144 0 65224 80
rect 65336 0 65416 80
rect 65528 0 65608 80
rect 65720 0 65800 80
rect 65912 0 65992 80
rect 66104 0 66184 80
rect 66296 0 66376 80
rect 66488 0 66568 80
rect 66680 0 66760 80
rect 66872 0 66952 80
rect 67064 0 67144 80
rect 67256 0 67336 80
rect 67448 0 67528 80
rect 67640 0 67720 80
rect 67832 0 67912 80
rect 68024 0 68104 80
rect 68216 0 68296 80
rect 68408 0 68488 80
rect 68600 0 68680 80
rect 68792 0 68872 80
rect 68984 0 69064 80
rect 69176 0 69256 80
rect 69368 0 69448 80
rect 69560 0 69640 80
rect 69752 0 69832 80
rect 69944 0 70024 80
rect 70136 0 70216 80
rect 70328 0 70408 80
rect 70520 0 70600 80
rect 70712 0 70792 80
rect 70904 0 70984 80
rect 71096 0 71176 80
rect 71288 0 71368 80
rect 71480 0 71560 80
rect 71672 0 71752 80
rect 71864 0 71944 80
rect 72056 0 72136 80
rect 72248 0 72328 80
rect 72440 0 72520 80
rect 72632 0 72712 80
rect 72824 0 72904 80
rect 73016 0 73096 80
rect 73208 0 73288 80
rect 73400 0 73480 80
rect 73592 0 73672 80
rect 73784 0 73864 80
rect 73976 0 74056 80
rect 74168 0 74248 80
rect 74360 0 74440 80
rect 74552 0 74632 80
rect 74744 0 74824 80
rect 74936 0 75016 80
rect 75128 0 75208 80
rect 75320 0 75400 80
rect 75512 0 75592 80
rect 75704 0 75784 80
rect 75896 0 75976 80
rect 76088 0 76168 80
rect 76280 0 76360 80
rect 76472 0 76552 80
rect 76664 0 76744 80
rect 76856 0 76936 80
rect 77048 0 77128 80
rect 77240 0 77320 80
rect 77432 0 77512 80
rect 77624 0 77704 80
rect 77816 0 77896 80
rect 78008 0 78088 80
rect 78200 0 78280 80
rect 78392 0 78472 80
rect 78584 0 78664 80
rect 78776 0 78856 80
rect 78968 0 79048 80
rect 79160 0 79240 80
rect 79352 0 79432 80
rect 79544 0 79624 80
rect 79736 0 79816 80
rect 79928 0 80008 80
rect 80120 0 80200 80
rect 80312 0 80392 80
rect 80504 0 80584 80
rect 80696 0 80776 80
rect 80888 0 80968 80
rect 81080 0 81160 80
rect 81272 0 81352 80
rect 81464 0 81544 80
rect 81656 0 81736 80
rect 81848 0 81928 80
rect 82040 0 82120 80
rect 82232 0 82312 80
rect 82424 0 82504 80
rect 82616 0 82696 80
rect 82808 0 82888 80
rect 83000 0 83080 80
rect 83192 0 83272 80
rect 83384 0 83464 80
rect 83576 0 83656 80
rect 83768 0 83848 80
rect 83960 0 84040 80
rect 84152 0 84232 80
rect 84344 0 84424 80
rect 84536 0 84616 80
rect 84728 0 84808 80
rect 84920 0 85000 80
rect 85112 0 85192 80
rect 85304 0 85384 80
rect 85496 0 85576 80
rect 85688 0 85768 80
rect 85880 0 85960 80
rect 86072 0 86152 80
rect 86264 0 86344 80
rect 86456 0 86536 80
rect 86648 0 86728 80
rect 86840 0 86920 80
rect 87032 0 87112 80
rect 87224 0 87304 80
rect 87416 0 87496 80
rect 87608 0 87688 80
rect 87800 0 87880 80
rect 87992 0 88072 80
rect 88184 0 88264 80
rect 88376 0 88456 80
rect 88568 0 88648 80
rect 88760 64 88780 80
rect 88820 80 88821 104
rect 88972 80 89012 1483
rect 89068 1373 89108 3928
rect 89164 3919 89204 3928
rect 89452 3928 89548 3968
rect 89452 3632 89492 3928
rect 89548 3919 89588 3928
rect 89644 3928 89932 3968
rect 89260 3592 89492 3632
rect 89163 3212 89205 3221
rect 89163 3172 89164 3212
rect 89204 3172 89205 3212
rect 89163 3163 89205 3172
rect 89164 3078 89204 3163
rect 89067 1364 89109 1373
rect 89067 1324 89068 1364
rect 89108 1324 89109 1364
rect 89067 1315 89109 1324
rect 89163 1280 89205 1289
rect 89163 1240 89164 1280
rect 89204 1240 89205 1280
rect 89163 1231 89205 1240
rect 89164 80 89204 1231
rect 89260 197 89300 3592
rect 89356 3464 89396 3473
rect 89356 2549 89396 3424
rect 89548 3212 89588 3221
rect 89355 2540 89397 2549
rect 89355 2500 89356 2540
rect 89396 2500 89397 2540
rect 89355 2491 89397 2500
rect 89355 2372 89397 2381
rect 89355 2332 89356 2372
rect 89396 2332 89397 2372
rect 89355 2323 89397 2332
rect 89259 188 89301 197
rect 89259 148 89260 188
rect 89300 148 89301 188
rect 89259 139 89301 148
rect 89356 80 89396 2323
rect 89548 1625 89588 3172
rect 89547 1616 89589 1625
rect 89547 1576 89548 1616
rect 89588 1576 89589 1616
rect 89547 1567 89589 1576
rect 89644 1289 89684 3928
rect 89932 3919 89972 3928
rect 89740 3464 89780 3473
rect 90028 3464 90068 9631
rect 92043 9008 92085 9017
rect 92043 8968 92044 9008
rect 92084 8968 92085 9008
rect 92043 8959 92085 8968
rect 90123 8420 90165 8429
rect 90123 8380 90124 8420
rect 90164 8380 90165 8420
rect 90123 8371 90165 8380
rect 90124 4136 90164 8371
rect 91947 7412 91989 7421
rect 91947 7372 91948 7412
rect 91988 7372 91989 7412
rect 91947 7363 91989 7372
rect 90507 7076 90549 7085
rect 90507 7036 90508 7076
rect 90548 7036 90549 7076
rect 90507 7027 90549 7036
rect 90124 4087 90164 4096
rect 90508 4136 90548 7027
rect 90891 6320 90933 6329
rect 90891 6280 90892 6320
rect 90932 6280 90933 6320
rect 90891 6271 90933 6280
rect 90508 4087 90548 4096
rect 90892 4136 90932 6271
rect 91275 5060 91317 5069
rect 91275 5020 91276 5060
rect 91316 5020 91317 5060
rect 91275 5011 91317 5020
rect 90892 4087 90932 4096
rect 91276 4136 91316 5011
rect 91948 4985 91988 7363
rect 91947 4976 91989 4985
rect 91947 4936 91948 4976
rect 91988 4936 91989 4976
rect 91947 4927 91989 4936
rect 91276 4087 91316 4096
rect 91659 4136 91701 4145
rect 91659 4096 91660 4136
rect 91700 4096 91701 4136
rect 91659 4087 91701 4096
rect 92044 4136 92084 8959
rect 92331 5228 92373 5237
rect 92331 5188 92332 5228
rect 92372 5188 92373 5228
rect 92331 5179 92373 5188
rect 92044 4087 92084 4096
rect 91660 4002 91700 4087
rect 90316 3968 90356 3977
rect 90700 3968 90740 3977
rect 90220 3928 90316 3968
rect 89780 3424 90068 3464
rect 90124 3464 90164 3473
rect 89740 3415 89780 3424
rect 89932 3212 89972 3221
rect 89932 1961 89972 3172
rect 90124 2129 90164 3424
rect 90123 2120 90165 2129
rect 90123 2080 90124 2120
rect 90164 2080 90165 2120
rect 90123 2071 90165 2080
rect 89931 1952 89973 1961
rect 89931 1912 89932 1952
rect 89972 1912 89973 1952
rect 89931 1903 89973 1912
rect 90220 1784 90260 3928
rect 90316 3919 90356 3928
rect 90604 3928 90700 3968
rect 90508 3464 90548 3473
rect 89740 1744 90260 1784
rect 90316 3212 90356 3221
rect 89643 1280 89685 1289
rect 89643 1240 89644 1280
rect 89684 1240 89685 1280
rect 89643 1231 89685 1240
rect 89740 1112 89780 1744
rect 89835 1616 89877 1625
rect 89835 1576 89836 1616
rect 89876 1576 89877 1616
rect 89835 1567 89877 1576
rect 90123 1616 90165 1625
rect 90123 1576 90124 1616
rect 90164 1576 90165 1616
rect 90123 1567 90165 1576
rect 89548 1072 89780 1112
rect 89548 80 89588 1072
rect 89836 944 89876 1567
rect 89931 1280 89973 1289
rect 89931 1240 89932 1280
rect 89972 1240 89973 1280
rect 89931 1231 89973 1240
rect 89740 904 89876 944
rect 89740 80 89780 904
rect 89932 80 89972 1231
rect 90124 80 90164 1567
rect 90316 1541 90356 3172
rect 90508 2297 90548 3424
rect 90507 2288 90549 2297
rect 90507 2248 90508 2288
rect 90548 2248 90549 2288
rect 90507 2239 90549 2248
rect 90604 1700 90644 3928
rect 90700 3900 90740 3928
rect 90795 3968 90837 3977
rect 91084 3968 91124 3977
rect 90795 3928 90796 3968
rect 90836 3928 90837 3968
rect 90795 3919 90837 3928
rect 90988 3928 91084 3968
rect 90700 3212 90740 3221
rect 90700 2381 90740 3172
rect 90699 2372 90741 2381
rect 90699 2332 90700 2372
rect 90740 2332 90741 2372
rect 90699 2323 90741 2332
rect 90412 1660 90644 1700
rect 90315 1532 90357 1541
rect 90315 1492 90316 1532
rect 90356 1492 90357 1532
rect 90315 1483 90357 1492
rect 90315 1364 90357 1373
rect 90315 1324 90316 1364
rect 90356 1324 90357 1364
rect 90315 1315 90357 1324
rect 90316 80 90356 1315
rect 90412 1289 90452 1660
rect 90507 1532 90549 1541
rect 90796 1532 90836 3919
rect 90892 3464 90932 3473
rect 90892 2633 90932 3424
rect 90891 2624 90933 2633
rect 90891 2584 90892 2624
rect 90932 2584 90933 2624
rect 90891 2575 90933 2584
rect 90891 1700 90933 1709
rect 90891 1660 90892 1700
rect 90932 1660 90933 1700
rect 90891 1651 90933 1660
rect 90507 1492 90508 1532
rect 90548 1492 90549 1532
rect 90507 1483 90549 1492
rect 90604 1492 90836 1532
rect 90411 1280 90453 1289
rect 90411 1240 90412 1280
rect 90452 1240 90453 1280
rect 90411 1231 90453 1240
rect 90508 80 90548 1483
rect 90604 440 90644 1492
rect 90604 400 90740 440
rect 90700 80 90740 400
rect 90892 80 90932 1651
rect 90988 1373 91028 3928
rect 91084 3919 91124 3928
rect 91467 3968 91509 3977
rect 91467 3928 91468 3968
rect 91508 3928 91509 3968
rect 91467 3919 91509 3928
rect 91755 3968 91797 3977
rect 91755 3928 91756 3968
rect 91796 3928 91797 3968
rect 91755 3919 91797 3928
rect 91852 3968 91892 3977
rect 91468 3834 91508 3919
rect 91179 3548 91221 3557
rect 91179 3508 91180 3548
rect 91220 3508 91221 3548
rect 91179 3499 91221 3508
rect 91084 3212 91124 3221
rect 91084 1793 91124 3172
rect 91083 1784 91125 1793
rect 91083 1744 91084 1784
rect 91124 1744 91125 1784
rect 91083 1735 91125 1744
rect 91180 1616 91220 3499
rect 91276 3464 91316 3473
rect 91276 2801 91316 3424
rect 91659 3464 91701 3473
rect 91659 3424 91660 3464
rect 91700 3424 91701 3464
rect 91659 3415 91701 3424
rect 91660 3330 91700 3415
rect 91468 3212 91508 3221
rect 91275 2792 91317 2801
rect 91275 2752 91276 2792
rect 91316 2752 91317 2792
rect 91275 2743 91317 2752
rect 91275 1784 91317 1793
rect 91275 1744 91276 1784
rect 91316 1744 91317 1784
rect 91275 1735 91317 1744
rect 91084 1576 91220 1616
rect 90987 1364 91029 1373
rect 90987 1324 90988 1364
rect 91028 1324 91029 1364
rect 90987 1315 91029 1324
rect 91084 80 91124 1576
rect 91276 80 91316 1735
rect 91468 1625 91508 3172
rect 91756 1784 91796 3919
rect 91852 3557 91892 3928
rect 92235 3968 92277 3977
rect 92235 3928 92236 3968
rect 92276 3928 92277 3968
rect 92235 3919 92277 3928
rect 92236 3834 92276 3919
rect 91947 3800 91989 3809
rect 91947 3760 91948 3800
rect 91988 3760 91989 3800
rect 91947 3751 91989 3760
rect 91851 3548 91893 3557
rect 91851 3508 91852 3548
rect 91892 3508 91893 3548
rect 91851 3499 91893 3508
rect 91564 1744 91796 1784
rect 91852 3212 91892 3221
rect 91467 1616 91509 1625
rect 91467 1576 91468 1616
rect 91508 1576 91509 1616
rect 91467 1567 91509 1576
rect 91564 1448 91604 1744
rect 91659 1616 91701 1625
rect 91659 1576 91660 1616
rect 91700 1576 91701 1616
rect 91659 1567 91701 1576
rect 91468 1408 91604 1448
rect 91468 80 91508 1408
rect 91660 80 91700 1567
rect 91852 1541 91892 3172
rect 91851 1532 91893 1541
rect 91851 1492 91852 1532
rect 91892 1492 91893 1532
rect 91851 1483 91893 1492
rect 91948 1364 91988 3751
rect 92043 3464 92085 3473
rect 92043 3424 92044 3464
rect 92084 3424 92085 3464
rect 92332 3464 92372 5179
rect 92428 4136 92468 10219
rect 92428 4087 92468 4096
rect 92812 4136 92852 10471
rect 93195 10100 93237 10109
rect 93195 10060 93196 10100
rect 93236 10060 93237 10100
rect 93195 10051 93237 10060
rect 93099 5396 93141 5405
rect 93099 5356 93100 5396
rect 93140 5356 93141 5396
rect 93099 5347 93141 5356
rect 92812 4087 92852 4096
rect 92620 3968 92660 3977
rect 93004 3968 93044 3977
rect 92620 3809 92660 3928
rect 92716 3928 93004 3968
rect 93100 3968 93140 5347
rect 93196 4136 93236 10051
rect 94408 9848 94776 9857
rect 94448 9808 94490 9848
rect 94530 9808 94572 9848
rect 94612 9808 94654 9848
rect 94694 9808 94736 9848
rect 94408 9799 94776 9808
rect 97227 9428 97269 9437
rect 97227 9388 97228 9428
rect 97268 9388 97269 9428
rect 97227 9379 97269 9388
rect 95648 9092 96016 9101
rect 95688 9052 95730 9092
rect 95770 9052 95812 9092
rect 95852 9052 95894 9092
rect 95934 9052 95976 9092
rect 95648 9043 96016 9052
rect 95787 8924 95829 8933
rect 95787 8884 95788 8924
rect 95828 8884 95829 8924
rect 95787 8875 95829 8884
rect 94408 8336 94776 8345
rect 94448 8296 94490 8336
rect 94530 8296 94572 8336
rect 94612 8296 94654 8336
rect 94694 8296 94736 8336
rect 94408 8287 94776 8296
rect 93963 8084 94005 8093
rect 93963 8044 93964 8084
rect 94004 8044 94005 8084
rect 93963 8035 94005 8044
rect 93483 5984 93525 5993
rect 93483 5944 93484 5984
rect 93524 5944 93525 5984
rect 93483 5935 93525 5944
rect 93291 4808 93333 4817
rect 93291 4768 93292 4808
rect 93332 4768 93333 4808
rect 93291 4759 93333 4768
rect 93292 4145 93332 4759
rect 93196 4087 93236 4096
rect 93291 4136 93333 4145
rect 93291 4096 93292 4136
rect 93332 4096 93333 4136
rect 93291 4087 93333 4096
rect 93388 3968 93428 3977
rect 93100 3928 93236 3968
rect 92619 3800 92661 3809
rect 92619 3760 92620 3800
rect 92660 3760 92661 3800
rect 92619 3751 92661 3760
rect 92428 3464 92468 3473
rect 92332 3424 92428 3464
rect 92043 3415 92085 3424
rect 92428 3415 92468 3424
rect 92044 3330 92084 3415
rect 92716 3380 92756 3928
rect 93004 3919 93044 3928
rect 92907 3800 92949 3809
rect 92907 3760 92908 3800
rect 92948 3760 92949 3800
rect 92907 3751 92949 3760
rect 92524 3340 92756 3380
rect 92812 3464 92852 3473
rect 92236 3212 92276 3221
rect 92236 1709 92276 3172
rect 92524 1868 92564 3340
rect 92332 1828 92564 1868
rect 92620 3212 92660 3221
rect 92235 1700 92277 1709
rect 92235 1660 92236 1700
rect 92276 1660 92277 1700
rect 92235 1651 92277 1660
rect 92043 1532 92085 1541
rect 92332 1532 92372 1828
rect 92620 1793 92660 3172
rect 92812 3137 92852 3424
rect 92811 3128 92853 3137
rect 92811 3088 92812 3128
rect 92852 3088 92853 3128
rect 92811 3079 92853 3088
rect 92908 1952 92948 3751
rect 93099 3632 93141 3641
rect 93099 3592 93100 3632
rect 93140 3592 93141 3632
rect 93099 3583 93141 3592
rect 92716 1912 92948 1952
rect 93004 3212 93044 3221
rect 92619 1784 92661 1793
rect 92619 1744 92620 1784
rect 92660 1744 92661 1784
rect 92619 1735 92661 1744
rect 92427 1700 92469 1709
rect 92427 1660 92428 1700
rect 92468 1660 92469 1700
rect 92427 1651 92469 1660
rect 92043 1492 92044 1532
rect 92084 1492 92085 1532
rect 92043 1483 92085 1492
rect 92236 1492 92372 1532
rect 91852 1324 91988 1364
rect 91852 80 91892 1324
rect 92044 80 92084 1483
rect 92236 80 92276 1492
rect 92428 80 92468 1651
rect 92716 1616 92756 1912
rect 92811 1784 92853 1793
rect 92811 1744 92812 1784
rect 92852 1744 92853 1784
rect 92811 1735 92853 1744
rect 92620 1576 92756 1616
rect 92620 80 92660 1576
rect 92812 80 92852 1735
rect 93004 1625 93044 3172
rect 93003 1616 93045 1625
rect 93003 1576 93004 1616
rect 93044 1576 93045 1616
rect 93003 1567 93045 1576
rect 93100 1448 93140 3583
rect 93196 3464 93236 3928
rect 93388 3809 93428 3928
rect 93387 3800 93429 3809
rect 93387 3760 93388 3800
rect 93428 3760 93429 3800
rect 93387 3751 93429 3760
rect 93484 3464 93524 5935
rect 93579 4556 93621 4565
rect 93579 4516 93580 4556
rect 93620 4516 93621 4556
rect 93579 4507 93621 4516
rect 93580 4136 93620 4507
rect 93580 4087 93620 4096
rect 93867 4136 93909 4145
rect 93867 4096 93868 4136
rect 93908 4096 93909 4136
rect 93867 4087 93909 4096
rect 93964 4136 94004 8035
rect 94251 8000 94293 8009
rect 94251 7960 94252 8000
rect 94292 7960 94293 8000
rect 94251 7951 94293 7960
rect 94252 5144 94292 7951
rect 95788 7757 95828 8875
rect 96651 7832 96693 7841
rect 96651 7792 96652 7832
rect 96692 7792 96693 7832
rect 96651 7783 96693 7792
rect 95787 7748 95829 7757
rect 95787 7708 95788 7748
rect 95828 7708 95829 7748
rect 95787 7699 95829 7708
rect 95648 7580 96016 7589
rect 95688 7540 95730 7580
rect 95770 7540 95812 7580
rect 95852 7540 95894 7580
rect 95934 7540 95976 7580
rect 95648 7531 96016 7540
rect 95499 7160 95541 7169
rect 95499 7120 95500 7160
rect 95540 7120 95541 7160
rect 95499 7111 95541 7120
rect 94408 6824 94776 6833
rect 94448 6784 94490 6824
rect 94530 6784 94572 6824
rect 94612 6784 94654 6824
rect 94694 6784 94736 6824
rect 94408 6775 94776 6784
rect 94408 5312 94776 5321
rect 94448 5272 94490 5312
rect 94530 5272 94572 5312
rect 94612 5272 94654 5312
rect 94694 5272 94736 5312
rect 94408 5263 94776 5272
rect 94252 5104 94388 5144
rect 93964 4087 94004 4096
rect 94348 4136 94388 5104
rect 95116 4145 95156 4230
rect 94348 4087 94388 4096
rect 94732 4136 94772 4145
rect 93772 3968 93812 3977
rect 93772 3641 93812 3928
rect 93771 3632 93813 3641
rect 93771 3592 93772 3632
rect 93812 3592 93813 3632
rect 93771 3583 93813 3592
rect 93580 3464 93620 3473
rect 93484 3424 93580 3464
rect 93868 3464 93908 4087
rect 94251 4052 94293 4061
rect 94251 4012 94252 4052
rect 94292 4012 94293 4052
rect 94251 4003 94293 4012
rect 94059 3968 94101 3977
rect 94059 3928 94060 3968
rect 94100 3928 94101 3968
rect 94059 3919 94101 3928
rect 94156 3968 94196 3977
rect 93964 3464 94004 3473
rect 93868 3424 93964 3464
rect 93196 3415 93236 3424
rect 93580 3415 93620 3424
rect 93964 3415 94004 3424
rect 93675 3380 93717 3389
rect 93675 3340 93676 3380
rect 93716 3340 93717 3380
rect 93675 3331 93717 3340
rect 93195 3212 93237 3221
rect 93195 3172 93196 3212
rect 93236 3172 93237 3212
rect 93195 3163 93237 3172
rect 93388 3212 93428 3221
rect 93004 1408 93140 1448
rect 93004 80 93044 1408
rect 93196 80 93236 3163
rect 93388 1541 93428 3172
rect 93676 1952 93716 3331
rect 93484 1912 93716 1952
rect 93772 3212 93812 3221
rect 93387 1532 93429 1541
rect 93387 1492 93388 1532
rect 93428 1492 93429 1532
rect 93387 1483 93429 1492
rect 93484 1364 93524 1912
rect 93772 1709 93812 3172
rect 94060 1868 94100 3919
rect 94156 3389 94196 3928
rect 94155 3380 94197 3389
rect 94155 3340 94156 3380
rect 94196 3340 94197 3380
rect 94155 3331 94197 3340
rect 93868 1828 94100 1868
rect 94156 3212 94196 3221
rect 93771 1700 93813 1709
rect 93771 1660 93772 1700
rect 93812 1660 93813 1700
rect 93771 1651 93813 1660
rect 93579 1616 93621 1625
rect 93579 1576 93580 1616
rect 93620 1576 93621 1616
rect 93579 1567 93621 1576
rect 93388 1324 93524 1364
rect 93388 80 93428 1324
rect 93580 80 93620 1567
rect 93868 1532 93908 1828
rect 94156 1793 94196 3172
rect 94155 1784 94197 1793
rect 94155 1744 94156 1784
rect 94196 1744 94197 1784
rect 94155 1735 94197 1744
rect 93963 1700 94005 1709
rect 93963 1660 93964 1700
rect 94004 1660 94005 1700
rect 93963 1651 94005 1660
rect 93772 1492 93908 1532
rect 93772 80 93812 1492
rect 93964 80 94004 1651
rect 94252 1616 94292 4003
rect 94540 3977 94580 4062
rect 94732 3977 94772 4096
rect 95115 4136 95157 4145
rect 95115 4096 95116 4136
rect 95156 4096 95157 4136
rect 95115 4087 95157 4096
rect 95500 4136 95540 7111
rect 95648 6068 96016 6077
rect 95688 6028 95730 6068
rect 95770 6028 95812 6068
rect 95852 6028 95894 6068
rect 95934 6028 95976 6068
rect 95648 6019 96016 6028
rect 96075 5816 96117 5825
rect 96075 5776 96076 5816
rect 96116 5776 96117 5816
rect 96075 5767 96117 5776
rect 95648 4556 96016 4565
rect 95688 4516 95730 4556
rect 95770 4516 95812 4556
rect 95852 4516 95894 4556
rect 95934 4516 95976 4556
rect 95648 4507 96016 4516
rect 95500 4087 95540 4096
rect 95884 4136 95924 4145
rect 96076 4136 96116 5767
rect 96267 5732 96309 5741
rect 96267 5692 96268 5732
rect 96308 5692 96309 5732
rect 96267 5683 96309 5692
rect 95924 4096 96116 4136
rect 96268 4136 96308 5683
rect 95884 4087 95924 4096
rect 96268 4087 96308 4096
rect 96652 4136 96692 7783
rect 97035 7664 97077 7673
rect 97035 7624 97036 7664
rect 97076 7624 97077 7664
rect 97035 7615 97077 7624
rect 96652 4087 96692 4096
rect 97036 4136 97076 7615
rect 97131 4976 97173 4985
rect 97131 4936 97132 4976
rect 97172 4936 97173 4976
rect 97131 4927 97173 4936
rect 97132 4842 97172 4927
rect 97228 4145 97268 9379
rect 97899 9344 97941 9353
rect 97899 9304 97900 9344
rect 97940 9304 97941 9344
rect 97899 9295 97941 9304
rect 97611 9176 97653 9185
rect 97611 9136 97612 9176
rect 97652 9136 97653 9176
rect 97611 9127 97653 9136
rect 97419 8840 97461 8849
rect 97419 8800 97420 8840
rect 97460 8800 97461 8840
rect 97419 8791 97461 8800
rect 97324 4724 97364 4733
rect 97036 4087 97076 4096
rect 97227 4136 97269 4145
rect 97227 4096 97228 4136
rect 97268 4096 97269 4136
rect 97227 4087 97269 4096
rect 94923 4052 94965 4061
rect 94923 4012 94924 4052
rect 94964 4012 94965 4052
rect 97324 4052 97364 4684
rect 97420 4149 97460 8791
rect 97515 5648 97557 5657
rect 97515 5608 97516 5648
rect 97556 5608 97557 5648
rect 97515 5599 97557 5608
rect 97516 5514 97556 5599
rect 97420 4100 97460 4109
rect 97516 4724 97556 4733
rect 97324 4012 97460 4052
rect 94923 4003 94965 4012
rect 94539 3968 94581 3977
rect 94539 3928 94540 3968
rect 94580 3928 94581 3968
rect 94539 3919 94581 3928
rect 94731 3968 94773 3977
rect 94731 3928 94732 3968
rect 94772 3928 94773 3968
rect 94731 3919 94773 3928
rect 94924 3918 94964 4003
rect 95308 3968 95348 3977
rect 95692 3968 95732 3977
rect 95020 3928 95308 3968
rect 94408 3800 94776 3809
rect 94448 3760 94490 3800
rect 94530 3760 94572 3800
rect 94612 3760 94654 3800
rect 94694 3760 94736 3800
rect 94408 3751 94776 3760
rect 94348 3464 94388 3473
rect 94348 3305 94388 3424
rect 94731 3464 94773 3473
rect 94731 3424 94732 3464
rect 94772 3424 94773 3464
rect 94731 3415 94773 3424
rect 94732 3330 94772 3415
rect 95020 3380 95060 3928
rect 95308 3919 95348 3928
rect 95404 3928 95692 3968
rect 95115 3464 95157 3473
rect 95115 3424 95116 3464
rect 95156 3424 95157 3464
rect 95115 3415 95157 3424
rect 94828 3340 95060 3380
rect 94347 3296 94389 3305
rect 94347 3256 94348 3296
rect 94388 3256 94389 3296
rect 94347 3247 94389 3256
rect 94539 3212 94581 3221
rect 94539 3172 94540 3212
rect 94580 3172 94581 3212
rect 94539 3163 94581 3172
rect 94540 3078 94580 3163
rect 94828 2036 94868 3340
rect 95116 3330 95156 3415
rect 95404 3380 95444 3928
rect 95692 3919 95732 3928
rect 96076 3968 96116 3977
rect 96076 3809 96116 3928
rect 96171 3968 96213 3977
rect 96460 3968 96500 3977
rect 96171 3928 96172 3968
rect 96212 3928 96213 3968
rect 96171 3919 96213 3928
rect 96364 3928 96460 3968
rect 95595 3800 95637 3809
rect 95595 3760 95596 3800
rect 95636 3760 95637 3800
rect 95595 3751 95637 3760
rect 96075 3800 96117 3809
rect 96075 3760 96076 3800
rect 96116 3760 96117 3800
rect 96075 3751 96117 3760
rect 95500 3473 95540 3558
rect 95499 3464 95541 3473
rect 95499 3424 95500 3464
rect 95540 3424 95541 3464
rect 95499 3415 95541 3424
rect 95212 3340 95444 3380
rect 94156 1576 94292 1616
rect 94540 1996 94868 2036
rect 94924 3212 94964 3221
rect 94156 80 94196 1576
rect 94347 1532 94389 1541
rect 94347 1492 94348 1532
rect 94388 1492 94389 1532
rect 94347 1483 94389 1492
rect 94348 80 94388 1483
rect 94540 80 94580 1996
rect 94731 1784 94773 1793
rect 94731 1744 94732 1784
rect 94772 1744 94773 1784
rect 94731 1735 94773 1744
rect 94732 80 94772 1735
rect 94924 1625 94964 3172
rect 95212 1784 95252 3340
rect 95596 3296 95636 3751
rect 95883 3464 95925 3473
rect 95883 3424 95884 3464
rect 95924 3424 95925 3464
rect 95883 3415 95925 3424
rect 95884 3330 95924 3415
rect 95404 3256 95636 3296
rect 95020 1744 95252 1784
rect 95308 3212 95348 3221
rect 94923 1616 94965 1625
rect 94923 1576 94924 1616
rect 94964 1576 94965 1616
rect 94923 1567 94965 1576
rect 95020 1448 95060 1744
rect 95308 1709 95348 3172
rect 95307 1700 95349 1709
rect 95307 1660 95308 1700
rect 95348 1660 95349 1700
rect 95307 1651 95349 1660
rect 95115 1616 95157 1625
rect 95115 1576 95116 1616
rect 95156 1576 95157 1616
rect 95115 1567 95157 1576
rect 94924 1408 95060 1448
rect 94924 80 94964 1408
rect 95116 80 95156 1567
rect 95404 1532 95444 3256
rect 95692 3212 95732 3221
rect 95500 3172 95692 3212
rect 95500 1541 95540 3172
rect 95692 3163 95732 3172
rect 96076 3212 96116 3221
rect 95648 3044 96016 3053
rect 95688 3004 95730 3044
rect 95770 3004 95812 3044
rect 95852 3004 95894 3044
rect 95934 3004 95976 3044
rect 95648 2995 96016 3004
rect 95691 2876 95733 2885
rect 95691 2836 95692 2876
rect 95732 2836 95733 2876
rect 95691 2827 95733 2836
rect 95308 1492 95444 1532
rect 95499 1532 95541 1541
rect 95499 1492 95500 1532
rect 95540 1492 95541 1532
rect 95308 80 95348 1492
rect 95499 1483 95541 1492
rect 95499 1364 95541 1373
rect 95499 1324 95500 1364
rect 95540 1324 95541 1364
rect 95499 1315 95541 1324
rect 95500 80 95540 1315
rect 95692 80 95732 2827
rect 96076 1793 96116 3172
rect 96075 1784 96117 1793
rect 96075 1744 96076 1784
rect 96116 1744 96117 1784
rect 96075 1735 96117 1744
rect 95883 1700 95925 1709
rect 95883 1660 95884 1700
rect 95924 1660 95925 1700
rect 95883 1651 95925 1660
rect 95884 80 95924 1651
rect 96172 1616 96212 3919
rect 96268 3464 96308 3473
rect 96268 2717 96308 3424
rect 96364 2885 96404 3928
rect 96460 3919 96500 3928
rect 96843 3968 96885 3977
rect 97228 3968 97268 3977
rect 96843 3928 96844 3968
rect 96884 3928 96885 3968
rect 96843 3919 96885 3928
rect 97132 3928 97228 3968
rect 96844 3834 96884 3919
rect 96651 3464 96693 3473
rect 96651 3424 96652 3464
rect 96692 3424 96693 3464
rect 96651 3415 96693 3424
rect 97036 3464 97076 3473
rect 96652 3330 96692 3415
rect 97036 3380 97076 3424
rect 96940 3340 97076 3380
rect 96460 3212 96500 3221
rect 96363 2876 96405 2885
rect 96363 2836 96364 2876
rect 96404 2836 96405 2876
rect 96363 2827 96405 2836
rect 96267 2708 96309 2717
rect 96267 2668 96268 2708
rect 96308 2668 96309 2708
rect 96267 2659 96309 2668
rect 96460 1625 96500 3172
rect 96844 3212 96884 3221
rect 96651 2540 96693 2549
rect 96651 2500 96652 2540
rect 96692 2500 96693 2540
rect 96651 2491 96693 2500
rect 96076 1576 96212 1616
rect 96459 1616 96501 1625
rect 96459 1576 96460 1616
rect 96500 1576 96501 1616
rect 96076 80 96116 1576
rect 96459 1567 96501 1576
rect 96267 1532 96309 1541
rect 96267 1492 96268 1532
rect 96308 1492 96309 1532
rect 96267 1483 96309 1492
rect 96268 80 96308 1483
rect 96459 1448 96501 1457
rect 96459 1408 96460 1448
rect 96500 1408 96501 1448
rect 96459 1399 96501 1408
rect 96460 80 96500 1399
rect 96652 80 96692 2491
rect 96844 1373 96884 3172
rect 96940 2969 96980 3340
rect 97035 3212 97077 3221
rect 97035 3172 97036 3212
rect 97076 3172 97077 3212
rect 97035 3163 97077 3172
rect 96939 2960 96981 2969
rect 96939 2920 96940 2960
rect 96980 2920 96981 2960
rect 96939 2911 96981 2920
rect 96939 2036 96981 2045
rect 96939 1996 96940 2036
rect 96980 1996 96981 2036
rect 96939 1987 96981 1996
rect 96843 1364 96885 1373
rect 96843 1324 96844 1364
rect 96884 1324 96885 1364
rect 96843 1315 96885 1324
rect 96940 1196 96980 1987
rect 96844 1156 96980 1196
rect 96844 80 96884 1156
rect 97036 80 97076 3163
rect 97132 1457 97172 3928
rect 97228 3919 97268 3928
rect 97420 3641 97460 4012
rect 97419 3632 97461 3641
rect 97419 3592 97420 3632
rect 97460 3592 97461 3632
rect 97419 3583 97461 3592
rect 97419 3464 97461 3473
rect 97419 3424 97420 3464
rect 97460 3424 97461 3464
rect 97419 3415 97461 3424
rect 97323 3380 97365 3389
rect 97323 3340 97324 3380
rect 97364 3340 97365 3380
rect 97323 3331 97365 3340
rect 97228 3212 97268 3221
rect 97228 1709 97268 3172
rect 97227 1700 97269 1709
rect 97227 1660 97228 1700
rect 97268 1660 97269 1700
rect 97227 1651 97269 1660
rect 97324 1532 97364 3331
rect 97420 3330 97460 3415
rect 97516 2372 97556 4684
rect 97612 4136 97652 9127
rect 97900 5648 97940 9295
rect 98187 7748 98229 7757
rect 98187 7708 98188 7748
rect 98228 7708 98229 7748
rect 98187 7699 98229 7708
rect 97900 5599 97940 5608
rect 97708 5480 97748 5489
rect 98092 5480 98132 5489
rect 97748 5440 97844 5480
rect 97708 5431 97748 5440
rect 97707 4976 97749 4985
rect 97707 4936 97708 4976
rect 97748 4936 97749 4976
rect 97707 4927 97749 4936
rect 97708 4842 97748 4927
rect 97804 4313 97844 5440
rect 97996 5440 98092 5480
rect 97900 4724 97940 4733
rect 97803 4304 97845 4313
rect 97803 4264 97804 4304
rect 97844 4264 97845 4304
rect 97803 4255 97845 4264
rect 97804 4136 97844 4145
rect 97612 4096 97804 4136
rect 97804 4087 97844 4096
rect 97612 3968 97652 3977
rect 97652 3928 97748 3968
rect 97612 3919 97652 3928
rect 97228 1492 97364 1532
rect 97420 2332 97556 2372
rect 97612 3212 97652 3221
rect 97131 1448 97173 1457
rect 97131 1408 97132 1448
rect 97172 1408 97173 1448
rect 97131 1399 97173 1408
rect 97228 80 97268 1492
rect 97420 80 97460 2332
rect 97612 1541 97652 3172
rect 97708 2045 97748 3928
rect 97803 3464 97845 3473
rect 97803 3424 97804 3464
rect 97844 3424 97845 3464
rect 97803 3415 97845 3424
rect 97804 3330 97844 3415
rect 97900 2372 97940 4684
rect 97996 4136 98036 5440
rect 98092 5431 98132 5440
rect 98091 4976 98133 4985
rect 98091 4936 98092 4976
rect 98132 4936 98133 4976
rect 98091 4927 98133 4936
rect 98092 4842 98132 4927
rect 98188 4136 98228 7699
rect 98475 6488 98517 6497
rect 98475 6448 98476 6488
rect 98516 6448 98517 6488
rect 98475 6439 98517 6448
rect 98476 6354 98516 6439
rect 98668 6236 98708 6245
rect 98476 5648 98516 5657
rect 98476 5489 98516 5608
rect 98284 5480 98324 5489
rect 98475 5480 98517 5489
rect 98324 5440 98420 5480
rect 98284 5431 98324 5440
rect 98283 4724 98325 4733
rect 98283 4684 98284 4724
rect 98324 4684 98325 4724
rect 98283 4675 98325 4684
rect 98284 4590 98324 4675
rect 98380 4136 98420 5440
rect 98475 5440 98476 5480
rect 98516 5440 98517 5480
rect 98475 5431 98517 5440
rect 98476 4985 98516 5070
rect 98475 4976 98517 4985
rect 98475 4936 98476 4976
rect 98516 4936 98517 4976
rect 98475 4927 98517 4936
rect 98475 4724 98517 4733
rect 98475 4684 98476 4724
rect 98516 4684 98517 4724
rect 98475 4675 98517 4684
rect 97996 4096 98132 4136
rect 97996 3968 98036 3977
rect 97996 3389 98036 3928
rect 97995 3380 98037 3389
rect 97995 3340 97996 3380
rect 98036 3340 98037 3380
rect 97995 3331 98037 3340
rect 97996 3212 98036 3221
rect 97996 2633 98036 3172
rect 98092 3053 98132 4096
rect 98188 4087 98228 4096
rect 98284 4096 98420 4136
rect 98187 3716 98229 3725
rect 98187 3676 98188 3716
rect 98228 3676 98229 3716
rect 98187 3667 98229 3676
rect 98188 3464 98228 3667
rect 98188 3415 98228 3424
rect 98091 3044 98133 3053
rect 98091 3004 98092 3044
rect 98132 3004 98133 3044
rect 98091 2995 98133 3004
rect 97995 2624 98037 2633
rect 97995 2584 97996 2624
rect 98036 2584 98037 2624
rect 97995 2575 98037 2584
rect 98284 2540 98324 4096
rect 98379 3968 98421 3977
rect 98379 3928 98380 3968
rect 98420 3928 98421 3968
rect 98379 3919 98421 3928
rect 98380 3834 98420 3919
rect 98380 3221 98420 3306
rect 98379 3212 98421 3221
rect 98379 3172 98380 3212
rect 98420 3172 98421 3212
rect 98379 3163 98421 3172
rect 98379 3044 98421 3053
rect 98379 3004 98380 3044
rect 98420 3004 98421 3044
rect 98379 2995 98421 3004
rect 98188 2500 98324 2540
rect 97804 2332 97940 2372
rect 97995 2372 98037 2381
rect 97995 2332 97996 2372
rect 98036 2332 98037 2372
rect 97707 2036 97749 2045
rect 97707 1996 97708 2036
rect 97748 1996 97749 2036
rect 97707 1987 97749 1996
rect 97611 1532 97653 1541
rect 97611 1492 97612 1532
rect 97652 1492 97653 1532
rect 97611 1483 97653 1492
rect 97611 1364 97653 1373
rect 97611 1324 97612 1364
rect 97652 1324 97653 1364
rect 97611 1315 97653 1324
rect 97612 80 97652 1315
rect 97804 80 97844 2332
rect 97995 2323 98037 2332
rect 97996 80 98036 2323
rect 98188 80 98228 2500
rect 98380 80 98420 2995
rect 98476 2381 98516 4675
rect 98571 4136 98613 4145
rect 98571 4096 98572 4136
rect 98612 4096 98613 4136
rect 98571 4087 98613 4096
rect 98572 4002 98612 4087
rect 98571 3464 98613 3473
rect 98571 3424 98572 3464
rect 98612 3424 98613 3464
rect 98571 3415 98613 3424
rect 98572 3330 98612 3415
rect 98668 2540 98708 6196
rect 98955 4304 98997 4313
rect 98955 4264 98956 4304
rect 98996 4264 98997 4304
rect 98955 4255 98997 4264
rect 98763 3968 98805 3977
rect 98763 3928 98764 3968
rect 98804 3928 98805 3968
rect 98763 3919 98805 3928
rect 98572 2500 98708 2540
rect 98475 2372 98517 2381
rect 98475 2332 98476 2372
rect 98516 2332 98517 2372
rect 98475 2323 98517 2332
rect 98572 80 98612 2500
rect 98764 1373 98804 3919
rect 98859 3632 98901 3641
rect 98859 3592 98860 3632
rect 98900 3592 98901 3632
rect 98859 3583 98901 3592
rect 98763 1364 98805 1373
rect 98763 1324 98764 1364
rect 98804 1324 98805 1364
rect 98763 1315 98805 1324
rect 98860 1196 98900 3583
rect 98764 1156 98900 1196
rect 98764 80 98804 1156
rect 98956 80 98996 4255
rect 88820 64 88840 80
rect 88760 0 88840 64
rect 88952 0 89032 80
rect 89144 0 89224 80
rect 89336 0 89416 80
rect 89528 0 89608 80
rect 89720 0 89800 80
rect 89912 0 89992 80
rect 90104 0 90184 80
rect 90296 0 90376 80
rect 90488 0 90568 80
rect 90680 0 90760 80
rect 90872 0 90952 80
rect 91064 0 91144 80
rect 91256 0 91336 80
rect 91448 0 91528 80
rect 91640 0 91720 80
rect 91832 0 91912 80
rect 92024 0 92104 80
rect 92216 0 92296 80
rect 92408 0 92488 80
rect 92600 0 92680 80
rect 92792 0 92872 80
rect 92984 0 93064 80
rect 93176 0 93256 80
rect 93368 0 93448 80
rect 93560 0 93640 80
rect 93752 0 93832 80
rect 93944 0 94024 80
rect 94136 0 94216 80
rect 94328 0 94408 80
rect 94520 0 94600 80
rect 94712 0 94792 80
rect 94904 0 94984 80
rect 95096 0 95176 80
rect 95288 0 95368 80
rect 95480 0 95560 80
rect 95672 0 95752 80
rect 95864 0 95944 80
rect 96056 0 96136 80
rect 96248 0 96328 80
rect 96440 0 96520 80
rect 96632 0 96712 80
rect 96824 0 96904 80
rect 97016 0 97096 80
rect 97208 0 97288 80
rect 97400 0 97480 80
rect 97592 0 97672 80
rect 97784 0 97864 80
rect 97976 0 98056 80
rect 98168 0 98248 80
rect 98360 0 98440 80
rect 98552 0 98632 80
rect 98744 0 98824 80
rect 98936 0 99016 80
<< via2 >>
rect 6220 11908 6260 11948
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 11980 10984 12020 11024
rect 10732 10816 10772 10856
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 7372 10144 7412 10184
rect 3436 9976 3476 10016
rect 3052 8800 3092 8840
rect 1996 8128 2036 8168
rect 1420 6448 1460 6488
rect 1708 5608 1748 5648
rect 1132 5440 1172 5480
rect 1036 3340 1076 3380
rect 1228 3424 1268 3464
rect 1900 5440 1940 5480
rect 1612 4852 1652 4892
rect 1708 4768 1748 4808
rect 1612 3424 1652 3464
rect 1420 3172 1460 3212
rect 1612 3172 1652 3212
rect 1612 2500 1652 2540
rect 2380 7708 2420 7748
rect 2092 5608 2132 5648
rect 2092 4936 2132 4976
rect 1996 3424 2036 3464
rect 1804 2500 1844 2540
rect 1708 1996 1748 2036
rect 1996 1996 2036 2036
rect 2764 6364 2804 6404
rect 2476 4936 2516 4976
rect 2380 3424 2420 3464
rect 2188 3172 2228 3212
rect 2380 3172 2420 3212
rect 2092 1912 2132 1952
rect 2668 4180 2708 4220
rect 2572 3340 2612 3380
rect 2572 3172 2612 3212
rect 2572 2332 2612 2372
rect 2380 2080 2420 2120
rect 2380 1912 2420 1952
rect 3148 6616 3188 6656
rect 3340 5440 3380 5480
rect 2956 2500 2996 2540
rect 2860 1156 2900 1196
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 6220 9472 6260 9512
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6124 8716 6164 8756
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5356 7120 5396 7160
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4780 6112 4820 6152
rect 4108 5692 4148 5732
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3820 5104 3860 5144
rect 4012 3928 4052 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3340 3424 3380 3464
rect 3532 3424 3572 3464
rect 3244 3088 3284 3128
rect 3628 3172 3668 3212
rect 3532 3088 3572 3128
rect 3340 2080 3380 2120
rect 3148 1408 3188 1448
rect 3052 1240 3092 1280
rect 3148 1156 3188 1196
rect 3436 1156 3476 1196
rect 4204 5020 4244 5060
rect 4588 4096 4628 4136
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 5068 4348 5108 4388
rect 4204 3928 4244 3968
rect 3724 1492 3764 1532
rect 4300 3424 4340 3464
rect 4108 1576 4148 1616
rect 4108 1240 4148 1280
rect 4492 1660 4532 1700
rect 4684 3760 4724 3800
rect 4684 3172 4724 3212
rect 5740 6868 5780 6908
rect 5452 6196 5492 6236
rect 5452 4348 5492 4388
rect 6508 6952 6548 6992
rect 6220 5020 6260 5060
rect 6892 6280 6932 6320
rect 7468 9892 7508 9932
rect 7372 6112 7412 6152
rect 7372 5356 7412 5396
rect 7276 4096 7316 4136
rect 4876 3172 4916 3212
rect 5260 3172 5300 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 5452 2416 5492 2456
rect 4684 1744 4724 1784
rect 4492 1156 4532 1196
rect 4876 1492 4916 1532
rect 5260 1576 5300 1616
rect 5548 1912 5588 1952
rect 5740 3172 5780 3212
rect 5836 2332 5876 2372
rect 5740 1996 5780 2036
rect 6220 2920 6260 2960
rect 5836 1912 5876 1952
rect 6028 1912 6068 1952
rect 5644 1828 5684 1868
rect 5644 1660 5684 1700
rect 6028 1744 6068 1784
rect 6412 1996 6452 2036
rect 6316 1660 6356 1700
rect 6796 1996 6836 2036
rect 6988 3424 7028 3464
rect 7180 2164 7220 2204
rect 6796 1828 6836 1868
rect 6700 1744 6740 1784
rect 7180 1912 7220 1952
rect 9196 9388 9236 9428
rect 7564 8968 7604 9008
rect 8812 8800 8852 8840
rect 8428 8212 8468 8252
rect 7564 7708 7604 7748
rect 8044 7708 8084 7748
rect 7468 5104 7508 5144
rect 7660 4264 7700 4304
rect 8812 8128 8852 8168
rect 8908 7876 8948 7916
rect 9100 7792 9140 7832
rect 9004 6112 9044 6152
rect 8908 5272 8948 5312
rect 8812 4936 8852 4976
rect 7372 3760 7412 3800
rect 7372 3088 7412 3128
rect 7372 2920 7412 2960
rect 7372 2080 7412 2120
rect 7756 3256 7796 3296
rect 7564 3172 7604 3212
rect 7948 2332 7988 2372
rect 7564 1660 7604 1700
rect 7948 1996 7988 2036
rect 8140 3424 8180 3464
rect 8524 3172 8564 3212
rect 8428 3004 8468 3044
rect 8332 2584 8372 2624
rect 8332 2164 8372 2204
rect 9580 9304 9620 9344
rect 9484 8296 9524 8336
rect 9292 8128 9332 8168
rect 9292 7876 9332 7916
rect 9196 5188 9236 5228
rect 9292 5104 9332 5144
rect 9196 4684 9236 4724
rect 9772 9220 9812 9260
rect 9676 8716 9716 8756
rect 9868 7960 9908 8000
rect 9676 7876 9716 7916
rect 10060 8716 10100 8756
rect 10156 8296 10196 8336
rect 10060 8128 10100 8168
rect 10252 7960 10292 8000
rect 10060 7372 10100 7412
rect 9484 7036 9524 7076
rect 9676 7204 9716 7244
rect 9868 7204 9908 7244
rect 10156 7288 10196 7328
rect 10636 8716 10676 8756
rect 10636 7960 10676 8000
rect 10348 7624 10388 7664
rect 10444 7540 10484 7580
rect 10636 7540 10676 7580
rect 10348 7288 10388 7328
rect 9964 7036 10004 7076
rect 9772 6952 9812 6992
rect 9676 5860 9716 5900
rect 9580 5608 9620 5648
rect 9580 5188 9620 5228
rect 9388 4600 9428 4640
rect 9100 2332 9140 2372
rect 8716 2164 8756 2204
rect 9196 1324 9236 1364
rect 10060 6700 10100 6740
rect 10252 6532 10292 6572
rect 10156 6448 10196 6488
rect 10252 4852 10292 4892
rect 10540 7204 10580 7244
rect 10828 10732 10868 10772
rect 11500 10732 11540 10772
rect 11788 10732 11828 10772
rect 10924 10564 10964 10604
rect 11212 10480 11252 10520
rect 11404 10228 11444 10268
rect 11404 9556 11444 9596
rect 11308 8884 11348 8924
rect 11116 8716 11156 8756
rect 11308 8548 11348 8588
rect 11020 8380 11060 8420
rect 10924 8296 10964 8336
rect 10828 7288 10868 7328
rect 10444 6532 10484 6572
rect 10444 6364 10484 6404
rect 10348 4768 10388 4808
rect 10732 4264 10772 4304
rect 10540 4096 10580 4136
rect 11020 7876 11060 7916
rect 11212 7204 11252 7244
rect 10924 6364 10964 6404
rect 11212 6952 11252 6992
rect 11116 6280 11156 6320
rect 11596 10648 11636 10688
rect 11596 10228 11636 10268
rect 12172 10900 12212 10940
rect 12364 10648 12404 10688
rect 12364 10480 12404 10520
rect 12172 10396 12212 10436
rect 12076 10228 12116 10268
rect 11788 10060 11828 10100
rect 11692 9556 11732 9596
rect 11692 9136 11732 9176
rect 11788 8884 11828 8924
rect 11596 8800 11636 8840
rect 11500 8716 11540 8756
rect 11980 8968 12020 9008
rect 11884 8716 11924 8756
rect 11692 7792 11732 7832
rect 11596 7708 11636 7748
rect 11692 7456 11732 7496
rect 11212 5020 11252 5060
rect 11020 4180 11060 4220
rect 11116 4096 11156 4136
rect 9484 2500 9524 2540
rect 9388 988 9428 1028
rect 9676 2164 9716 2204
rect 9580 1576 9620 1616
rect 10060 3424 10100 3464
rect 9868 1660 9908 1700
rect 10444 3088 10484 3128
rect 10252 1492 10292 1532
rect 10252 1324 10292 1364
rect 9676 988 9716 1028
rect 10828 3256 10868 3296
rect 10636 1744 10676 1784
rect 10636 1576 10676 1616
rect 11596 5188 11636 5228
rect 11020 1828 11060 1868
rect 11020 1660 11060 1700
rect 11980 8128 12020 8168
rect 12748 10900 12788 10940
rect 12556 10396 12596 10436
rect 14572 10732 14612 10772
rect 15148 10732 15188 10772
rect 14476 10564 14516 10604
rect 12940 10396 12980 10436
rect 14956 10648 14996 10688
rect 14764 10564 14804 10604
rect 14572 10228 14612 10268
rect 12844 10144 12884 10184
rect 14476 10144 14516 10184
rect 12748 10060 12788 10100
rect 12364 9052 12404 9092
rect 12460 8884 12500 8924
rect 13036 9220 13076 9260
rect 12556 8800 12596 8840
rect 12268 8716 12308 8756
rect 12460 8716 12500 8756
rect 12652 8716 12692 8756
rect 12076 7960 12116 8000
rect 12076 7792 12116 7832
rect 12172 7708 12212 7748
rect 11884 7456 11924 7496
rect 11884 7288 11924 7328
rect 11788 6952 11828 6992
rect 12460 8044 12500 8084
rect 12364 7876 12404 7916
rect 12556 7456 12596 7496
rect 12940 8212 12980 8252
rect 12748 8128 12788 8168
rect 12940 7876 12980 7916
rect 12748 7456 12788 7496
rect 12268 7120 12308 7160
rect 13324 8716 13364 8756
rect 13132 8128 13172 8168
rect 13708 8632 13748 8672
rect 13516 8128 13556 8168
rect 13324 8044 13364 8084
rect 12844 7120 12884 7160
rect 12076 6952 12116 6992
rect 12268 6532 12308 6572
rect 11980 4936 12020 4976
rect 12556 6448 12596 6488
rect 12556 6196 12596 6236
rect 12748 6952 12788 6992
rect 12652 4684 12692 4724
rect 12364 4600 12404 4640
rect 11404 1660 11444 1700
rect 11404 1492 11444 1532
rect 11980 3592 12020 3632
rect 11788 1912 11828 1952
rect 11788 1744 11828 1784
rect 13132 7120 13172 7160
rect 13036 4432 13076 4472
rect 12172 2248 12212 2288
rect 12172 1828 12212 1868
rect 12556 1660 12596 1700
rect 12460 484 12500 524
rect 12748 1660 12788 1700
rect 13324 7624 13364 7664
rect 13228 6364 13268 6404
rect 13708 7624 13748 7664
rect 13612 7372 13652 7412
rect 13708 7288 13748 7328
rect 13612 7204 13652 7244
rect 13420 6952 13460 6992
rect 13708 6112 13748 6152
rect 13900 4936 13940 4976
rect 14476 9136 14516 9176
rect 14380 8548 14420 8588
rect 14188 8128 14228 8168
rect 14284 7792 14324 7832
rect 14188 7372 14228 7412
rect 12940 1912 12980 1952
rect 12844 568 12884 608
rect 13132 1660 13172 1700
rect 13036 1492 13076 1532
rect 13804 4348 13844 4388
rect 13516 3004 13556 3044
rect 13324 2248 13364 2288
rect 13228 1240 13268 1280
rect 13132 736 13172 776
rect 13132 568 13172 608
rect 13420 1576 13460 1616
rect 13612 2500 13652 2540
rect 13900 3088 13940 3128
rect 13900 2836 13940 2876
rect 13708 1240 13748 1280
rect 14668 9388 14708 9428
rect 14860 10060 14900 10100
rect 14572 8800 14612 8840
rect 15724 10816 15764 10856
rect 15628 10732 15668 10772
rect 15532 10648 15572 10688
rect 15532 10312 15572 10352
rect 15340 10228 15380 10268
rect 15148 9808 15188 9848
rect 15148 9640 15188 9680
rect 14956 8800 14996 8840
rect 14476 6112 14516 6152
rect 14764 6112 14804 6152
rect 14668 4936 14708 4976
rect 14188 3928 14228 3968
rect 14092 3172 14132 3212
rect 14668 4516 14708 4556
rect 14572 4180 14612 4220
rect 14380 3340 14420 3380
rect 14380 3172 14420 3212
rect 13996 1324 14036 1364
rect 13804 988 13844 1028
rect 13900 484 13940 524
rect 14284 2416 14324 2456
rect 14764 4096 14804 4136
rect 14764 3928 14804 3968
rect 15436 10060 15476 10100
rect 15724 10228 15764 10268
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 28396 11404 28436 11444
rect 19564 11068 19604 11108
rect 21196 11068 21236 11108
rect 24364 11068 24404 11108
rect 19276 10984 19316 11024
rect 17452 10900 17492 10940
rect 18604 10732 18644 10772
rect 16300 10396 16340 10436
rect 15916 10228 15956 10268
rect 16108 10228 16148 10268
rect 19084 10648 19124 10688
rect 18796 10396 18836 10436
rect 19180 10480 19220 10520
rect 17644 10144 17684 10184
rect 16204 10060 16244 10100
rect 15916 9388 15956 9428
rect 15436 9304 15476 9344
rect 15532 8884 15572 8924
rect 15436 8800 15476 8840
rect 15244 8716 15284 8756
rect 15724 8548 15764 8588
rect 15244 6700 15284 6740
rect 15148 6532 15188 6572
rect 15052 6364 15092 6404
rect 15148 6196 15188 6236
rect 15052 4768 15092 4808
rect 15340 5776 15380 5816
rect 15532 6868 15572 6908
rect 15628 6532 15668 6572
rect 15820 6616 15860 6656
rect 16300 9640 16340 9680
rect 16108 9388 16148 9428
rect 16300 8800 16340 8840
rect 16780 8800 16820 8840
rect 16588 6868 16628 6908
rect 16204 6700 16244 6740
rect 16396 6532 16436 6572
rect 15820 6364 15860 6404
rect 15724 6196 15764 6236
rect 16012 6364 16052 6404
rect 16300 6364 16340 6404
rect 16108 6280 16148 6320
rect 16397 6280 16437 6320
rect 16012 6028 16052 6068
rect 15916 5944 15956 5984
rect 15724 5608 15764 5648
rect 15724 5104 15764 5144
rect 15340 5020 15380 5060
rect 15535 5020 15575 5060
rect 15436 4852 15476 4892
rect 16108 5776 16148 5816
rect 16684 6028 16724 6068
rect 16396 5944 16436 5984
rect 16108 5272 16148 5312
rect 16300 5188 16340 5228
rect 16108 5020 16148 5060
rect 15052 3844 15092 3884
rect 15148 3760 15188 3800
rect 15052 3676 15092 3716
rect 14764 3340 14804 3380
rect 14476 1660 14516 1700
rect 14476 1492 14516 1532
rect 14380 1072 14420 1112
rect 15148 3256 15188 3296
rect 15052 1576 15092 1616
rect 14860 1492 14900 1532
rect 14860 1324 14900 1364
rect 14764 1240 14804 1280
rect 15244 1576 15284 1616
rect 15628 4684 15668 4724
rect 15436 3676 15476 3716
rect 15436 3172 15476 3212
rect 15724 4264 15764 4304
rect 16492 5692 16532 5732
rect 16492 5440 16532 5480
rect 17164 7204 17204 7244
rect 17260 6280 17300 6320
rect 17068 5944 17108 5984
rect 16972 5860 17012 5900
rect 16876 5776 16916 5816
rect 16492 5104 16532 5144
rect 16108 3928 16148 3968
rect 15628 3760 15668 3800
rect 15916 3760 15956 3800
rect 15724 3676 15764 3716
rect 15532 2584 15572 2624
rect 15820 3424 15860 3464
rect 15916 3340 15956 3380
rect 15916 3172 15956 3212
rect 15628 1324 15668 1364
rect 15436 1240 15476 1280
rect 15340 1156 15380 1196
rect 15628 988 15668 1028
rect 16780 5020 16820 5060
rect 17164 5860 17204 5900
rect 17452 5944 17492 5984
rect 17260 5692 17300 5732
rect 19180 10144 19220 10184
rect 18988 10060 19028 10100
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19180 9640 19220 9680
rect 18700 9472 18740 9512
rect 18988 9388 19028 9428
rect 18412 8968 18452 9008
rect 17836 8296 17876 8336
rect 17836 8044 17876 8084
rect 18028 7876 18068 7916
rect 18220 7876 18260 7916
rect 19564 10816 19604 10856
rect 19948 10900 19988 10940
rect 19660 10732 19700 10772
rect 19948 10564 19988 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 19852 10480 19892 10520
rect 19372 10060 19412 10100
rect 19948 10228 19988 10268
rect 19756 10060 19796 10100
rect 20332 10312 20372 10352
rect 20131 10060 20171 10100
rect 19564 9724 19604 9764
rect 19468 9472 19508 9512
rect 19372 9388 19412 9428
rect 19468 9304 19508 9344
rect 19948 9388 19988 9428
rect 18700 8800 18740 8840
rect 19084 8800 19124 8840
rect 18604 8716 18644 8756
rect 18796 8632 18836 8672
rect 19372 8632 19412 8672
rect 18604 8380 18644 8420
rect 19276 8380 19316 8420
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 18796 8128 18836 8168
rect 19180 8128 19220 8168
rect 17932 7792 17972 7832
rect 17740 6868 17780 6908
rect 18220 6616 18260 6656
rect 18604 7876 18644 7916
rect 18412 7456 18452 7496
rect 18988 7876 19028 7916
rect 18796 7792 18836 7832
rect 19564 8464 19604 8504
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 19564 7960 19604 8000
rect 19372 7876 19412 7916
rect 18892 7708 18932 7748
rect 18892 7540 18932 7580
rect 18700 7372 18740 7412
rect 19276 7792 19316 7832
rect 19276 7456 19316 7496
rect 19084 7036 19124 7076
rect 18796 6952 18836 6992
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 18316 6532 18356 6572
rect 17260 5524 17300 5564
rect 17164 5356 17204 5396
rect 17740 5356 17780 5396
rect 18220 6196 18260 6236
rect 18316 5944 18356 5984
rect 18124 5692 18164 5732
rect 17836 5104 17876 5144
rect 17356 4852 17396 4892
rect 17548 4852 17588 4892
rect 16588 3928 16628 3968
rect 16396 2416 16436 2456
rect 16300 1240 16340 1280
rect 15916 316 15956 356
rect 16204 1072 16244 1112
rect 16588 2668 16628 2708
rect 16876 3928 16916 3968
rect 16780 3424 16820 3464
rect 16684 2584 16724 2624
rect 16492 1660 16532 1700
rect 16588 1156 16628 1196
rect 16492 400 16532 440
rect 16684 904 16724 944
rect 16972 3424 17012 3464
rect 16972 2416 17012 2456
rect 16876 1156 16916 1196
rect 16780 568 16820 608
rect 16780 400 16820 440
rect 17164 4600 17204 4640
rect 17356 4600 17396 4640
rect 17548 4432 17588 4472
rect 17740 4600 17780 4640
rect 17644 4180 17684 4220
rect 17644 4012 17684 4052
rect 17164 3424 17204 3464
rect 17164 3172 17204 3212
rect 17548 3760 17588 3800
rect 17356 3424 17396 3464
rect 17740 3844 17780 3884
rect 17260 3088 17300 3128
rect 17548 2584 17588 2624
rect 18220 5104 18260 5144
rect 18700 6448 18740 6488
rect 19468 6700 19508 6740
rect 20044 7960 20084 8000
rect 20428 7876 20468 7916
rect 19756 7624 19796 7664
rect 19948 7792 19988 7832
rect 19852 7540 19892 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 19468 6532 19508 6572
rect 18604 6196 18644 6236
rect 18892 6196 18932 6236
rect 19180 6112 19220 6152
rect 19084 6028 19124 6068
rect 18604 5692 18644 5732
rect 18796 5692 18836 5732
rect 19084 5776 19124 5816
rect 19180 5692 19220 5732
rect 18508 5356 18548 5396
rect 18892 5440 18932 5480
rect 19084 5440 19124 5480
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18892 5104 18932 5144
rect 18604 5020 18644 5060
rect 18796 4852 18836 4892
rect 18316 4684 18356 4724
rect 18508 4684 18548 4724
rect 18124 4516 18164 4556
rect 18124 4096 18164 4136
rect 17164 1492 17204 1532
rect 17068 820 17108 860
rect 17356 1156 17396 1196
rect 17740 1576 17780 1616
rect 17932 820 17972 860
rect 18220 1324 18260 1364
rect 18124 1240 18164 1280
rect 18028 652 18068 692
rect 19185 4936 19225 4976
rect 19084 4768 19124 4808
rect 18988 4600 19028 4640
rect 19180 4432 19220 4472
rect 18604 3508 18644 3548
rect 18508 3424 18548 3464
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19372 6196 19412 6236
rect 19660 6364 19700 6404
rect 20620 9388 20660 9428
rect 24076 10816 24116 10856
rect 21292 10732 21332 10772
rect 21484 10732 21524 10772
rect 21292 10396 21332 10436
rect 23404 10648 23444 10688
rect 23884 10648 23924 10688
rect 21676 10480 21716 10520
rect 21484 10312 21524 10352
rect 21580 9892 21620 9932
rect 21964 9472 22004 9512
rect 20620 7792 20660 7832
rect 20812 7792 20852 7832
rect 21004 7036 21044 7076
rect 20716 6952 20756 6992
rect 19756 6280 19796 6320
rect 19564 5860 19604 5900
rect 19372 5188 19412 5228
rect 19564 5440 19604 5480
rect 19372 4684 19412 4724
rect 18892 3508 18932 3548
rect 18316 1240 18356 1280
rect 18604 1912 18644 1952
rect 19468 4264 19508 4304
rect 19564 4180 19604 4220
rect 19372 3508 19412 3548
rect 19276 3424 19316 3464
rect 19852 6196 19892 6236
rect 20428 6196 20468 6236
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 19948 5860 19988 5900
rect 19756 5776 19796 5816
rect 20332 5776 20372 5816
rect 20236 5608 20276 5648
rect 19756 5524 19796 5564
rect 20140 5524 20180 5564
rect 20524 5692 20564 5732
rect 20332 5440 20372 5480
rect 20524 5440 20564 5480
rect 19948 5020 19988 5060
rect 20332 4936 20372 4976
rect 20121 4852 20161 4892
rect 19948 4684 19988 4724
rect 19852 4600 19892 4640
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20332 4264 20372 4304
rect 20145 4180 20185 4220
rect 20524 4180 20564 4220
rect 19756 3928 19796 3968
rect 19948 3928 19988 3968
rect 20428 3844 20468 3884
rect 20044 3424 20084 3464
rect 20524 3508 20564 3548
rect 20716 5776 20756 5816
rect 20716 5272 20756 5312
rect 21100 6700 21140 6740
rect 20908 5188 20948 5228
rect 20908 4852 20948 4892
rect 20716 4684 20756 4724
rect 20716 4516 20756 4556
rect 20812 4432 20852 4472
rect 19084 1576 19124 1616
rect 18796 1072 18836 1112
rect 18700 988 18740 1028
rect 19084 904 19124 944
rect 18892 316 18932 356
rect 19660 3172 19700 3212
rect 19468 1492 19508 1532
rect 19468 568 19508 608
rect 20236 3172 20276 3212
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20044 2416 20084 2456
rect 19852 1324 19892 1364
rect 19852 652 19892 692
rect 20236 1240 20276 1280
rect 20620 1828 20660 1868
rect 20620 1072 20660 1112
rect 20908 3676 20948 3716
rect 21484 6196 21524 6236
rect 21388 5188 21428 5228
rect 21292 4852 21332 4892
rect 21100 4600 21140 4640
rect 21292 4516 21332 4556
rect 21196 4348 21236 4388
rect 21196 4180 21236 4220
rect 21100 4012 21140 4052
rect 21484 4768 21524 4808
rect 21484 4432 21524 4472
rect 21484 4180 21524 4220
rect 21388 3844 21428 3884
rect 21196 3424 21236 3464
rect 20812 3256 20852 3296
rect 20716 904 20756 944
rect 21004 3172 21044 3212
rect 20908 3088 20948 3128
rect 20908 1156 20948 1196
rect 21004 988 21044 1028
rect 22348 8548 22388 8588
rect 22636 7876 22676 7916
rect 23308 7876 23348 7916
rect 23020 7792 23060 7832
rect 23212 7792 23252 7832
rect 22540 7624 22580 7664
rect 22636 7372 22676 7412
rect 22828 7372 22868 7412
rect 23020 7372 23060 7412
rect 22732 7204 22772 7244
rect 22924 7204 22964 7244
rect 23116 7204 23156 7244
rect 22924 6364 22964 6404
rect 23212 7120 23252 7160
rect 23308 7036 23348 7076
rect 23788 10564 23828 10604
rect 23980 10060 24020 10100
rect 23788 9724 23828 9764
rect 24460 10984 24500 11024
rect 24364 10816 24404 10856
rect 24748 10900 24788 10940
rect 25420 11068 25460 11108
rect 24844 10396 24884 10436
rect 24172 10060 24212 10100
rect 24076 9640 24116 9680
rect 24364 9892 24404 9932
rect 24268 9556 24308 9596
rect 24172 9388 24212 9428
rect 23500 9304 23540 9344
rect 23404 6700 23444 6740
rect 23212 6364 23252 6404
rect 23404 6364 23444 6404
rect 23020 6028 23060 6068
rect 22924 5944 22964 5984
rect 23116 5944 23156 5984
rect 22732 5524 22772 5564
rect 21964 5020 22004 5060
rect 22444 5020 22484 5060
rect 21868 4852 21908 4892
rect 21676 4432 21716 4472
rect 21580 3508 21620 3548
rect 21484 2500 21524 2540
rect 22252 4852 22292 4892
rect 22924 5272 22964 5312
rect 22828 5104 22868 5144
rect 22540 4768 22580 4808
rect 23020 5104 23060 5144
rect 22348 4684 22388 4724
rect 22828 4684 22868 4724
rect 22252 4600 22292 4640
rect 22156 4516 22196 4556
rect 21868 4180 21908 4220
rect 21772 3508 21812 3548
rect 22060 3844 22100 3884
rect 22828 4432 22868 4472
rect 22732 4264 22772 4304
rect 22252 4180 22292 4220
rect 22636 4180 22676 4220
rect 22924 4180 22964 4220
rect 22540 3844 22580 3884
rect 22444 3760 22484 3800
rect 21964 3424 22004 3464
rect 21580 1576 21620 1616
rect 21484 988 21524 1028
rect 21964 2164 22004 2204
rect 21868 1660 21908 1700
rect 22348 3592 22388 3632
rect 23308 6028 23348 6068
rect 23404 5860 23444 5900
rect 23308 5692 23348 5732
rect 24268 9304 24308 9344
rect 24748 10228 24788 10268
rect 24652 9472 24692 9512
rect 24556 9388 24596 9428
rect 24460 9052 24500 9092
rect 25228 10900 25268 10940
rect 25420 10900 25460 10940
rect 33928 11320 33968 11360
rect 34010 11320 34050 11360
rect 34092 11320 34132 11360
rect 34174 11320 34214 11360
rect 34256 11320 34296 11360
rect 25132 10732 25172 10772
rect 29260 10648 29300 10688
rect 25420 10480 25460 10520
rect 25324 9808 25364 9848
rect 27724 9556 27764 9596
rect 25228 9388 25268 9428
rect 25324 9052 25364 9092
rect 25036 8968 25076 9008
rect 24940 8884 24980 8924
rect 24076 8716 24116 8756
rect 24364 8716 24404 8756
rect 24172 8380 24212 8420
rect 23596 7876 23636 7916
rect 24076 7876 24116 7916
rect 24268 7540 24308 7580
rect 24172 7456 24212 7496
rect 23596 7288 23636 7328
rect 24076 7204 24116 7244
rect 25036 8800 25076 8840
rect 24556 8716 24596 8756
rect 24940 8716 24980 8756
rect 24748 8632 24788 8672
rect 24556 8128 24596 8168
rect 24556 7876 24596 7916
rect 24748 7876 24788 7916
rect 24460 7372 24500 7412
rect 23788 6616 23828 6656
rect 23788 6448 23828 6488
rect 23596 6364 23636 6404
rect 24364 7204 24404 7244
rect 24460 7036 24500 7076
rect 24364 6952 24404 6992
rect 24268 6868 24308 6908
rect 24172 6784 24212 6824
rect 24076 6364 24116 6404
rect 23692 5860 23732 5900
rect 23980 5860 24020 5900
rect 23980 5692 24020 5732
rect 24268 6196 24308 6236
rect 24556 6700 24596 6740
rect 24748 7288 24788 7328
rect 24748 6952 24788 6992
rect 24460 6196 24500 6236
rect 23788 5440 23828 5480
rect 23212 4684 23252 4724
rect 23116 3676 23156 3716
rect 22732 3592 22772 3632
rect 22636 3508 22676 3548
rect 22252 1996 22292 2036
rect 21964 1492 22004 1532
rect 22156 1492 22196 1532
rect 22348 1324 22388 1364
rect 22156 1156 22196 1196
rect 22540 1072 22580 1112
rect 22540 904 22580 944
rect 23116 3424 23156 3464
rect 23116 3172 23156 3212
rect 23020 1828 23060 1868
rect 22924 1744 22964 1784
rect 23596 5020 23636 5060
rect 24364 5188 24404 5228
rect 24172 4852 24212 4892
rect 23404 4768 23444 4808
rect 23788 4768 23828 4808
rect 23404 4264 23444 4304
rect 23596 4180 23636 4220
rect 23500 3424 23540 3464
rect 23308 3340 23348 3380
rect 23788 4180 23828 4220
rect 24652 6112 24692 6152
rect 24748 6028 24788 6068
rect 23980 4180 24020 4220
rect 23980 4012 24020 4052
rect 23884 3592 23924 3632
rect 24364 4600 24404 4640
rect 24268 4348 24308 4388
rect 24172 4180 24212 4220
rect 24268 4096 24308 4136
rect 24652 4936 24692 4976
rect 24556 4852 24596 4892
rect 24748 4516 24788 4556
rect 24652 4348 24692 4388
rect 24556 3928 24596 3968
rect 24652 3760 24692 3800
rect 25420 8716 25460 8756
rect 26860 8800 26900 8840
rect 25612 8464 25652 8504
rect 25324 8296 25364 8336
rect 25132 8212 25172 8252
rect 25132 7960 25172 8000
rect 24940 7876 24980 7916
rect 25900 8044 25940 8084
rect 25516 7876 25556 7916
rect 25708 7876 25748 7916
rect 25036 7792 25076 7832
rect 25228 7708 25268 7748
rect 25132 7204 25172 7244
rect 25036 7036 25076 7076
rect 25036 6700 25076 6740
rect 25132 6616 25172 6656
rect 25036 6364 25076 6404
rect 25708 7540 25748 7580
rect 25036 5356 25076 5396
rect 25132 5188 25172 5228
rect 25132 5020 25172 5060
rect 24940 4852 24980 4892
rect 25324 6364 25364 6404
rect 25516 6364 25556 6404
rect 26476 7792 26516 7832
rect 25420 5104 25460 5144
rect 25324 4852 25364 4892
rect 25228 4768 25268 4808
rect 25516 4768 25556 4808
rect 25036 4684 25076 4724
rect 25324 4684 25364 4724
rect 25132 3844 25172 3884
rect 25516 4264 25556 4304
rect 25900 5020 25940 5060
rect 26188 6364 26228 6404
rect 26380 6364 26420 6404
rect 26188 5944 26228 5984
rect 26380 6196 26420 6236
rect 23692 2500 23732 2540
rect 23308 1576 23348 1616
rect 22924 820 22964 860
rect 22828 736 22868 776
rect 23692 1660 23732 1700
rect 23500 1240 23540 1280
rect 23404 1156 23444 1196
rect 23500 988 23540 1028
rect 23884 1492 23924 1532
rect 24076 1324 24116 1364
rect 24076 1156 24116 1196
rect 24748 1744 24788 1784
rect 24460 1492 24500 1532
rect 24652 1240 24692 1280
rect 25420 3592 25460 3632
rect 25420 3424 25460 3464
rect 25228 3172 25268 3212
rect 25228 2416 25268 2456
rect 25132 2248 25172 2288
rect 24844 1660 24884 1700
rect 25036 1576 25076 1616
rect 24460 1072 24500 1112
rect 25420 1324 25460 1364
rect 25708 4096 25748 4136
rect 25612 2500 25652 2540
rect 25516 1240 25556 1280
rect 25804 1492 25844 1532
rect 26092 4012 26132 4052
rect 25996 3340 26036 3380
rect 26188 3340 26228 3380
rect 25996 1744 26036 1784
rect 25996 1240 26036 1280
rect 25900 1156 25940 1196
rect 26572 6448 26612 6488
rect 26764 6364 26804 6404
rect 26572 6196 26612 6236
rect 26572 5860 26612 5900
rect 26476 4768 26516 4808
rect 26668 4852 26708 4892
rect 27628 8716 27668 8756
rect 27436 8380 27476 8420
rect 26956 7204 26996 7244
rect 27148 6616 27188 6656
rect 26956 6364 26996 6404
rect 27052 6280 27092 6320
rect 26956 5860 26996 5900
rect 27340 6868 27380 6908
rect 28108 9304 28148 9344
rect 27916 8800 27956 8840
rect 27820 8716 27860 8756
rect 28684 9136 28724 9176
rect 28300 8884 28340 8924
rect 28204 8716 28244 8756
rect 28588 8716 28628 8756
rect 28396 8632 28436 8672
rect 28684 8632 28724 8672
rect 28108 8548 28148 8588
rect 28588 8296 28628 8336
rect 28012 8212 28052 8252
rect 28204 8128 28244 8168
rect 27628 7876 27668 7916
rect 27820 7708 27860 7748
rect 28012 7876 28052 7916
rect 27916 6784 27956 6824
rect 27532 6364 27572 6404
rect 27436 6280 27476 6320
rect 27916 6448 27956 6488
rect 27724 6028 27764 6068
rect 27724 5692 27764 5732
rect 27244 5440 27284 5480
rect 27148 5104 27188 5144
rect 26956 4852 26996 4892
rect 26572 3592 26612 3632
rect 26668 3508 26708 3548
rect 26860 4348 26900 4388
rect 26860 4180 26900 4220
rect 26380 3340 26420 3380
rect 26380 1828 26420 1868
rect 26380 1660 26420 1700
rect 26284 988 26324 1028
rect 26572 1156 26612 1196
rect 26956 3172 26996 3212
rect 26860 1492 26900 1532
rect 27244 4432 27284 4472
rect 27244 3928 27284 3968
rect 27628 5608 27668 5648
rect 27628 4852 27668 4892
rect 27436 4180 27476 4220
rect 27628 4180 27668 4220
rect 27820 5272 27860 5312
rect 28396 7876 28436 7916
rect 28684 8212 28724 8252
rect 28972 8044 29012 8084
rect 28876 7960 28916 8000
rect 28204 7540 28244 7580
rect 28396 6784 28436 6824
rect 28108 5860 28148 5900
rect 28108 5272 28148 5312
rect 27820 4852 27860 4892
rect 27820 4600 27860 4640
rect 28012 4852 28052 4892
rect 27916 4432 27956 4472
rect 28108 4684 28148 4724
rect 28204 4516 28244 4556
rect 28204 4264 28244 4304
rect 28012 4180 28052 4220
rect 27724 4096 27764 4136
rect 28012 4012 28052 4052
rect 28780 7876 28820 7916
rect 28972 7876 29012 7916
rect 28588 7708 28628 7748
rect 28492 6364 28532 6404
rect 28492 5692 28532 5732
rect 28492 5440 28532 5480
rect 28396 5272 28436 5312
rect 28684 6364 28724 6404
rect 28780 5692 28820 5732
rect 28684 5272 28724 5312
rect 28396 5020 28436 5060
rect 28396 4768 28436 4808
rect 28396 4096 28436 4136
rect 27628 3760 27668 3800
rect 27436 3424 27476 3464
rect 27628 3424 27668 3464
rect 27052 2668 27092 2708
rect 27148 1324 27188 1364
rect 27148 988 27188 1028
rect 27724 3256 27764 3296
rect 28108 3424 28148 3464
rect 27916 3172 27956 3212
rect 28588 4516 28628 4556
rect 28588 4096 28628 4136
rect 28492 3844 28532 3884
rect 28492 3676 28532 3716
rect 27532 2416 27572 2456
rect 27436 1576 27476 1616
rect 28108 1744 28148 1784
rect 28492 2668 28532 2708
rect 28396 988 28436 1028
rect 29164 6448 29204 6488
rect 28972 5692 29012 5732
rect 30604 11068 30644 11108
rect 31372 11068 31412 11108
rect 30508 10900 30548 10940
rect 29644 9472 29684 9512
rect 29356 8716 29396 8756
rect 29548 8716 29588 8756
rect 29548 7372 29588 7412
rect 30220 10396 30260 10436
rect 30412 10396 30452 10436
rect 30316 10228 30356 10268
rect 30412 10060 30452 10100
rect 30316 9892 30356 9932
rect 30988 10984 31028 11024
rect 30796 10900 30836 10940
rect 30604 10816 30644 10856
rect 31180 10900 31220 10940
rect 36172 10984 36212 11024
rect 31084 10816 31124 10856
rect 30796 10648 30836 10688
rect 30988 10648 31028 10688
rect 30796 10228 30836 10268
rect 30700 10060 30740 10100
rect 30604 9976 30644 10016
rect 30508 9556 30548 9596
rect 31180 10312 31220 10352
rect 30988 9976 31028 10016
rect 30892 9724 30932 9764
rect 31084 9556 31124 9596
rect 30892 9472 30932 9512
rect 30796 9388 30836 9428
rect 30028 8716 30068 8756
rect 30220 8716 30260 8756
rect 30028 7456 30068 7496
rect 30028 7204 30068 7244
rect 29836 7120 29876 7160
rect 29740 6784 29780 6824
rect 30028 6364 30068 6404
rect 29836 6280 29876 6320
rect 28972 5188 29012 5228
rect 28876 4852 28916 4892
rect 28780 4768 28820 4808
rect 28972 4684 29012 4724
rect 29164 4516 29204 4556
rect 28876 4348 28916 4388
rect 28780 4180 28820 4220
rect 28684 3760 28724 3800
rect 29452 5272 29492 5312
rect 29356 4684 29396 4724
rect 28684 2668 28724 2708
rect 28684 1828 28724 1868
rect 28588 1240 28628 1280
rect 28876 1492 28916 1532
rect 29261 3928 29301 3968
rect 29260 3760 29300 3800
rect 29068 2752 29108 2792
rect 29548 5104 29588 5144
rect 29452 4012 29492 4052
rect 30604 9220 30644 9260
rect 30700 9052 30740 9092
rect 30988 9220 31028 9260
rect 31084 8968 31124 9008
rect 30316 6112 30356 6152
rect 30316 5860 30356 5900
rect 30124 5692 30164 5732
rect 30604 5692 30644 5732
rect 30412 5608 30452 5648
rect 30508 5524 30548 5564
rect 30412 5440 30452 5480
rect 29068 1324 29108 1364
rect 28972 1156 29012 1196
rect 29644 3424 29684 3464
rect 29452 1744 29492 1784
rect 29452 1576 29492 1616
rect 29836 4684 29876 4724
rect 29932 4180 29972 4220
rect 30316 4684 30356 4724
rect 30220 4600 30260 4640
rect 30124 4180 30164 4220
rect 30316 4180 30356 4220
rect 30028 3340 30068 3380
rect 29932 1324 29972 1364
rect 29836 1240 29876 1280
rect 29740 904 29780 944
rect 30316 3424 30356 3464
rect 30604 5188 30644 5228
rect 30508 4852 30548 4892
rect 30796 8212 30836 8252
rect 36076 10900 36116 10940
rect 31372 10648 31412 10688
rect 31564 10564 31604 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 31948 10480 31988 10520
rect 31564 10144 31604 10184
rect 31372 9976 31412 10016
rect 31756 8632 31796 8672
rect 31276 8044 31316 8084
rect 30796 7876 30836 7916
rect 30988 7876 31028 7916
rect 31180 7876 31220 7916
rect 30892 7792 30932 7832
rect 31276 7792 31316 7832
rect 31564 7876 31604 7916
rect 31660 7792 31700 7832
rect 31372 7708 31412 7748
rect 30988 7456 31028 7496
rect 35596 10396 35636 10436
rect 36172 10480 36212 10520
rect 32044 9976 32084 10016
rect 35788 10228 35828 10268
rect 35980 10228 36020 10268
rect 36460 10648 36500 10688
rect 36652 10732 36692 10772
rect 36652 10564 36692 10604
rect 36364 10228 36404 10268
rect 35884 10060 35924 10100
rect 35692 9976 35732 10016
rect 34540 9892 34580 9932
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 35116 9640 35156 9680
rect 32236 9388 32276 9428
rect 33388 9136 33428 9176
rect 32620 8884 32660 8924
rect 32140 8380 32180 8420
rect 32140 7960 32180 8000
rect 31948 7876 31988 7916
rect 32044 7792 32084 7832
rect 32524 8548 32564 8588
rect 32428 7960 32468 8000
rect 32332 7792 32372 7832
rect 32908 8296 32948 8336
rect 32908 8128 32948 8168
rect 32812 7876 32852 7916
rect 32716 7792 32756 7832
rect 31660 7120 31700 7160
rect 30988 6952 31028 6992
rect 31180 6952 31220 6992
rect 30892 5860 30932 5900
rect 31084 5860 31124 5900
rect 30796 5692 30836 5732
rect 30700 5104 30740 5144
rect 30700 4936 30740 4976
rect 31660 6784 31700 6824
rect 31564 6700 31604 6740
rect 31660 6616 31700 6656
rect 31660 6280 31700 6320
rect 31468 6196 31508 6236
rect 31276 5776 31316 5816
rect 31084 5440 31124 5480
rect 30892 4852 30932 4892
rect 30796 4684 30836 4724
rect 30796 4432 30836 4472
rect 30700 4348 30740 4388
rect 30508 3844 30548 3884
rect 30508 3676 30548 3716
rect 30892 4180 30932 4220
rect 30892 4012 30932 4052
rect 31660 5692 31700 5732
rect 31660 5440 31700 5480
rect 31948 7204 31988 7244
rect 32140 7204 32180 7244
rect 32332 7204 32372 7244
rect 32332 7036 32372 7076
rect 32140 6952 32180 6992
rect 32044 6868 32084 6908
rect 31852 6616 31892 6656
rect 32236 6784 32276 6824
rect 32044 6364 32084 6404
rect 32236 6532 32276 6572
rect 31852 6028 31892 6068
rect 31852 5776 31892 5816
rect 32044 5692 32084 5732
rect 31948 5440 31988 5480
rect 31852 5356 31892 5396
rect 31660 5020 31700 5060
rect 31564 4852 31604 4892
rect 31564 4684 31604 4724
rect 31084 4432 31124 4472
rect 31084 4264 31124 4304
rect 31468 4264 31508 4304
rect 31276 4180 31316 4220
rect 30220 3172 30260 3212
rect 30316 3088 30356 3128
rect 30220 1744 30260 1784
rect 30220 1240 30260 1280
rect 30604 2836 30644 2876
rect 31276 3928 31316 3968
rect 30892 2248 30932 2288
rect 31660 4180 31700 4220
rect 31276 3088 31316 3128
rect 31276 2752 31316 2792
rect 31180 2668 31220 2708
rect 30988 1576 31028 1616
rect 30412 1156 30452 1196
rect 30124 1072 30164 1112
rect 30988 1072 31028 1112
rect 30796 988 30836 1028
rect 30604 904 30644 944
rect 31564 3172 31604 3212
rect 31852 4012 31892 4052
rect 32332 6280 32372 6320
rect 32332 5944 32372 5984
rect 33196 7876 33236 7916
rect 33100 7792 33140 7832
rect 33292 7624 33332 7664
rect 32812 7540 32852 7580
rect 33292 7372 33332 7412
rect 33196 7120 33236 7160
rect 32620 6364 32660 6404
rect 32716 6112 32756 6152
rect 32428 5692 32468 5732
rect 32524 5608 32564 5648
rect 32332 5524 32372 5564
rect 32236 5440 32276 5480
rect 32428 5440 32468 5480
rect 32620 5524 32660 5564
rect 32812 5692 32852 5732
rect 32812 5272 32852 5312
rect 32236 4264 32276 4304
rect 32044 4096 32084 4136
rect 31948 3592 31988 3632
rect 31948 3424 31988 3464
rect 31756 3340 31796 3380
rect 32140 2920 32180 2960
rect 32044 2836 32084 2876
rect 31756 2752 31796 2792
rect 31660 1996 31700 2036
rect 31756 1324 31796 1364
rect 31564 1240 31604 1280
rect 31372 1156 31412 1196
rect 32332 1996 32372 2036
rect 32236 736 32276 776
rect 32716 4768 32756 4808
rect 33292 7036 33332 7076
rect 33004 6448 33044 6488
rect 33196 6448 33236 6488
rect 33100 6364 33140 6404
rect 33484 8968 33524 9008
rect 33388 5944 33428 5984
rect 33100 5860 33140 5900
rect 33292 5440 33332 5480
rect 33676 8632 33716 8672
rect 33580 7876 33620 7916
rect 34156 8716 34196 8756
rect 34348 8716 34388 8756
rect 34060 8464 34100 8504
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33772 8044 33812 8084
rect 34540 8548 34580 8588
rect 34444 8296 34484 8336
rect 34924 9304 34964 9344
rect 34828 9220 34868 9260
rect 34828 8884 34868 8924
rect 34732 8716 34772 8756
rect 35116 9220 35156 9260
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35692 8800 35732 8840
rect 35116 8716 35156 8756
rect 35500 8716 35540 8756
rect 35308 8632 35348 8672
rect 35692 8632 35732 8672
rect 35020 8380 35060 8420
rect 34828 8212 34868 8252
rect 35020 8212 35060 8252
rect 34636 8128 34676 8168
rect 35308 8128 35348 8168
rect 34924 7960 34964 8000
rect 34444 7876 34484 7916
rect 33868 7792 33908 7832
rect 33676 7540 33716 7580
rect 33868 7372 33908 7412
rect 33868 7204 33908 7244
rect 34060 7204 34100 7244
rect 34348 7204 34388 7244
rect 34252 7120 34292 7160
rect 33964 6952 34004 6992
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33676 6700 33716 6740
rect 34060 6616 34100 6656
rect 33868 6364 33908 6404
rect 34828 7876 34868 7916
rect 35020 7792 35060 7832
rect 34636 7708 34676 7748
rect 35596 8464 35636 8504
rect 36556 10144 36596 10184
rect 49900 11404 49940 11444
rect 49048 11320 49088 11360
rect 49130 11320 49170 11360
rect 49212 11320 49252 11360
rect 49294 11320 49334 11360
rect 49376 11320 49416 11360
rect 37036 10816 37076 10856
rect 37420 10816 37460 10856
rect 37996 10816 38036 10856
rect 36940 10312 36980 10352
rect 36748 10228 36788 10268
rect 36940 10144 36980 10184
rect 36652 9808 36692 9848
rect 36844 9724 36884 9764
rect 36364 9556 36404 9596
rect 36460 9472 36500 9512
rect 36268 9388 36308 9428
rect 36652 9388 36692 9428
rect 36844 9304 36884 9344
rect 36940 9220 36980 9260
rect 36844 8968 36884 9008
rect 36748 8212 36788 8252
rect 35020 7624 35060 7664
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 34636 7372 34676 7412
rect 34636 7204 34676 7244
rect 34540 7036 34580 7076
rect 34444 6784 34484 6824
rect 34732 7120 34772 7160
rect 34636 6532 34676 6572
rect 34348 6364 34388 6404
rect 34156 6280 34196 6320
rect 33772 6196 33812 6236
rect 33772 5944 33812 5984
rect 34156 5860 34196 5900
rect 34540 6196 34580 6236
rect 34540 5776 34580 5816
rect 34348 5692 34388 5732
rect 34828 6868 34868 6908
rect 35500 6532 35540 6572
rect 35020 6364 35060 6404
rect 34732 6028 34772 6068
rect 34732 5692 34772 5732
rect 33004 4936 33044 4976
rect 33484 5272 33524 5312
rect 33388 4936 33428 4976
rect 32716 4264 32756 4304
rect 32716 4096 32756 4136
rect 32524 2668 32564 2708
rect 32428 1240 32468 1280
rect 33004 4096 33044 4136
rect 32812 1744 32852 1784
rect 32716 1576 32756 1616
rect 33100 3592 33140 3632
rect 33100 3340 33140 3380
rect 32908 904 32948 944
rect 32908 736 32948 776
rect 33196 1996 33236 2036
rect 33964 5440 34004 5480
rect 34348 5440 34388 5480
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 34156 5104 34196 5144
rect 33580 4936 33620 4976
rect 33772 4936 33812 4976
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 36172 7876 36212 7916
rect 36748 7876 36788 7916
rect 36460 7120 36500 7160
rect 36172 6952 36212 6992
rect 35596 5860 35636 5900
rect 34924 5608 34964 5648
rect 34924 5272 34964 5312
rect 34828 5104 34868 5144
rect 34252 4852 34292 4892
rect 34540 4852 34580 4892
rect 34732 4852 34772 4892
rect 33580 4684 33620 4724
rect 33772 4684 33812 4724
rect 33580 3928 33620 3968
rect 33868 4516 33908 4556
rect 33868 4180 33908 4220
rect 34060 4600 34100 4640
rect 34348 4516 34388 4556
rect 34252 4348 34292 4388
rect 34060 4096 34100 4136
rect 34252 4096 34292 4136
rect 34444 4180 34484 4220
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 33580 3424 33620 3464
rect 33868 2836 33908 2876
rect 33292 1156 33332 1196
rect 33484 1240 33524 1280
rect 33388 904 33428 944
rect 33772 988 33812 1028
rect 34252 3592 34292 3632
rect 34060 2752 34100 2792
rect 33964 2332 34004 2372
rect 34636 4432 34676 4472
rect 34732 4180 34772 4220
rect 34636 4012 34676 4052
rect 35404 5692 35444 5732
rect 35878 6364 35884 6404
rect 35884 6364 35918 6404
rect 35980 6364 36020 6404
rect 36844 7624 36884 7664
rect 36748 7540 36788 7580
rect 36652 6952 36692 6992
rect 36844 6784 36884 6824
rect 36364 6364 36404 6404
rect 36844 6364 36884 6404
rect 35308 5356 35348 5396
rect 35116 5104 35156 5144
rect 35404 5188 35444 5228
rect 35116 4852 35156 4892
rect 35308 4768 35348 4808
rect 35020 4684 35060 4724
rect 35500 4684 35540 4724
rect 35884 4852 35924 4892
rect 36268 5692 36308 5732
rect 36556 5692 36596 5732
rect 36460 5608 36500 5648
rect 36268 4852 36308 4892
rect 35692 4684 35732 4724
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35596 4516 35636 4556
rect 35020 4348 35060 4388
rect 35020 4180 35060 4220
rect 35500 4180 35540 4220
rect 35788 4348 35828 4388
rect 35116 4096 35156 4136
rect 35020 3676 35060 3716
rect 34924 3508 34964 3548
rect 35596 3844 35636 3884
rect 35308 3760 35348 3800
rect 35116 3592 35156 3632
rect 34636 2920 34676 2960
rect 34444 2332 34484 2372
rect 34348 2248 34388 2288
rect 34252 1744 34292 1784
rect 34156 1072 34196 1112
rect 34540 1576 34580 1616
rect 34828 1996 34868 2036
rect 34732 1240 34772 1280
rect 35500 3172 35540 3212
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35212 2668 35252 2708
rect 35020 2248 35060 2288
rect 34924 1324 34964 1364
rect 35404 1156 35444 1196
rect 35692 3424 35732 3464
rect 36172 4684 36212 4724
rect 36076 4264 36116 4304
rect 36172 4012 36212 4052
rect 36460 4936 36500 4976
rect 37036 8716 37076 8756
rect 37324 10480 37364 10520
rect 37324 10228 37364 10268
rect 38092 10564 38132 10604
rect 37996 10312 38036 10352
rect 37612 10228 37652 10268
rect 37804 10228 37844 10268
rect 38764 10480 38804 10520
rect 38380 10396 38420 10436
rect 38188 10228 38228 10268
rect 38764 10312 38804 10352
rect 38572 10228 38612 10268
rect 37900 10060 37940 10100
rect 38092 10060 38132 10100
rect 38956 10228 38996 10268
rect 39148 10144 39188 10184
rect 38380 10060 38420 10100
rect 37900 9640 37940 9680
rect 37516 9472 37556 9512
rect 37324 9388 37364 9428
rect 37900 9388 37940 9428
rect 38188 9388 38228 9428
rect 37804 9220 37844 9260
rect 37996 9220 38036 9260
rect 37324 8716 37364 8756
rect 37324 8464 37364 8504
rect 37228 7456 37268 7496
rect 37708 8044 37748 8084
rect 37420 7876 37460 7916
rect 37420 7540 37460 7580
rect 37612 7540 37652 7580
rect 37516 7456 37556 7496
rect 37324 7204 37364 7244
rect 37324 6448 37364 6488
rect 37324 6196 37364 6236
rect 37228 6112 37268 6152
rect 37036 5776 37076 5816
rect 36652 4936 36692 4976
rect 36556 4852 36596 4892
rect 36748 4516 36788 4556
rect 35884 3760 35924 3800
rect 36076 3424 36116 3464
rect 35788 3256 35828 3296
rect 35788 2920 35828 2960
rect 35884 1660 35924 1700
rect 35788 1240 35828 1280
rect 36172 904 36212 944
rect 35980 820 36020 860
rect 36844 3760 36884 3800
rect 37324 5440 37364 5480
rect 37036 4852 37076 4892
rect 37228 4852 37268 4892
rect 36940 3256 36980 3296
rect 36940 3088 36980 3128
rect 36748 1996 36788 2036
rect 36748 1576 36788 1616
rect 36652 1408 36692 1448
rect 36364 1240 36404 1280
rect 36556 1072 36596 1112
rect 36364 988 36404 1028
rect 36268 148 36308 188
rect 37228 3256 37268 3296
rect 37228 2416 37268 2456
rect 37132 2080 37172 2120
rect 37132 1240 37172 1280
rect 37036 1156 37076 1196
rect 37516 7204 37556 7244
rect 37516 6952 37556 6992
rect 37708 7288 37748 7328
rect 37708 7120 37748 7160
rect 38092 9136 38132 9176
rect 38476 9304 38516 9344
rect 38380 9220 38420 9260
rect 38572 9052 38612 9092
rect 38380 8968 38420 9008
rect 37996 8884 38036 8924
rect 37900 7204 37940 7244
rect 37900 6532 37940 6572
rect 37804 6448 37844 6488
rect 37516 5776 37556 5816
rect 37708 5692 37748 5732
rect 37516 5524 37556 5564
rect 37708 5440 37748 5480
rect 37516 4936 37556 4976
rect 37612 4768 37652 4808
rect 37612 4264 37652 4304
rect 37420 3340 37460 3380
rect 37516 3172 37556 3212
rect 37516 3004 37556 3044
rect 37900 6280 37940 6320
rect 37900 6028 37940 6068
rect 37900 5440 37940 5480
rect 38188 8212 38228 8252
rect 38284 8044 38324 8084
rect 38284 7204 38324 7244
rect 38092 6700 38132 6740
rect 38092 6364 38132 6404
rect 38956 9388 38996 9428
rect 38860 9052 38900 9092
rect 38764 8968 38804 9008
rect 38668 8296 38708 8336
rect 39052 8128 39092 8168
rect 40780 10900 40820 10940
rect 40588 10732 40628 10772
rect 40684 10144 40724 10184
rect 40204 9892 40244 9932
rect 40012 9808 40052 9848
rect 39340 9388 39380 9428
rect 39916 8548 39956 8588
rect 39628 8380 39668 8420
rect 39244 7456 39284 7496
rect 38668 6784 38708 6824
rect 38668 6616 38708 6656
rect 38764 6448 38804 6488
rect 39340 7036 39380 7076
rect 39148 6364 39188 6404
rect 39532 7288 39572 7328
rect 39436 6868 39476 6908
rect 38284 6280 38324 6320
rect 38860 6280 38900 6320
rect 38188 6028 38228 6068
rect 38092 5608 38132 5648
rect 38092 5272 38132 5312
rect 38956 6028 38996 6068
rect 38572 5692 38612 5732
rect 38764 5692 38804 5732
rect 38572 5440 38612 5480
rect 37804 4348 37844 4388
rect 37804 4180 37844 4220
rect 37804 3928 37844 3968
rect 37996 4516 38036 4556
rect 37996 3676 38036 3716
rect 37708 1996 37748 2036
rect 37516 1660 37556 1700
rect 37420 1576 37460 1616
rect 38188 4180 38228 4220
rect 38188 3928 38228 3968
rect 38092 2332 38132 2372
rect 38380 4684 38420 4724
rect 38668 4768 38708 4808
rect 38572 4180 38612 4220
rect 38572 4012 38612 4052
rect 38764 4348 38804 4388
rect 39148 5860 39188 5900
rect 39148 5692 39188 5732
rect 39052 5608 39092 5648
rect 39340 5608 39380 5648
rect 38956 4516 38996 4556
rect 39340 4852 39380 4892
rect 38956 4180 38996 4220
rect 38764 4096 38804 4136
rect 38668 3928 38708 3968
rect 38764 3760 38804 3800
rect 38380 3424 38420 3464
rect 38284 3004 38324 3044
rect 39052 3592 39092 3632
rect 38956 3424 38996 3464
rect 38860 3340 38900 3380
rect 38476 2920 38516 2960
rect 38476 2332 38516 2372
rect 38284 2080 38324 2120
rect 38188 1744 38228 1784
rect 37996 1660 38036 1700
rect 38092 64 38132 104
rect 38572 1492 38612 1532
rect 38668 1408 38708 1448
rect 39148 3088 39188 3128
rect 39052 2836 39092 2876
rect 39340 4180 39380 4220
rect 39340 3928 39380 3968
rect 39244 2752 39284 2792
rect 39244 1576 39284 1616
rect 39052 1156 39092 1196
rect 38956 1072 38996 1112
rect 39340 568 39380 608
rect 39724 8044 39764 8084
rect 39724 7708 39764 7748
rect 39724 5356 39764 5396
rect 39820 5188 39860 5228
rect 39628 4852 39668 4892
rect 39820 4432 39860 4472
rect 39532 3592 39572 3632
rect 39532 3256 39572 3296
rect 39532 1660 39572 1700
rect 39724 1576 39764 1616
rect 39628 1240 39668 1280
rect 40300 9304 40340 9344
rect 40588 8716 40628 8756
rect 40396 7960 40436 8000
rect 40108 7204 40148 7244
rect 40204 6616 40244 6656
rect 41260 10648 41300 10688
rect 48652 10648 48692 10688
rect 40876 8464 40916 8504
rect 40108 4600 40148 4640
rect 40300 4096 40340 4136
rect 39916 3172 39956 3212
rect 40012 1744 40052 1784
rect 40300 3760 40340 3800
rect 40108 1660 40148 1700
rect 40204 1492 40244 1532
rect 40300 1156 40340 1196
rect 40588 4096 40628 4136
rect 41164 7876 41204 7916
rect 41548 10396 41588 10436
rect 49804 10396 49844 10436
rect 49420 10312 49460 10352
rect 42796 10228 42836 10268
rect 48652 10228 48692 10268
rect 41836 10060 41876 10100
rect 42316 9724 42356 9764
rect 46252 9724 46292 9764
rect 43660 9640 43700 9680
rect 43084 9556 43124 9596
rect 42700 9136 42740 9176
rect 41548 8968 41588 9008
rect 42508 8632 42548 8672
rect 42412 8380 42452 8420
rect 41356 7708 41396 7748
rect 42124 7876 42164 7916
rect 42028 7624 42068 7664
rect 41932 7120 41972 7160
rect 41740 6784 41780 6824
rect 41644 6364 41684 6404
rect 41260 5944 41300 5984
rect 40780 5692 40820 5732
rect 40876 5188 40916 5228
rect 40588 3508 40628 3548
rect 40492 3340 40532 3380
rect 40684 3256 40724 3296
rect 40972 5020 41012 5060
rect 41740 5440 41780 5480
rect 41548 5020 41588 5060
rect 40876 4096 40916 4136
rect 40876 3508 40916 3548
rect 40780 2332 40820 2372
rect 40876 1408 40916 1448
rect 40780 1240 40820 1280
rect 40588 1072 40628 1112
rect 40492 736 40532 776
rect 41068 4096 41108 4136
rect 41068 3760 41108 3800
rect 41836 4684 41876 4724
rect 41356 4348 41396 4388
rect 41452 4096 41492 4136
rect 41260 3760 41300 3800
rect 41356 3508 41396 3548
rect 41164 2500 41204 2540
rect 41164 2332 41204 2372
rect 41548 3088 41588 3128
rect 41548 2668 41588 2708
rect 41356 1996 41396 2036
rect 41548 1156 41588 1196
rect 41356 568 41396 608
rect 41260 316 41300 356
rect 41836 3424 41876 3464
rect 41740 2668 41780 2708
rect 42604 5356 42644 5396
rect 42988 7372 43028 7412
rect 42892 7036 42932 7076
rect 43276 9304 43316 9344
rect 43372 8716 43412 8756
rect 43756 9052 43796 9092
rect 43372 7876 43412 7916
rect 43468 7204 43508 7244
rect 43468 6532 43508 6572
rect 43276 5608 43316 5648
rect 43660 5608 43700 5648
rect 42700 5104 42740 5144
rect 42508 5020 42548 5060
rect 42988 5020 43028 5060
rect 42220 4768 42260 4808
rect 42220 3844 42260 3884
rect 42028 3508 42068 3548
rect 42124 3340 42164 3380
rect 41740 2500 41780 2540
rect 41932 2500 41972 2540
rect 41644 904 41684 944
rect 41932 1576 41972 1616
rect 42028 988 42068 1028
rect 42220 2668 42260 2708
rect 42604 4096 42644 4136
rect 42988 4096 43028 4136
rect 42796 4012 42836 4052
rect 42988 3844 43028 3884
rect 42604 3592 42644 3632
rect 42892 3592 42932 3632
rect 42508 2668 42548 2708
rect 42700 1996 42740 2036
rect 42508 1660 42548 1700
rect 42412 1576 42452 1616
rect 42316 232 42356 272
rect 43372 4096 43412 4136
rect 43180 3928 43220 3968
rect 43276 3760 43316 3800
rect 43180 3004 43220 3044
rect 42892 2920 42932 2960
rect 43084 2920 43124 2960
rect 42892 2500 42932 2540
rect 42796 1240 42836 1280
rect 43084 736 43124 776
rect 43564 3760 43604 3800
rect 43468 3676 43508 3716
rect 43372 3424 43412 3464
rect 43468 2920 43508 2960
rect 43564 2836 43604 2876
rect 44140 8800 44180 8840
rect 44620 8380 44660 8420
rect 44140 8212 44180 8252
rect 44620 8212 44660 8252
rect 44044 7876 44084 7916
rect 43948 7204 43988 7244
rect 44236 7792 44276 7832
rect 44332 7624 44372 7664
rect 44908 8800 44948 8840
rect 48460 9556 48500 9596
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 48940 9556 48980 9596
rect 47596 9472 47636 9512
rect 47020 9220 47060 9260
rect 44908 8548 44948 8588
rect 44620 7540 44660 7580
rect 44428 7204 44468 7244
rect 44524 6952 44564 6992
rect 44140 5860 44180 5900
rect 45004 7876 45044 7916
rect 44908 7204 44948 7244
rect 44428 6448 44468 6488
rect 44332 6028 44372 6068
rect 44332 5776 44372 5816
rect 44044 5440 44084 5480
rect 44140 5188 44180 5228
rect 44236 5020 44276 5060
rect 44332 4600 44372 4640
rect 43948 3340 43988 3380
rect 44332 3508 44372 3548
rect 45196 8548 45236 8588
rect 45388 7960 45428 8000
rect 45580 7960 45620 8000
rect 46252 8716 46292 8756
rect 46540 8548 46580 8588
rect 46924 8464 46964 8504
rect 45580 7708 45620 7748
rect 45868 7876 45908 7916
rect 46156 7876 46196 7916
rect 45868 7708 45908 7748
rect 45292 7540 45332 7580
rect 45772 7540 45812 7580
rect 45196 7204 45236 7244
rect 44812 6448 44852 6488
rect 45100 6448 45140 6488
rect 44716 6364 44756 6404
rect 44716 5776 44756 5816
rect 45100 6112 45140 6152
rect 45196 5776 45236 5816
rect 44620 5440 44660 5480
rect 44524 4600 44564 4640
rect 44620 4180 44660 4220
rect 44716 3424 44756 3464
rect 44236 3088 44276 3128
rect 43948 2920 43988 2960
rect 43852 2584 43892 2624
rect 43660 1408 43700 1448
rect 44332 2752 44372 2792
rect 44236 316 44276 356
rect 44620 3340 44660 3380
rect 44716 2584 44756 2624
rect 45676 6364 45716 6404
rect 45964 7372 46004 7412
rect 45676 5944 45716 5984
rect 45292 5608 45332 5648
rect 45388 5440 45428 5480
rect 45964 5944 46004 5984
rect 46060 5776 46100 5816
rect 45868 5440 45908 5480
rect 45676 5272 45716 5312
rect 45580 5104 45620 5144
rect 45580 4684 45620 4724
rect 45484 4348 45524 4388
rect 45580 4180 45620 4220
rect 45388 4012 45428 4052
rect 45100 3340 45140 3380
rect 44908 2416 44948 2456
rect 45292 2668 45332 2708
rect 45100 1156 45140 1196
rect 45196 988 45236 1028
rect 44812 904 44852 944
rect 45004 232 45044 272
rect 45484 2500 45524 2540
rect 46540 7876 46580 7916
rect 46924 7876 46964 7916
rect 46540 7708 46580 7748
rect 46444 7540 46484 7580
rect 46636 7372 46676 7412
rect 46348 7120 46388 7160
rect 46636 7120 46676 7160
rect 46636 6952 46676 6992
rect 47116 8632 47156 8672
rect 47308 7960 47348 8000
rect 47212 7708 47252 7748
rect 47116 7540 47156 7580
rect 46732 6784 46772 6824
rect 46348 6112 46388 6152
rect 46828 5944 46868 5984
rect 46156 4936 46196 4976
rect 45868 4684 45908 4724
rect 45964 4348 46004 4388
rect 45772 3928 45812 3968
rect 45580 2416 45620 2456
rect 45580 1576 45620 1616
rect 46636 5188 46676 5228
rect 46636 4936 46676 4976
rect 46828 4936 46868 4976
rect 46540 4768 46580 4808
rect 46444 4096 46484 4136
rect 46060 4012 46100 4052
rect 46156 3760 46196 3800
rect 45868 2668 45908 2708
rect 45964 1240 46004 1280
rect 46252 3340 46292 3380
rect 46636 4432 46676 4472
rect 46828 3760 46868 3800
rect 46732 3592 46772 3632
rect 47020 5944 47060 5984
rect 47212 6784 47252 6824
rect 47500 8128 47540 8168
rect 47404 6448 47444 6488
rect 47020 4768 47060 4808
rect 47116 4684 47156 4724
rect 47116 4180 47156 4220
rect 46636 3256 46676 3296
rect 46348 3004 46388 3044
rect 46636 3004 46676 3044
rect 46540 2836 46580 2876
rect 46636 2584 46676 2624
rect 46924 2920 46964 2960
rect 47116 2752 47156 2792
rect 47308 4936 47348 4976
rect 47308 4180 47348 4220
rect 48172 9136 48212 9176
rect 48076 8548 48116 8588
rect 49804 9472 49844 9512
rect 48844 8968 48884 9008
rect 48460 8800 48500 8840
rect 48364 8716 48404 8756
rect 48268 8632 48308 8672
rect 48748 8716 48788 8756
rect 48268 8128 48308 8168
rect 48172 7204 48212 7244
rect 48364 7204 48404 7244
rect 47980 6868 48020 6908
rect 47884 6532 47924 6572
rect 47692 6448 47732 6488
rect 48076 6364 48116 6404
rect 48748 7792 48788 7832
rect 49612 9220 49652 9260
rect 49324 8968 49364 9008
rect 49612 8968 49652 9008
rect 49420 8800 49460 8840
rect 48940 8632 48980 8672
rect 53164 11908 53204 11948
rect 59692 11908 59732 11948
rect 52108 10816 52148 10856
rect 50284 10732 50324 10772
rect 51244 10732 51284 10772
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 50284 10396 50324 10436
rect 51148 10396 51188 10436
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 49708 8800 49748 8840
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 49516 8212 49556 8252
rect 49420 8128 49460 8168
rect 49132 7708 49172 7748
rect 49996 8716 50036 8756
rect 50764 8212 50804 8252
rect 49612 7876 49652 7916
rect 50092 7876 50132 7916
rect 49516 7708 49556 7748
rect 49228 7540 49268 7580
rect 48652 7120 48692 7160
rect 48556 6868 48596 6908
rect 48460 6784 48500 6824
rect 49324 7204 49364 7244
rect 49996 7792 50036 7832
rect 49900 7540 49940 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 51148 8212 51188 8252
rect 50764 7456 50804 7496
rect 50956 7456 50996 7496
rect 50572 7372 50612 7412
rect 49036 6952 49076 6992
rect 49324 6952 49364 6992
rect 48748 6784 48788 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 47884 5944 47924 5984
rect 48268 5860 48308 5900
rect 47884 5608 47924 5648
rect 48652 5692 48692 5732
rect 47500 4768 47540 4808
rect 47596 4264 47636 4304
rect 47500 3760 47540 3800
rect 47212 1072 47252 1112
rect 47404 3004 47444 3044
rect 47500 2920 47540 2960
rect 47788 4936 47828 4976
rect 47788 4684 47828 4724
rect 47980 4516 48020 4556
rect 48364 4936 48404 4976
rect 48748 4936 48788 4976
rect 48460 4684 48500 4724
rect 48172 3508 48212 3548
rect 47980 3424 48020 3464
rect 48364 2752 48404 2792
rect 48268 2584 48308 2624
rect 48172 1576 48212 1616
rect 47692 1240 47732 1280
rect 48076 1240 48116 1280
rect 47884 1156 47924 1196
rect 47692 1072 47732 1112
rect 48556 3676 48596 3716
rect 48748 3088 48788 3128
rect 48652 3004 48692 3044
rect 48748 2668 48788 2708
rect 48556 1492 48596 1532
rect 49324 6364 49364 6404
rect 50380 6364 50420 6404
rect 50188 6280 50228 6320
rect 49612 5692 49652 5732
rect 50764 7204 50804 7244
rect 50668 6700 50708 6740
rect 50860 6448 50900 6488
rect 50764 6364 50804 6404
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 52492 10480 52532 10520
rect 53068 10480 53108 10520
rect 52108 9556 52148 9596
rect 52300 9556 52340 9596
rect 51436 9388 51476 9428
rect 51820 9388 51860 9428
rect 52012 9388 52052 9428
rect 51436 9220 51476 9260
rect 51340 8212 51380 8252
rect 51340 7960 51380 8000
rect 51244 7372 51284 7412
rect 52012 9220 52052 9260
rect 51532 7372 51572 7412
rect 51244 7204 51284 7244
rect 51436 7204 51476 7244
rect 51436 6784 51476 6824
rect 51244 6532 51284 6572
rect 51436 6448 51476 6488
rect 51628 7204 51668 7244
rect 51532 6364 51572 6404
rect 51916 7372 51956 7412
rect 51916 7204 51956 7244
rect 51724 7120 51764 7160
rect 51820 7036 51860 7076
rect 53068 9556 53108 9596
rect 52396 9304 52436 9344
rect 52588 9220 52628 9260
rect 52876 8716 52916 8756
rect 52396 8632 52436 8672
rect 52684 8632 52724 8672
rect 52204 7372 52244 7412
rect 52108 7120 52148 7160
rect 52108 6952 52148 6992
rect 52300 7204 52340 7244
rect 52300 6532 52340 6572
rect 52012 6448 52052 6488
rect 51916 6364 51956 6404
rect 51052 6280 51092 6320
rect 52684 8212 52724 8252
rect 52588 6868 52628 6908
rect 52876 7540 52916 7580
rect 52780 7120 52820 7160
rect 52588 6448 52628 6488
rect 50956 5776 50996 5816
rect 51532 6196 51572 6236
rect 51436 5692 51476 5732
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 49036 5020 49076 5060
rect 48940 4936 48980 4976
rect 50476 4936 50516 4976
rect 50956 4936 50996 4976
rect 49516 4852 49556 4892
rect 49708 4852 49748 4892
rect 49900 4852 49940 4892
rect 49996 4768 50036 4808
rect 49228 4684 49268 4724
rect 49036 4264 49076 4304
rect 49612 4684 49652 4724
rect 49804 4684 49844 4724
rect 49516 4217 49556 4220
rect 49516 4180 49556 4217
rect 49228 3928 49268 3968
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 49516 3760 49556 3800
rect 48940 3592 48980 3632
rect 49420 3592 49460 3632
rect 49036 3508 49076 3548
rect 48940 3172 48980 3212
rect 49132 3424 49172 3464
rect 49324 3340 49364 3380
rect 49228 3256 49268 3296
rect 49228 3004 49268 3044
rect 50572 4768 50612 4808
rect 50188 4684 50228 4724
rect 50380 4684 50420 4724
rect 50188 4516 50228 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 49996 4180 50036 4220
rect 49708 3928 49748 3968
rect 49900 3844 49940 3884
rect 49516 3340 49556 3380
rect 49612 3256 49652 3296
rect 50284 4096 50324 4136
rect 50188 4012 50228 4052
rect 50092 3760 50132 3800
rect 50860 4684 50900 4724
rect 52684 6364 52724 6404
rect 53068 7204 53108 7244
rect 52492 6280 52532 6320
rect 52588 6112 52628 6152
rect 52204 5356 52244 5396
rect 52108 5020 52148 5060
rect 51724 4852 51764 4892
rect 52396 4936 52436 4976
rect 52204 4348 52244 4388
rect 50956 4096 50996 4136
rect 52108 4180 52148 4220
rect 51244 4012 51284 4052
rect 51628 4012 51668 4052
rect 50188 3172 50228 3212
rect 49804 1576 49844 1616
rect 49996 1492 50036 1532
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 50476 2836 50516 2876
rect 50572 1996 50612 2036
rect 52204 3676 52244 3716
rect 51436 3508 51476 3548
rect 51820 3424 51860 3464
rect 50956 2836 50996 2876
rect 50860 1996 50900 2036
rect 51916 1660 51956 1700
rect 51532 1576 51572 1616
rect 51724 1240 51764 1280
rect 52876 6280 52916 6320
rect 52780 5104 52820 5144
rect 57676 10564 57716 10604
rect 56236 10312 56276 10352
rect 57580 10312 57620 10352
rect 53452 10060 53492 10100
rect 58060 10396 58100 10436
rect 57292 10060 57332 10100
rect 58156 10312 58196 10352
rect 58636 10312 58676 10352
rect 58828 10312 58868 10352
rect 58444 10060 58484 10100
rect 58636 10060 58676 10100
rect 56620 9640 56660 9680
rect 55852 9556 55892 9596
rect 54796 9388 54836 9428
rect 53452 8716 53492 8756
rect 55660 9388 55700 9428
rect 55468 9052 55508 9092
rect 54995 8800 55035 8840
rect 54316 8632 54356 8672
rect 53836 8464 53876 8504
rect 53356 6700 53396 6740
rect 53356 6448 53396 6488
rect 53260 6280 53300 6320
rect 53164 5104 53204 5144
rect 52876 4936 52916 4976
rect 53452 6112 53492 6152
rect 53260 4684 53300 4724
rect 53260 4516 53300 4556
rect 52396 4180 52436 4220
rect 52972 4264 53012 4304
rect 52684 4180 52724 4220
rect 52876 4180 52916 4220
rect 52588 4096 52628 4136
rect 52492 3676 52532 3716
rect 52492 3508 52532 3548
rect 52396 3424 52436 3464
rect 52780 3928 52820 3968
rect 52012 1576 52052 1616
rect 52876 3760 52916 3800
rect 52492 1744 52532 1784
rect 52300 1576 52340 1616
rect 53356 4180 53396 4220
rect 53356 3676 53396 3716
rect 53740 5944 53780 5984
rect 53548 4264 53588 4304
rect 53740 3928 53780 3968
rect 53644 3844 53684 3884
rect 54910 8724 54932 8756
rect 54932 8724 54950 8756
rect 54910 8716 54950 8724
rect 54700 8464 54740 8504
rect 54604 8296 54644 8336
rect 54124 6196 54164 6236
rect 53932 5944 53972 5984
rect 53932 5692 53972 5732
rect 53932 4768 53972 4808
rect 54028 4600 54068 4640
rect 54124 4096 54164 4136
rect 54028 3928 54068 3968
rect 53644 3340 53684 3380
rect 53452 3172 53492 3212
rect 53356 1660 53396 1700
rect 53068 1408 53108 1448
rect 52972 1240 53012 1280
rect 53260 1240 53300 1280
rect 53740 1576 53780 1616
rect 53836 1324 53876 1364
rect 54124 3760 54164 3800
rect 54412 7960 54452 8000
rect 54700 7960 54740 8000
rect 54316 7372 54356 7412
rect 54796 7876 54836 7916
rect 55372 7876 55412 7916
rect 54412 6280 54452 6320
rect 54316 6196 54356 6236
rect 54892 7708 54932 7748
rect 55372 7624 55412 7664
rect 56140 9388 56180 9428
rect 55948 9304 55988 9344
rect 56332 9304 56372 9344
rect 56716 9304 56756 9344
rect 56812 8800 56852 8840
rect 55948 8716 55988 8756
rect 57196 8800 57236 8840
rect 56044 8548 56084 8588
rect 56140 8464 56180 8504
rect 56140 7876 56180 7916
rect 55852 7456 55892 7496
rect 55756 7372 55796 7412
rect 55660 6784 55700 6824
rect 54796 6364 54836 6404
rect 54700 6280 54740 6320
rect 54316 5692 54356 5732
rect 54316 4516 54356 4556
rect 55180 6532 55220 6572
rect 54988 6364 55028 6404
rect 54892 6196 54932 6236
rect 54604 5944 54644 5984
rect 54508 5692 54548 5732
rect 54508 4600 54548 4640
rect 54508 4348 54548 4388
rect 54988 5692 55028 5732
rect 54892 5608 54932 5648
rect 54604 2752 54644 2792
rect 55564 6364 55604 6404
rect 56140 7372 56180 7412
rect 55468 6196 55508 6236
rect 55372 6112 55412 6152
rect 55660 6112 55700 6152
rect 55276 6028 55316 6068
rect 55852 5776 55892 5816
rect 55756 5692 55796 5732
rect 55660 5524 55700 5564
rect 55372 5272 55412 5312
rect 54796 4852 54836 4892
rect 54796 4180 54836 4220
rect 54796 4012 54836 4052
rect 54796 3592 54836 3632
rect 54796 3256 54836 3296
rect 54124 1744 54164 1784
rect 54220 1576 54260 1616
rect 54604 2332 54644 2372
rect 55180 4852 55220 4892
rect 55276 4348 55316 4388
rect 54988 4264 55028 4304
rect 55084 4180 55124 4220
rect 54988 4096 55028 4136
rect 55276 3760 55316 3800
rect 55372 3592 55412 3632
rect 55468 3340 55508 3380
rect 54988 3256 55028 3296
rect 55276 3256 55316 3296
rect 54988 1492 55028 1532
rect 55276 2836 55316 2876
rect 55372 2248 55412 2288
rect 55180 1660 55220 1700
rect 55084 1408 55124 1448
rect 56236 7288 56276 7328
rect 56236 7120 56276 7160
rect 56044 6784 56084 6824
rect 56140 6280 56180 6320
rect 56428 8548 56468 8588
rect 56716 8548 56756 8588
rect 57004 8548 57044 8588
rect 57196 8548 57236 8588
rect 56620 8044 56660 8084
rect 56908 7708 56948 7748
rect 56812 7624 56852 7664
rect 56524 7540 56564 7580
rect 56332 6196 56372 6236
rect 56140 6028 56180 6068
rect 56140 5860 56180 5900
rect 56332 5860 56372 5900
rect 56524 6784 56564 6824
rect 57196 6868 57236 6908
rect 57676 8716 57716 8756
rect 57388 8464 57428 8504
rect 57772 8380 57812 8420
rect 57772 8128 57812 8168
rect 57868 7876 57908 7916
rect 57676 7624 57716 7664
rect 57772 7540 57812 7580
rect 57868 6952 57908 6992
rect 57676 6868 57716 6908
rect 56620 6532 56660 6572
rect 56524 6364 56564 6404
rect 57100 6532 57140 6572
rect 57292 6532 57332 6572
rect 57484 6448 57524 6488
rect 57004 6364 57044 6404
rect 56716 6280 56756 6320
rect 57580 6364 57620 6404
rect 57388 6280 57428 6320
rect 57196 6196 57236 6236
rect 56620 6112 56660 6152
rect 57868 6448 57908 6488
rect 57676 6028 57716 6068
rect 56524 5860 56564 5900
rect 56812 5860 56852 5900
rect 57676 5776 57716 5816
rect 56524 5524 56564 5564
rect 55948 4852 55988 4892
rect 55756 4516 55796 4556
rect 55660 4096 55700 4136
rect 55852 3928 55892 3968
rect 55852 3172 55892 3212
rect 55756 2332 55796 2372
rect 55468 1240 55508 1280
rect 55756 736 55796 776
rect 55564 232 55604 272
rect 56908 5692 56948 5732
rect 56332 4852 56372 4892
rect 56715 4936 56755 4976
rect 56908 4936 56948 4976
rect 57100 5188 57140 5228
rect 57388 5692 57428 5732
rect 57292 5272 57332 5312
rect 57484 5020 57524 5060
rect 56620 4768 56660 4808
rect 56044 4264 56084 4304
rect 56236 4432 56276 4472
rect 56140 4012 56180 4052
rect 56044 3592 56084 3632
rect 56236 1324 56276 1364
rect 56140 988 56180 1028
rect 56524 4684 56564 4724
rect 56524 4180 56564 4220
rect 56524 4012 56564 4052
rect 57100 4684 57140 4724
rect 57292 4684 57332 4724
rect 56716 4432 56756 4472
rect 57004 4432 57044 4472
rect 57100 4180 57140 4220
rect 57676 4852 57716 4892
rect 57388 4432 57428 4472
rect 57580 4432 57620 4472
rect 56428 3928 56468 3968
rect 57388 3928 57428 3968
rect 56908 3424 56948 3464
rect 56812 3172 56852 3212
rect 56716 1744 56756 1784
rect 56620 1576 56660 1616
rect 56524 1072 56564 1112
rect 57196 3340 57236 3380
rect 57580 4012 57620 4052
rect 57964 6196 58004 6236
rect 58636 9640 58676 9680
rect 58732 9556 58772 9596
rect 58156 9388 58196 9428
rect 59020 10060 59060 10100
rect 59404 9640 59444 9680
rect 59212 9556 59252 9596
rect 57868 5524 57908 5564
rect 57868 5272 57908 5312
rect 58444 8044 58484 8084
rect 58348 7960 58388 8000
rect 58252 7876 58292 7916
rect 58348 7624 58388 7664
rect 58540 6952 58580 6992
rect 58252 6364 58292 6404
rect 58444 6364 58484 6404
rect 59116 9388 59156 9428
rect 59596 9388 59636 9428
rect 58924 8716 58964 8756
rect 58732 8128 58772 8168
rect 58828 7876 58868 7916
rect 58828 7708 58868 7748
rect 58252 5440 58292 5480
rect 58156 5272 58196 5312
rect 57964 4936 58004 4976
rect 57868 4768 57908 4808
rect 58060 4684 58100 4724
rect 57964 4180 58004 4220
rect 58060 4096 58100 4136
rect 57772 3424 57812 3464
rect 57100 3172 57140 3212
rect 57100 2752 57140 2792
rect 57292 2164 57332 2204
rect 57484 1576 57524 1616
rect 57868 2752 57908 2792
rect 57676 2668 57716 2708
rect 57580 1492 57620 1532
rect 58252 4852 58292 4892
rect 58444 4852 58484 4892
rect 58444 4684 58484 4724
rect 58444 4516 58484 4556
rect 58348 4264 58388 4304
rect 58924 6364 58964 6404
rect 59308 8464 59348 8504
rect 59212 8044 59252 8084
rect 59596 9052 59636 9092
rect 59500 8044 59540 8084
rect 59500 7624 59540 7664
rect 64168 11320 64208 11360
rect 64250 11320 64290 11360
rect 64332 11320 64372 11360
rect 64414 11320 64454 11360
rect 64496 11320 64536 11360
rect 60076 10396 60116 10436
rect 60364 10396 60404 10436
rect 60076 10060 60116 10100
rect 59884 9640 59924 9680
rect 59884 9388 59924 9428
rect 60460 9724 60500 9764
rect 60364 9388 60404 9428
rect 59884 9052 59924 9092
rect 60172 9052 60212 9092
rect 59692 8800 59732 8840
rect 60076 8716 60116 8756
rect 59404 7372 59444 7412
rect 59884 7708 59924 7748
rect 59692 7372 59732 7412
rect 59212 6784 59252 6824
rect 59308 6616 59348 6656
rect 59116 6280 59156 6320
rect 59116 5944 59156 5984
rect 58732 5104 58772 5144
rect 58540 4096 58580 4136
rect 58540 3844 58580 3884
rect 58252 3760 58292 3800
rect 58156 3592 58196 3632
rect 58156 3424 58196 3464
rect 58060 2248 58100 2288
rect 57964 1660 58004 1700
rect 57868 1408 57908 1448
rect 58156 2164 58196 2204
rect 58444 2164 58484 2204
rect 58348 232 58388 272
rect 58828 4348 58868 4388
rect 58828 4180 58868 4220
rect 58732 3760 58772 3800
rect 59788 7204 59828 7244
rect 59788 6952 59828 6992
rect 59596 6112 59636 6152
rect 60364 9052 60404 9092
rect 60844 9556 60884 9596
rect 60844 9388 60884 9428
rect 60460 8800 60500 8840
rect 60556 8380 60596 8420
rect 60652 7540 60692 7580
rect 60844 8716 60884 8756
rect 60748 7456 60788 7496
rect 60364 7372 60404 7412
rect 59980 7204 60020 7244
rect 59980 6952 60020 6992
rect 59212 4936 59252 4976
rect 59020 4852 59060 4892
rect 58636 1240 58676 1280
rect 58540 988 58580 1028
rect 58924 3088 58964 3128
rect 58828 2668 58868 2708
rect 59116 4684 59156 4724
rect 58828 2500 58868 2540
rect 58732 736 58772 776
rect 59020 2332 59060 2372
rect 58924 1072 58964 1112
rect 59212 3508 59252 3548
rect 59500 5272 59540 5312
rect 59404 4936 59444 4976
rect 59500 4264 59540 4304
rect 59404 4180 59444 4220
rect 59500 3172 59540 3212
rect 59788 5440 59828 5480
rect 59692 4936 59732 4976
rect 59692 3592 59732 3632
rect 59692 3172 59732 3212
rect 59500 2584 59540 2624
rect 59884 4180 59924 4220
rect 60076 6364 60116 6404
rect 60076 5440 60116 5480
rect 60556 7372 60596 7412
rect 60268 7204 60308 7244
rect 60369 7204 60404 7244
rect 60404 7204 60409 7244
rect 60268 6616 60308 6656
rect 60652 7204 60692 7244
rect 60556 6952 60596 6992
rect 60460 6364 60500 6404
rect 60364 6280 60404 6320
rect 60556 6280 60596 6320
rect 60364 6112 60404 6152
rect 60268 5524 60308 5564
rect 60172 5020 60212 5060
rect 61036 6952 61076 6992
rect 61036 6616 61076 6656
rect 60748 6532 60788 6572
rect 60652 5608 60692 5648
rect 60076 4852 60116 4892
rect 60172 4684 60212 4724
rect 61324 10900 61364 10940
rect 79288 11320 79328 11360
rect 79370 11320 79410 11360
rect 79452 11320 79492 11360
rect 79534 11320 79574 11360
rect 79616 11320 79656 11360
rect 93772 11908 93812 11948
rect 94408 11320 94448 11360
rect 94490 11320 94530 11360
rect 94572 11320 94612 11360
rect 94654 11320 94694 11360
rect 94736 11320 94776 11360
rect 61228 8548 61268 8588
rect 61228 8380 61268 8420
rect 68428 10648 68468 10688
rect 65408 10564 65448 10604
rect 65490 10564 65530 10604
rect 65572 10564 65612 10604
rect 65654 10564 65694 10604
rect 65736 10564 65776 10604
rect 69772 10396 69812 10436
rect 71308 10396 71348 10436
rect 69580 10228 69620 10268
rect 69100 10060 69140 10100
rect 64168 9808 64208 9848
rect 64250 9808 64290 9848
rect 64332 9808 64372 9848
rect 64414 9808 64454 9848
rect 64496 9808 64536 9848
rect 67948 9556 67988 9596
rect 66892 9472 66932 9512
rect 65164 9388 65204 9428
rect 63724 9220 63764 9260
rect 62092 8968 62132 9008
rect 62956 8968 62996 9008
rect 62092 8296 62132 8336
rect 63628 8212 63668 8252
rect 62092 7960 62132 8000
rect 61708 7372 61748 7412
rect 62668 7876 62708 7916
rect 62380 7540 62420 7580
rect 61324 6532 61364 6572
rect 61900 7204 61940 7244
rect 61900 6532 61940 6572
rect 61900 6364 61940 6404
rect 62188 7204 62228 7244
rect 61420 6280 61460 6320
rect 61228 6196 61268 6236
rect 61324 5944 61364 5984
rect 61228 5692 61268 5732
rect 62092 6280 62132 6320
rect 61804 5944 61844 5984
rect 61996 5944 62036 5984
rect 61132 5608 61172 5648
rect 62284 6364 62324 6404
rect 61900 5524 61940 5564
rect 60940 5188 60980 5228
rect 60172 4264 60212 4304
rect 60076 4012 60116 4052
rect 60268 3508 60308 3548
rect 60268 3172 60308 3212
rect 59980 2668 60020 2708
rect 60460 4169 60500 4209
rect 60460 4012 60500 4052
rect 63052 7204 63092 7244
rect 62476 7120 62516 7160
rect 62668 6364 62708 6404
rect 63148 6364 63188 6404
rect 61996 5356 62036 5396
rect 61804 5188 61844 5228
rect 62668 5440 62708 5480
rect 62764 5356 62804 5396
rect 62956 5524 62996 5564
rect 62860 5188 62900 5228
rect 62764 5020 62804 5060
rect 62956 5020 62996 5060
rect 61228 4516 61268 4556
rect 61228 4348 61268 4388
rect 60652 4012 60692 4052
rect 60652 3760 60692 3800
rect 59980 2500 60020 2540
rect 59308 2248 59348 2288
rect 59116 2164 59156 2204
rect 59404 1996 59444 2036
rect 59212 1072 59252 1112
rect 60364 2500 60404 2540
rect 59788 1156 59828 1196
rect 60460 2332 60500 2372
rect 60364 1828 60404 1868
rect 60172 820 60212 860
rect 60556 1744 60596 1784
rect 61132 3676 61172 3716
rect 60748 3424 60788 3464
rect 61228 3508 61268 3548
rect 60748 3172 60788 3212
rect 61228 2836 61268 2876
rect 61132 2416 61172 2456
rect 60940 1576 60980 1616
rect 60940 988 60980 1028
rect 61612 4684 61652 4724
rect 61900 4516 61940 4556
rect 61996 4096 62036 4136
rect 61516 3676 61556 3716
rect 61516 3004 61556 3044
rect 61420 1996 61460 2036
rect 61324 1408 61364 1448
rect 61324 904 61364 944
rect 61612 2164 61652 2204
rect 62476 4516 62516 4556
rect 62380 4432 62420 4472
rect 62284 4180 62324 4220
rect 62092 3844 62132 3884
rect 62284 3508 62324 3548
rect 61804 3088 61844 3128
rect 61996 3088 62036 3128
rect 61900 2836 61940 2876
rect 61708 1240 61748 1280
rect 61996 1156 62036 1196
rect 62188 3088 62228 3128
rect 62092 1072 62132 1112
rect 62284 2920 62324 2960
rect 62284 2332 62324 2372
rect 62380 820 62420 860
rect 62572 3760 62612 3800
rect 62572 3340 62612 3380
rect 62860 4684 62900 4724
rect 62764 4600 62804 4640
rect 62764 3340 62804 3380
rect 62668 2416 62708 2456
rect 62668 1156 62708 1196
rect 63052 4516 63092 4556
rect 63052 3844 63092 3884
rect 63532 5608 63572 5648
rect 65408 9052 65448 9092
rect 65490 9052 65530 9092
rect 65572 9052 65612 9092
rect 65654 9052 65694 9092
rect 65736 9052 65776 9092
rect 66124 9052 66164 9092
rect 64012 8800 64052 8840
rect 64972 8632 65012 8672
rect 64168 8296 64208 8336
rect 64250 8296 64290 8336
rect 64332 8296 64372 8336
rect 64414 8296 64454 8336
rect 64496 8296 64536 8336
rect 64684 8044 64724 8084
rect 64012 7288 64052 7328
rect 64492 7204 64532 7244
rect 66412 8128 66452 8168
rect 65260 7876 65300 7916
rect 65836 7792 65876 7832
rect 65408 7540 65448 7580
rect 65490 7540 65530 7580
rect 65572 7540 65612 7580
rect 65654 7540 65694 7580
rect 65736 7540 65776 7580
rect 64012 7036 64052 7076
rect 64972 6868 65012 6908
rect 64168 6784 64208 6824
rect 64250 6784 64290 6824
rect 64332 6784 64372 6824
rect 64414 6784 64454 6824
rect 64496 6784 64536 6824
rect 65164 6784 65204 6824
rect 64780 6448 64820 6488
rect 65260 6364 65300 6404
rect 64780 6280 64820 6320
rect 64972 6280 65012 6320
rect 65068 6112 65108 6152
rect 63916 5860 63956 5900
rect 65408 6028 65448 6068
rect 65490 6028 65530 6068
rect 65572 6028 65612 6068
rect 65654 6028 65694 6068
rect 65736 6028 65776 6068
rect 65260 5944 65300 5984
rect 63244 5440 63284 5480
rect 63244 4852 63284 4892
rect 63436 4852 63476 4892
rect 63532 4432 63572 4472
rect 63436 4348 63476 4388
rect 63340 3844 63380 3884
rect 63724 4432 63764 4472
rect 63628 4012 63668 4052
rect 63244 3424 63284 3464
rect 63148 3256 63188 3296
rect 64588 5692 64628 5732
rect 64012 5608 64052 5648
rect 64168 5272 64208 5312
rect 64250 5272 64290 5312
rect 64332 5272 64372 5312
rect 64414 5272 64454 5312
rect 64496 5272 64536 5312
rect 64012 5188 64052 5228
rect 63916 3508 63956 3548
rect 63532 3256 63572 3296
rect 63436 3172 63476 3212
rect 63340 2332 63380 2372
rect 63244 1828 63284 1868
rect 63244 1660 63284 1700
rect 64780 5020 64820 5060
rect 64108 4684 64148 4724
rect 64204 4432 64244 4472
rect 64396 4936 64436 4976
rect 64588 4936 64628 4976
rect 64396 4684 64436 4724
rect 64300 4348 64340 4388
rect 64588 4180 64628 4220
rect 64780 4180 64820 4220
rect 64588 3928 64628 3968
rect 64168 3760 64208 3800
rect 64250 3760 64290 3800
rect 64332 3760 64372 3800
rect 64414 3760 64454 3800
rect 64496 3760 64536 3800
rect 63916 3088 63956 3128
rect 63916 2920 63956 2960
rect 63820 2752 63860 2792
rect 63724 988 63764 1028
rect 63916 2668 63956 2708
rect 65452 5524 65492 5564
rect 65408 4516 65448 4556
rect 65490 4516 65530 4556
rect 65572 4516 65612 4556
rect 65654 4516 65694 4556
rect 65736 4516 65776 4556
rect 66220 7624 66260 7664
rect 66220 7120 66260 7160
rect 66796 7204 66836 7244
rect 66604 6448 66644 6488
rect 66412 5692 66452 5732
rect 64780 4012 64820 4052
rect 64684 3844 64724 3884
rect 64876 3844 64916 3884
rect 64780 3760 64820 3800
rect 64396 3172 64436 3212
rect 64300 2920 64340 2960
rect 64012 1240 64052 1280
rect 64396 2164 64436 2204
rect 64588 3172 64628 3212
rect 64588 2836 64628 2876
rect 64204 1576 64244 1616
rect 64108 904 64148 944
rect 64780 3256 64820 3296
rect 64972 3676 65012 3716
rect 65260 3760 65300 3800
rect 65452 3760 65492 3800
rect 64972 3508 65012 3548
rect 64972 2920 65012 2960
rect 64684 1156 64724 1196
rect 65164 3424 65204 3464
rect 65644 4180 65684 4220
rect 65836 3928 65876 3968
rect 66028 4348 66068 4388
rect 66028 4096 66068 4136
rect 65932 3760 65972 3800
rect 66508 5440 66548 5480
rect 66412 4096 66452 4136
rect 66220 3928 66260 3968
rect 66220 3676 66260 3716
rect 65740 3172 65780 3212
rect 65408 3004 65448 3044
rect 65490 3004 65530 3044
rect 65572 3004 65612 3044
rect 65654 3004 65694 3044
rect 65736 3004 65776 3044
rect 65356 2584 65396 2624
rect 65068 1240 65108 1280
rect 65932 3424 65972 3464
rect 66028 3172 66068 3212
rect 65932 2668 65972 2708
rect 66124 2752 66164 2792
rect 66316 3508 66356 3548
rect 66508 3340 66548 3380
rect 66316 3172 66356 3212
rect 66028 1660 66068 1700
rect 65932 1240 65972 1280
rect 66508 2752 66548 2792
rect 66412 1576 66452 1616
rect 66988 8716 67028 8756
rect 67180 8716 67220 8756
rect 67852 7960 67892 8000
rect 67180 7876 67220 7916
rect 67660 7876 67700 7916
rect 67372 7708 67412 7748
rect 70060 9220 70100 9260
rect 68716 8884 68756 8924
rect 70732 9388 70772 9428
rect 70540 9136 70580 9176
rect 71212 9136 71252 9176
rect 70156 8716 70196 8756
rect 70924 8800 70964 8840
rect 68908 7876 68948 7916
rect 69772 7876 69812 7916
rect 69964 7876 70004 7916
rect 69772 7540 69812 7580
rect 68044 7204 68084 7244
rect 66988 7036 67028 7076
rect 67084 6868 67124 6908
rect 67180 6532 67220 6572
rect 67084 6364 67124 6404
rect 67372 6364 67412 6404
rect 66988 5608 67028 5648
rect 67180 4936 67220 4976
rect 67756 6364 67796 6404
rect 67948 7036 67988 7076
rect 68044 6784 68084 6824
rect 68236 7120 68276 7160
rect 68140 6364 68180 6404
rect 67372 4852 67412 4892
rect 66892 4768 66932 4808
rect 66892 4432 66932 4472
rect 66700 3676 66740 3716
rect 67564 5272 67604 5312
rect 67852 5776 67892 5816
rect 68044 5692 68084 5732
rect 68236 6196 68276 6236
rect 68140 5608 68180 5648
rect 67756 5188 67796 5228
rect 67660 5020 67700 5060
rect 67564 4600 67604 4640
rect 67084 4264 67124 4304
rect 67276 4264 67316 4304
rect 67084 3760 67124 3800
rect 66988 3424 67028 3464
rect 66700 3340 66740 3380
rect 67084 3340 67124 3380
rect 66796 2836 66836 2876
rect 66988 2836 67028 2876
rect 67468 4264 67508 4304
rect 67756 4852 67796 4892
rect 68044 5104 68084 5144
rect 67948 4936 67988 4976
rect 68140 4936 68180 4976
rect 67756 4432 67796 4472
rect 67948 4264 67988 4304
rect 68044 4180 68084 4220
rect 68145 4180 68180 4220
rect 68180 4180 68185 4220
rect 67276 2920 67316 2960
rect 66892 1324 66932 1364
rect 68140 3928 68180 3968
rect 67756 3844 67796 3884
rect 67852 3760 67892 3800
rect 67468 3424 67508 3464
rect 68140 3676 68180 3716
rect 68044 2668 68084 2708
rect 67660 2584 67700 2624
rect 68716 7204 68756 7244
rect 68332 5944 68372 5984
rect 68332 5692 68372 5732
rect 68332 5440 68372 5480
rect 68620 6616 68660 6656
rect 68524 6364 68564 6404
rect 68812 6532 68852 6572
rect 69196 7204 69236 7244
rect 68908 6280 68948 6320
rect 68716 6112 68756 6152
rect 68908 6112 68948 6152
rect 68716 5944 68756 5984
rect 68428 5020 68468 5060
rect 68524 4852 68564 4892
rect 68332 4768 68372 4808
rect 68908 5608 68948 5648
rect 69100 6448 69140 6488
rect 69676 6532 69716 6572
rect 70348 7960 70388 8000
rect 70156 7876 70196 7916
rect 70636 8632 70676 8672
rect 70732 8044 70772 8084
rect 70540 7876 70580 7916
rect 71020 8548 71060 8588
rect 71116 8212 71156 8252
rect 70924 7876 70964 7916
rect 70252 7792 70292 7832
rect 70732 7708 70772 7748
rect 70060 6700 70100 6740
rect 69196 6196 69236 6236
rect 69388 6196 69428 6236
rect 69388 5776 69428 5816
rect 68812 4768 68852 4808
rect 68332 4264 68372 4304
rect 68524 4516 68564 4556
rect 68428 4096 68468 4136
rect 68524 4012 68564 4052
rect 68716 4264 68756 4304
rect 68524 3676 68564 3716
rect 69004 4348 69044 4388
rect 68908 4264 68948 4304
rect 69004 4096 69044 4136
rect 68428 3172 68468 3212
rect 68236 2920 68276 2960
rect 69100 4012 69140 4052
rect 69388 5440 69428 5480
rect 69292 5356 69332 5396
rect 69292 4684 69332 4724
rect 69292 4264 69332 4304
rect 68812 2752 68852 2792
rect 68812 2584 68852 2624
rect 67372 1240 67412 1280
rect 67468 1072 67508 1112
rect 67660 820 67700 860
rect 68236 1828 68276 1868
rect 68044 1576 68084 1616
rect 68620 1156 68660 1196
rect 69196 1324 69236 1364
rect 69196 988 69236 1028
rect 69772 5692 69812 5732
rect 69580 5524 69620 5564
rect 69580 5104 69620 5144
rect 69772 5272 69812 5312
rect 69676 4936 69716 4976
rect 69772 4852 69812 4892
rect 69964 5860 70004 5900
rect 69964 5440 70004 5480
rect 70156 6196 70196 6236
rect 70156 5776 70196 5816
rect 70636 6028 70676 6068
rect 70060 5356 70100 5396
rect 69580 4432 69620 4472
rect 69484 4096 69524 4136
rect 69580 4012 69620 4052
rect 69388 3424 69428 3464
rect 69580 2836 69620 2876
rect 69388 1240 69428 1280
rect 69292 820 69332 860
rect 70156 4852 70196 4892
rect 69964 4600 70004 4640
rect 69868 4516 69908 4556
rect 70060 4516 70100 4556
rect 70060 4264 70100 4304
rect 70060 3760 70100 3800
rect 70348 5020 70388 5060
rect 70540 5440 70580 5480
rect 70636 5356 70676 5396
rect 71020 6280 71060 6320
rect 72172 9724 72212 9764
rect 72076 9556 72116 9596
rect 71788 9388 71828 9428
rect 71596 9304 71636 9344
rect 71980 9304 72020 9344
rect 72172 8968 72212 9008
rect 72076 8128 72116 8168
rect 71500 7372 71540 7412
rect 71500 6616 71540 6656
rect 71404 6364 71444 6404
rect 71308 6280 71348 6320
rect 71308 5692 71348 5732
rect 70924 5440 70964 5480
rect 70828 5356 70868 5396
rect 70924 4936 70964 4976
rect 70540 4852 70580 4892
rect 70828 4852 70868 4892
rect 70444 4768 70484 4808
rect 70732 4684 70772 4724
rect 70252 4180 70292 4220
rect 70156 3592 70196 3632
rect 70252 3508 70292 3548
rect 70444 4180 70484 4220
rect 70444 4012 70484 4052
rect 70636 4012 70676 4052
rect 70636 3844 70676 3884
rect 69772 2332 69812 2372
rect 69676 1828 69716 1868
rect 69964 1072 70004 1112
rect 69964 904 70004 944
rect 71116 4852 71156 4892
rect 71308 4852 71348 4892
rect 70924 4684 70964 4724
rect 71212 4684 71252 4724
rect 71500 5944 71540 5984
rect 71500 5356 71540 5396
rect 71692 7876 71732 7916
rect 71884 7372 71924 7412
rect 71788 6616 71828 6656
rect 71788 6364 71828 6404
rect 71692 5860 71732 5900
rect 71692 5608 71732 5648
rect 71596 5188 71636 5228
rect 71692 5020 71732 5060
rect 71020 4348 71060 4388
rect 70828 4180 70868 4220
rect 71212 4180 71252 4220
rect 71308 4096 71348 4136
rect 71404 4012 71444 4052
rect 71020 3928 71060 3968
rect 71404 3760 71444 3800
rect 70924 3592 70964 3632
rect 71692 4852 71732 4892
rect 71596 4600 71636 4640
rect 71596 4432 71636 4472
rect 71788 4180 71828 4220
rect 71788 3928 71828 3968
rect 71788 3592 71828 3632
rect 70550 3256 70590 3296
rect 83116 10900 83156 10940
rect 80528 10564 80568 10604
rect 80610 10564 80650 10604
rect 80692 10564 80732 10604
rect 80774 10564 80814 10604
rect 80856 10564 80896 10604
rect 95648 10564 95688 10604
rect 95730 10564 95770 10604
rect 95812 10564 95852 10604
rect 95894 10564 95934 10604
rect 95976 10564 96016 10604
rect 73804 10480 73844 10520
rect 73996 10480 74036 10520
rect 77068 10480 77108 10520
rect 78028 10480 78068 10520
rect 82828 10480 82868 10520
rect 84076 10480 84116 10520
rect 88300 10480 88340 10520
rect 92812 10480 92852 10520
rect 73132 10312 73172 10352
rect 73324 10228 73364 10268
rect 73516 10228 73556 10268
rect 76492 10312 76532 10352
rect 73132 10060 73172 10100
rect 72940 9976 72980 10016
rect 73228 9976 73268 10016
rect 73804 9640 73844 9680
rect 73036 9472 73076 9512
rect 73228 9472 73268 9512
rect 73708 9472 73748 9512
rect 72940 9304 72980 9344
rect 72940 8968 72980 9008
rect 72556 8128 72596 8168
rect 72748 7876 72788 7916
rect 72844 7456 72884 7496
rect 72364 7204 72404 7244
rect 71980 6616 72020 6656
rect 72844 6868 72884 6908
rect 72652 6616 72692 6656
rect 71980 6196 72020 6236
rect 72364 6196 72404 6236
rect 73036 8884 73076 8924
rect 74188 9640 74228 9680
rect 73324 9052 73364 9092
rect 73708 8884 73748 8924
rect 73420 8380 73460 8420
rect 73324 8296 73364 8336
rect 73420 7624 73460 7664
rect 73036 6280 73076 6320
rect 72940 6196 72980 6236
rect 73516 6196 73556 6236
rect 73228 6028 73268 6068
rect 72748 5944 72788 5984
rect 73516 5944 73556 5984
rect 72076 5860 72116 5900
rect 71980 5356 72020 5396
rect 72364 5440 72404 5480
rect 72556 5440 72596 5480
rect 72748 5524 72788 5564
rect 72652 5356 72692 5396
rect 72652 5188 72692 5228
rect 72172 5020 72212 5060
rect 72556 5020 72596 5060
rect 72364 4936 72404 4976
rect 72076 4768 72116 4808
rect 72172 4684 72212 4724
rect 72076 4516 72116 4556
rect 71980 4432 72020 4472
rect 72268 4348 72308 4388
rect 72172 4180 72212 4220
rect 72172 3928 72212 3968
rect 71980 3760 72020 3800
rect 71884 3340 71924 3380
rect 71308 3256 71348 3296
rect 71788 3256 71828 3296
rect 70444 2332 70484 2372
rect 70348 1576 70388 1616
rect 70348 484 70388 524
rect 71212 3172 71252 3212
rect 71116 2584 71156 2624
rect 70924 1996 70964 2036
rect 70828 1576 70868 1616
rect 70732 1156 70772 1196
rect 71308 1660 71348 1700
rect 71596 2584 71636 2624
rect 71500 988 71540 1028
rect 71692 1492 71732 1532
rect 71884 1240 71924 1280
rect 72076 3508 72116 3548
rect 72364 4180 72404 4220
rect 72076 2668 72116 2708
rect 72556 4516 72596 4556
rect 73420 5692 73460 5732
rect 73612 5692 73652 5732
rect 73228 5608 73268 5648
rect 72940 5440 72980 5480
rect 73516 5608 73556 5648
rect 73228 5356 73268 5396
rect 73516 5104 73556 5144
rect 72844 5020 72884 5060
rect 73132 4936 73172 4976
rect 74476 10228 74516 10268
rect 74380 10060 74420 10100
rect 74284 9472 74324 9512
rect 75436 9136 75476 9176
rect 74668 8968 74708 9008
rect 75052 8800 75092 8840
rect 74764 8716 74804 8756
rect 74572 8548 74612 8588
rect 74380 8296 74420 8336
rect 77644 10396 77684 10436
rect 77260 10228 77300 10268
rect 77452 10144 77492 10184
rect 76684 9220 76724 9260
rect 76588 8884 76628 8924
rect 76012 8800 76052 8840
rect 75148 8716 75188 8756
rect 75532 8716 75572 8756
rect 75340 8632 75380 8672
rect 75148 8464 75188 8504
rect 74956 8212 74996 8252
rect 75052 8128 75092 8168
rect 73996 7960 74036 8000
rect 74188 7876 74228 7916
rect 73996 7708 74036 7748
rect 74380 8044 74420 8084
rect 74572 7876 74612 7916
rect 74860 7540 74900 7580
rect 74764 7456 74804 7496
rect 74476 7372 74516 7412
rect 74284 7036 74324 7076
rect 74188 6952 74228 6992
rect 74284 6784 74324 6824
rect 73996 6616 74036 6656
rect 74188 6616 74228 6656
rect 74092 6532 74132 6572
rect 75052 7540 75092 7580
rect 74956 7372 74996 7412
rect 74565 7120 74605 7160
rect 74476 6952 74516 6992
rect 74956 6784 74996 6824
rect 73900 6196 73940 6236
rect 74092 6364 74132 6404
rect 74668 6448 74708 6488
rect 74572 6364 74612 6404
rect 74380 6280 74420 6320
rect 73804 6028 73844 6068
rect 73996 6028 74036 6068
rect 73900 5944 73940 5984
rect 73996 5692 74036 5732
rect 74668 6280 74708 6320
rect 74284 5776 74324 5816
rect 74476 5692 74516 5732
rect 73900 5272 73940 5312
rect 74188 5356 74228 5396
rect 73996 5104 74036 5144
rect 72940 4852 72980 4892
rect 73612 4852 73652 4892
rect 73324 4768 73364 4808
rect 72844 4684 72884 4724
rect 72748 4600 72788 4640
rect 72940 4516 72980 4556
rect 72748 4180 72788 4220
rect 73228 4432 73268 4472
rect 72556 4096 72596 4136
rect 73132 4096 73172 4136
rect 73132 3592 73172 3632
rect 72556 3340 72596 3380
rect 73516 4348 73556 4388
rect 73324 4180 73364 4220
rect 73516 4012 73556 4052
rect 72460 3256 72500 3296
rect 72844 3256 72884 3296
rect 73132 3256 73172 3296
rect 72460 2080 72500 2120
rect 72268 904 72308 944
rect 72556 1996 72596 2036
rect 72748 3088 72788 3128
rect 72652 484 72692 524
rect 72844 1744 72884 1784
rect 73516 3592 73556 3632
rect 73420 3172 73460 3212
rect 73900 4684 73940 4724
rect 73708 4516 73748 4556
rect 73900 4096 73940 4136
rect 73900 3760 73940 3800
rect 73708 3508 73748 3548
rect 74188 4936 74228 4976
rect 74476 5524 74516 5564
rect 74476 5272 74516 5312
rect 74092 4600 74132 4640
rect 74476 4264 74516 4304
rect 74380 4096 74420 4136
rect 74668 5692 74708 5732
rect 74668 4264 74708 4304
rect 74188 3424 74228 3464
rect 73324 1828 73364 1868
rect 73036 1576 73076 1616
rect 73228 1240 73268 1280
rect 73036 1156 73076 1196
rect 74188 2584 74228 2624
rect 74956 6196 74996 6236
rect 75244 8128 75284 8168
rect 75916 8128 75956 8168
rect 75244 7624 75284 7664
rect 75916 7792 75956 7832
rect 75820 7624 75860 7664
rect 75436 7540 75476 7580
rect 77356 9976 77396 10016
rect 82444 10312 82484 10352
rect 77836 10144 77876 10184
rect 78028 10144 78068 10184
rect 77644 10060 77684 10100
rect 82732 10060 82772 10100
rect 77452 9640 77492 9680
rect 76972 9388 77012 9428
rect 76780 8464 76820 8504
rect 76876 8380 76916 8420
rect 76876 8128 76916 8168
rect 76300 7792 76340 7832
rect 75244 7120 75284 7160
rect 75148 6868 75188 6908
rect 75628 6952 75668 6992
rect 75340 6700 75380 6740
rect 75340 6448 75380 6488
rect 75148 6280 75188 6320
rect 74956 5692 74996 5732
rect 75052 5524 75092 5564
rect 75052 5272 75092 5312
rect 74860 4768 74900 4808
rect 75340 6112 75380 6152
rect 75244 5692 75284 5732
rect 75148 4852 75188 4892
rect 75148 4600 75188 4640
rect 75532 5608 75572 5648
rect 75532 4600 75572 4640
rect 75052 4096 75092 4136
rect 74860 4012 74900 4052
rect 74380 3004 74420 3044
rect 74284 2080 74324 2120
rect 73804 1660 73844 1700
rect 74188 1660 74228 1700
rect 73804 1408 73844 1448
rect 73612 904 73652 944
rect 73996 820 74036 860
rect 74764 2920 74804 2960
rect 74572 1492 74612 1532
rect 74572 1072 74612 1112
rect 74956 2668 74996 2708
rect 74956 2500 74996 2540
rect 75244 4096 75284 4136
rect 75148 3424 75188 3464
rect 75916 5524 75956 5564
rect 75820 5020 75860 5060
rect 75928 5020 75968 5060
rect 75724 4684 75764 4724
rect 76780 7624 76820 7664
rect 76876 7120 76916 7160
rect 76780 6532 76820 6572
rect 76684 5860 76724 5900
rect 76876 5608 76916 5648
rect 76108 5440 76148 5480
rect 76396 5356 76436 5396
rect 76108 5104 76148 5144
rect 76012 4516 76052 4556
rect 75820 4348 75860 4388
rect 75628 4096 75668 4136
rect 75532 4012 75572 4052
rect 75628 3844 75668 3884
rect 75532 3760 75572 3800
rect 75436 3592 75476 3632
rect 75340 3172 75380 3212
rect 75244 3004 75284 3044
rect 75148 2752 75188 2792
rect 75052 1156 75092 1196
rect 75532 2416 75572 2456
rect 75820 4180 75860 4220
rect 76012 4180 76052 4220
rect 76300 4936 76340 4976
rect 76396 4852 76436 4892
rect 76204 4768 76244 4808
rect 76300 4684 76340 4724
rect 76396 4264 76436 4304
rect 76108 4096 76148 4136
rect 76396 4096 76436 4136
rect 75628 1996 75668 2036
rect 75916 3004 75956 3044
rect 75916 2248 75956 2288
rect 75724 1744 75764 1784
rect 75724 988 75764 1028
rect 76108 2500 76148 2540
rect 76012 1240 76052 1280
rect 76876 5272 76916 5312
rect 76780 5104 76820 5144
rect 76588 4936 76628 4976
rect 77164 9220 77204 9260
rect 79288 9808 79328 9848
rect 79370 9808 79410 9848
rect 79452 9808 79492 9848
rect 79534 9808 79574 9848
rect 79616 9808 79656 9848
rect 77932 9724 77972 9764
rect 80620 9724 80660 9764
rect 77740 9556 77780 9596
rect 77548 9220 77588 9260
rect 77356 9052 77396 9092
rect 78412 9052 78452 9092
rect 78220 8884 78260 8924
rect 77932 8716 77972 8756
rect 77164 8464 77204 8504
rect 77068 7540 77108 7580
rect 77068 6532 77108 6572
rect 77068 6196 77108 6236
rect 77068 5608 77108 5648
rect 77548 7960 77588 8000
rect 77740 7876 77780 7916
rect 77452 7624 77492 7664
rect 77260 7204 77300 7244
rect 77548 7204 77588 7244
rect 77356 6868 77396 6908
rect 77548 6616 77588 6656
rect 77740 7288 77780 7328
rect 77740 6868 77780 6908
rect 77644 6532 77684 6572
rect 77452 6448 77492 6488
rect 77740 6448 77780 6488
rect 78220 8716 78260 8756
rect 78124 8212 78164 8252
rect 78507 8548 78547 8588
rect 78412 8464 78452 8504
rect 78412 7876 78452 7916
rect 78028 7792 78068 7832
rect 77932 7708 77972 7748
rect 80236 9388 80276 9428
rect 81868 9556 81908 9596
rect 80812 9388 80852 9428
rect 81004 9388 81044 9428
rect 82060 9472 82100 9512
rect 80528 9052 80568 9092
rect 80610 9052 80650 9092
rect 80692 9052 80732 9092
rect 80774 9052 80814 9092
rect 80856 9052 80896 9092
rect 81196 9304 81236 9344
rect 81484 9304 81524 9344
rect 81100 9052 81140 9092
rect 78796 8800 78836 8840
rect 78988 8800 79028 8840
rect 80908 8800 80948 8840
rect 78892 8716 78932 8756
rect 78700 8632 78740 8672
rect 80812 8716 80852 8756
rect 78988 8296 79028 8336
rect 79288 8296 79328 8336
rect 79370 8296 79410 8336
rect 79452 8296 79492 8336
rect 79534 8296 79574 8336
rect 79616 8296 79656 8336
rect 78988 8044 79028 8084
rect 78316 7624 78356 7664
rect 78028 7120 78068 7160
rect 77164 5104 77204 5144
rect 76780 4684 76820 4724
rect 76684 4516 76724 4556
rect 76588 4348 76628 4388
rect 76780 4348 76820 4388
rect 76780 4180 76820 4220
rect 76684 4096 76724 4136
rect 76684 3592 76724 3632
rect 76300 3424 76340 3464
rect 76300 1156 76340 1196
rect 76204 820 76244 860
rect 76492 2836 76532 2876
rect 76396 904 76436 944
rect 77452 5440 77492 5480
rect 77356 5356 77396 5396
rect 77836 5440 77876 5480
rect 77548 5188 77588 5228
rect 77740 5188 77780 5228
rect 77452 5104 77492 5144
rect 76972 4852 77012 4892
rect 77260 4852 77300 4892
rect 77164 4348 77204 4388
rect 77164 4096 77204 4136
rect 77068 3844 77108 3884
rect 77356 4180 77396 4220
rect 77356 3592 77396 3632
rect 76972 3256 77012 3296
rect 76588 2416 76628 2456
rect 76780 2416 76820 2456
rect 76684 2332 76724 2372
rect 76876 1408 76916 1448
rect 77164 2248 77204 2288
rect 77260 1660 77300 1700
rect 77836 4852 77876 4892
rect 77644 4264 77684 4304
rect 77740 3760 77780 3800
rect 77068 988 77108 1028
rect 77452 1240 77492 1280
rect 78220 6532 78260 6572
rect 78028 6448 78068 6488
rect 78028 5440 78068 5480
rect 78028 5104 78068 5144
rect 78028 3844 78068 3884
rect 78508 7288 78548 7328
rect 78796 7876 78836 7916
rect 80908 8464 80948 8504
rect 81004 8380 81044 8420
rect 81004 8212 81044 8252
rect 80908 8128 80948 8168
rect 80716 7876 80756 7916
rect 81292 8884 81332 8924
rect 81196 8716 81236 8756
rect 81676 9220 81716 9260
rect 81484 8800 81524 8840
rect 81868 9136 81908 9176
rect 82060 8968 82100 9008
rect 81580 8716 81620 8756
rect 81388 8632 81428 8672
rect 81964 8716 82004 8756
rect 82156 8716 82196 8756
rect 81772 8548 81812 8588
rect 81580 8296 81620 8336
rect 81772 8128 81812 8168
rect 81676 8044 81716 8084
rect 80812 7792 80852 7832
rect 78892 7372 78932 7412
rect 78700 7288 78740 7328
rect 78604 7204 78644 7244
rect 78508 7036 78548 7076
rect 78412 6280 78452 6320
rect 78988 6952 79028 6992
rect 78700 6868 78740 6908
rect 78604 6616 78644 6656
rect 78508 6112 78548 6152
rect 78412 6028 78452 6068
rect 78508 5944 78548 5984
rect 78412 5692 78452 5732
rect 78316 5608 78356 5648
rect 78412 5440 78452 5480
rect 78220 3760 78260 3800
rect 78220 3508 78260 3548
rect 77740 3088 77780 3128
rect 78028 2920 78068 2960
rect 78508 5020 78548 5060
rect 80528 7540 80568 7580
rect 80610 7540 80650 7580
rect 80692 7540 80732 7580
rect 80774 7540 80814 7580
rect 80856 7540 80896 7580
rect 80428 7456 80468 7496
rect 79180 7372 79220 7412
rect 79180 6952 79220 6992
rect 79180 6784 79220 6824
rect 79288 6784 79328 6824
rect 79370 6784 79410 6824
rect 79452 6784 79492 6824
rect 79534 6784 79574 6824
rect 79616 6784 79656 6824
rect 78796 6448 78836 6488
rect 78700 6364 78740 6404
rect 78796 6112 78836 6152
rect 78892 6028 78932 6068
rect 78892 5860 78932 5900
rect 78796 5692 78836 5732
rect 78700 5440 78740 5480
rect 78796 5104 78836 5144
rect 79468 6616 79508 6656
rect 79276 6532 79316 6572
rect 79852 6532 79892 6572
rect 79084 6028 79124 6068
rect 79660 6196 79700 6236
rect 79372 6028 79412 6068
rect 79084 5692 79124 5732
rect 79468 5692 79508 5732
rect 80140 6448 80180 6488
rect 80044 6028 80084 6068
rect 79852 5692 79892 5732
rect 80044 5692 80084 5732
rect 79276 5608 79316 5648
rect 79756 5440 79796 5480
rect 79084 5272 79124 5312
rect 79288 5272 79328 5312
rect 79370 5272 79410 5312
rect 79452 5272 79492 5312
rect 79534 5272 79574 5312
rect 79616 5272 79656 5312
rect 78412 4180 78452 4220
rect 78795 4096 78835 4136
rect 78700 3592 78740 3632
rect 78604 3424 78644 3464
rect 78796 3424 78836 3464
rect 78988 4432 79028 4472
rect 79372 5104 79412 5144
rect 79276 4936 79316 4976
rect 79564 5104 79604 5144
rect 79468 5020 79508 5060
rect 79276 4432 79316 4472
rect 79084 4264 79124 4304
rect 78988 4096 79028 4136
rect 78988 3760 79028 3800
rect 79564 3928 79604 3968
rect 79852 5188 79892 5228
rect 79852 5020 79892 5060
rect 80044 5020 80084 5060
rect 80044 4096 80084 4136
rect 80332 6448 80372 6488
rect 82156 8044 82196 8084
rect 81099 7876 81100 7916
rect 81100 7876 81139 7916
rect 80812 7288 80852 7328
rect 80236 6280 80276 6320
rect 80236 5776 80276 5816
rect 80428 6280 80468 6320
rect 81484 7876 81524 7916
rect 82060 7960 82100 8000
rect 81868 7876 81908 7916
rect 81388 7792 81428 7832
rect 81292 7708 81332 7748
rect 81292 6700 81332 6740
rect 80528 6028 80568 6068
rect 80610 6028 80650 6068
rect 80692 6028 80732 6068
rect 80774 6028 80814 6068
rect 80856 6028 80896 6068
rect 81100 6028 81140 6068
rect 80428 5692 80468 5732
rect 80908 5860 80948 5900
rect 80812 5776 80852 5816
rect 80620 5608 80660 5648
rect 80620 5440 80660 5480
rect 80908 5692 80948 5732
rect 80812 5104 80852 5144
rect 80908 4936 80948 4976
rect 81100 5272 81140 5312
rect 81964 6448 82004 6488
rect 81971 6196 82011 6236
rect 81388 5860 81428 5900
rect 81292 5692 81332 5732
rect 81484 5692 81524 5732
rect 81388 5608 81428 5648
rect 79288 3760 79328 3800
rect 79370 3760 79410 3800
rect 79452 3760 79492 3800
rect 79534 3760 79574 3800
rect 79616 3760 79656 3800
rect 79852 3928 79892 3968
rect 79276 3508 79316 3548
rect 79180 3340 79220 3380
rect 78412 2752 78452 2792
rect 78028 2332 78068 2372
rect 78220 2332 78260 2372
rect 77644 1072 77684 1112
rect 77644 904 77684 944
rect 77836 736 77876 776
rect 78412 2248 78452 2288
rect 78604 2164 78644 2204
rect 78892 2752 78932 2792
rect 78796 820 78836 860
rect 79180 1156 79220 1196
rect 79372 3424 79412 3464
rect 79564 2836 79604 2876
rect 79756 3340 79796 3380
rect 79660 2332 79700 2372
rect 79756 1240 79796 1280
rect 79564 1072 79604 1112
rect 79372 148 79412 188
rect 79948 1240 79988 1280
rect 79852 988 79892 1028
rect 79756 652 79796 692
rect 80140 3424 80180 3464
rect 80428 4516 80468 4556
rect 80528 4516 80568 4556
rect 80610 4516 80650 4556
rect 80692 4516 80732 4556
rect 80774 4516 80814 4556
rect 80856 4516 80896 4556
rect 80428 4096 80468 4136
rect 80908 4348 80948 4388
rect 80620 4264 80660 4304
rect 80332 3928 80372 3968
rect 80236 2164 80276 2204
rect 80140 1156 80180 1196
rect 80044 736 80084 776
rect 80620 3844 80660 3884
rect 81004 4264 81044 4304
rect 80908 4096 80948 4136
rect 80716 3760 80756 3800
rect 80524 3424 80564 3464
rect 80528 3004 80568 3044
rect 80610 3004 80650 3044
rect 80692 3004 80732 3044
rect 80774 3004 80814 3044
rect 80856 3004 80896 3044
rect 80428 2248 80468 2288
rect 81484 5272 81524 5312
rect 81676 5440 81716 5480
rect 81676 5272 81716 5312
rect 81292 4684 81332 4724
rect 81580 5104 81620 5144
rect 81964 6028 82004 6068
rect 81868 5608 81908 5648
rect 81868 5440 81908 5480
rect 81964 5104 82004 5144
rect 81772 4852 81812 4892
rect 81484 4432 81524 4472
rect 81580 4264 81620 4304
rect 81292 4180 81332 4220
rect 81196 3760 81236 3800
rect 81100 3424 81140 3464
rect 81100 3172 81140 3212
rect 81004 2080 81044 2120
rect 80908 1408 80948 1448
rect 80524 1240 80564 1280
rect 80332 904 80372 944
rect 80332 736 80372 776
rect 80716 400 80756 440
rect 81772 4348 81812 4388
rect 81676 3256 81716 3296
rect 81196 1996 81236 2036
rect 81292 1912 81332 1952
rect 81484 1492 81524 1532
rect 81292 1324 81332 1364
rect 81292 988 81332 1028
rect 81868 1660 81908 1700
rect 82156 6868 82196 6908
rect 82348 8800 82388 8840
rect 82444 8548 82484 8588
rect 82732 9472 82772 9512
rect 83212 10312 83252 10352
rect 87148 10396 87188 10436
rect 83596 10228 83636 10268
rect 83980 10144 84020 10184
rect 83404 10060 83444 10100
rect 83788 10060 83828 10100
rect 83308 9976 83348 10016
rect 83212 9640 83252 9680
rect 83596 9052 83636 9092
rect 83884 9976 83924 10016
rect 83020 8632 83060 8672
rect 83692 8716 83732 8756
rect 83500 8632 83540 8672
rect 83404 8380 83444 8420
rect 82444 7899 82484 7916
rect 82444 7876 82484 7899
rect 82252 6616 82292 6656
rect 82348 6532 82388 6572
rect 82252 6448 82292 6488
rect 82156 5860 82196 5900
rect 82156 5524 82196 5564
rect 82156 4684 82196 4724
rect 82156 3928 82196 3968
rect 82060 3424 82100 3464
rect 82060 2332 82100 2372
rect 82060 1660 82100 1700
rect 81964 736 82004 776
rect 82348 6364 82388 6404
rect 82348 5776 82388 5816
rect 82348 5440 82388 5480
rect 82636 7792 82676 7832
rect 82636 7204 82676 7244
rect 82828 8044 82868 8084
rect 83020 8044 83060 8084
rect 83116 7960 83156 8000
rect 82828 7876 82868 7916
rect 83020 7792 83060 7832
rect 82924 7540 82964 7580
rect 83212 7876 83252 7916
rect 83404 7876 83444 7916
rect 83020 7204 83060 7244
rect 83308 7624 83348 7664
rect 83596 8128 83636 8168
rect 83788 8128 83828 8168
rect 83788 7960 83828 8000
rect 82828 7120 82868 7160
rect 82924 6952 82964 6992
rect 82828 6784 82868 6824
rect 83404 7204 83444 7244
rect 83788 7540 83828 7580
rect 84172 10060 84212 10100
rect 83980 9472 84020 9512
rect 83980 8800 84020 8840
rect 86860 9388 86900 9428
rect 89644 10396 89684 10436
rect 89932 10396 89972 10436
rect 89164 10312 89204 10352
rect 87532 9556 87572 9596
rect 86764 9304 86804 9344
rect 85996 9220 86036 9260
rect 85036 8884 85076 8924
rect 84364 8716 84404 8756
rect 84268 8632 84308 8672
rect 84268 8464 84308 8504
rect 83980 7876 84020 7916
rect 84172 7876 84212 7916
rect 83980 7624 84020 7664
rect 83884 7456 83924 7496
rect 84172 7624 84212 7664
rect 84076 7540 84116 7580
rect 84172 7456 84212 7496
rect 84844 7960 84884 8000
rect 84556 7876 84596 7916
rect 84460 7792 84500 7832
rect 84940 7876 84980 7916
rect 84748 7708 84788 7748
rect 84940 7708 84980 7748
rect 84076 7120 84116 7160
rect 83500 6952 83540 6992
rect 83116 6784 83156 6824
rect 83788 6784 83828 6824
rect 83116 6448 83156 6488
rect 82924 6364 82964 6404
rect 82636 6280 82676 6320
rect 82828 6280 82868 6320
rect 83020 6280 83060 6320
rect 82540 5944 82580 5984
rect 83116 5944 83156 5984
rect 82924 5860 82964 5900
rect 82828 5776 82868 5816
rect 82636 5608 82676 5648
rect 82540 5524 82580 5564
rect 82636 5188 82676 5228
rect 82252 3676 82292 3716
rect 82252 2668 82292 2708
rect 82444 4684 82484 4724
rect 82540 4096 82580 4136
rect 82732 5104 82772 5144
rect 83116 5188 83156 5228
rect 83020 5020 83060 5060
rect 82924 4852 82964 4892
rect 82732 4516 82772 4556
rect 82732 4096 82772 4136
rect 82444 3928 82484 3968
rect 82444 3676 82484 3716
rect 82636 3508 82676 3548
rect 82348 1408 82388 1448
rect 82636 1408 82676 1448
rect 82252 1324 82292 1364
rect 82156 652 82196 692
rect 82060 568 82100 608
rect 82444 820 82484 860
rect 83308 6532 83348 6572
rect 83404 6448 83444 6488
rect 83596 6448 83636 6488
rect 83308 6280 83348 6320
rect 83308 6112 83348 6152
rect 83692 6280 83732 6320
rect 83500 6112 83540 6152
rect 83884 6700 83924 6740
rect 84652 7036 84692 7076
rect 83980 6280 84020 6320
rect 83884 6112 83924 6152
rect 84172 6028 84212 6068
rect 83692 5860 83732 5900
rect 83884 5776 83924 5816
rect 83500 5440 83540 5480
rect 83500 4852 83540 4892
rect 83788 5692 83828 5732
rect 83884 5524 83924 5564
rect 84076 5944 84116 5984
rect 83980 5272 84020 5312
rect 84076 5020 84116 5060
rect 83404 4684 83444 4724
rect 83884 4684 83924 4724
rect 83788 4516 83828 4556
rect 83212 4096 83252 4136
rect 83212 3592 83252 3632
rect 82924 3508 82964 3548
rect 82828 3424 82868 3464
rect 83404 4348 83444 4388
rect 83692 4348 83732 4388
rect 83404 3676 83444 3716
rect 82732 1240 82772 1280
rect 83308 1996 83348 2036
rect 83020 1576 83060 1616
rect 82924 1072 82964 1112
rect 82828 232 82868 272
rect 83212 1072 83252 1112
rect 83404 1156 83444 1196
rect 83596 3760 83636 3800
rect 84076 4516 84116 4556
rect 83980 4264 84020 4304
rect 83884 3424 83924 3464
rect 84364 5692 84404 5732
rect 84844 6280 84884 6320
rect 85132 8464 85172 8504
rect 85900 8296 85940 8336
rect 85228 8044 85268 8084
rect 85324 7708 85364 7748
rect 85516 7372 85556 7412
rect 85708 7372 85748 7412
rect 85612 7204 85652 7244
rect 85708 7120 85748 7160
rect 85420 6532 85460 6572
rect 85324 6448 85364 6488
rect 84364 5272 84404 5312
rect 84268 5104 84308 5144
rect 84268 4852 84308 4892
rect 84268 4684 84308 4724
rect 84268 4516 84308 4556
rect 84652 4852 84692 4892
rect 84556 4516 84596 4556
rect 84460 4180 84500 4220
rect 84364 4096 84404 4136
rect 84364 3928 84404 3968
rect 84460 3760 84500 3800
rect 83692 2164 83732 2204
rect 83500 988 83540 1028
rect 83596 736 83636 776
rect 84172 3172 84212 3212
rect 85132 5860 85172 5900
rect 84556 1492 84596 1532
rect 83980 1240 84020 1280
rect 83788 484 83828 524
rect 83692 400 83732 440
rect 84172 1156 84212 1196
rect 84556 652 84596 692
rect 85036 4768 85076 4808
rect 84940 4684 84980 4724
rect 85132 4012 85172 4052
rect 85036 3928 85076 3968
rect 84940 3592 84980 3632
rect 85132 3592 85172 3632
rect 85132 3340 85172 3380
rect 84940 2416 84980 2456
rect 84844 1072 84884 1112
rect 85516 5776 85556 5816
rect 85324 5020 85364 5060
rect 85420 4516 85460 4556
rect 85324 4264 85364 4304
rect 85612 4852 85652 4892
rect 85516 4012 85556 4052
rect 85420 3340 85460 3380
rect 85804 7036 85844 7076
rect 85804 5524 85844 5564
rect 86092 8968 86132 9008
rect 85996 7120 86036 7160
rect 85996 4852 86036 4892
rect 85804 4684 85844 4724
rect 85708 4264 85748 4304
rect 85708 3340 85748 3380
rect 85324 2332 85364 2372
rect 85516 1996 85556 2036
rect 85228 1240 85268 1280
rect 85516 1240 85556 1280
rect 85324 988 85364 1028
rect 85900 3844 85940 3884
rect 87052 9304 87092 9344
rect 86956 8884 86996 8924
rect 86860 8716 86900 8756
rect 86860 7708 86900 7748
rect 86380 7204 86420 7244
rect 86284 7120 86324 7160
rect 86188 5608 86228 5648
rect 86860 7036 86900 7076
rect 86572 6952 86612 6992
rect 86476 6532 86516 6572
rect 86668 6280 86708 6320
rect 86572 5776 86612 5816
rect 86380 4348 86420 4388
rect 86572 4600 86612 4640
rect 86284 4096 86324 4136
rect 86956 5020 86996 5060
rect 87436 8800 87476 8840
rect 88012 10228 88052 10268
rect 88396 10228 88436 10268
rect 88204 10144 88244 10184
rect 87916 10060 87956 10100
rect 88108 9724 88148 9764
rect 87916 9472 87956 9512
rect 87820 9388 87860 9428
rect 87724 9304 87764 9344
rect 87724 8968 87764 9008
rect 87916 8800 87956 8840
rect 87628 8716 87668 8756
rect 87244 8632 87284 8672
rect 87532 8632 87572 8672
rect 87052 4936 87092 4976
rect 86764 4684 86804 4724
rect 86668 4516 86708 4556
rect 86860 4516 86900 4556
rect 86764 4264 86804 4304
rect 86092 3340 86132 3380
rect 85996 2584 86036 2624
rect 85900 2500 85940 2540
rect 85900 2332 85940 2372
rect 85612 568 85652 608
rect 86092 1492 86132 1532
rect 86860 3760 86900 3800
rect 86860 3508 86900 3548
rect 86860 3340 86900 3380
rect 86188 1324 86228 1364
rect 86668 2920 86708 2960
rect 86668 2584 86708 2624
rect 86572 2500 86612 2540
rect 86476 1408 86516 1448
rect 86668 1324 86708 1364
rect 87436 8464 87476 8504
rect 87340 7120 87380 7160
rect 87340 6952 87380 6992
rect 87532 8128 87572 8168
rect 87628 7792 87668 7832
rect 87532 7204 87572 7244
rect 87820 8296 87860 8336
rect 88012 8716 88052 8756
rect 88204 9472 88244 9512
rect 88684 10228 88724 10268
rect 88972 10144 89012 10184
rect 88588 9556 88628 9596
rect 88204 9220 88244 9260
rect 88108 8464 88148 8504
rect 88204 8296 88244 8336
rect 88204 8128 88244 8168
rect 87820 7708 87860 7748
rect 87724 7288 87764 7328
rect 87628 7120 87668 7160
rect 87436 6532 87476 6572
rect 88396 9220 88436 9260
rect 88396 8716 88436 8756
rect 88780 9220 88820 9260
rect 89068 10060 89108 10100
rect 89452 10144 89492 10184
rect 89068 9304 89108 9344
rect 89548 9220 89588 9260
rect 88972 9136 89012 9176
rect 88876 8800 88916 8840
rect 89068 8800 89108 8840
rect 88684 8128 88724 8168
rect 88396 7876 88436 7916
rect 88300 7792 88340 7832
rect 88204 7456 88244 7496
rect 88012 7036 88052 7076
rect 88204 7036 88244 7076
rect 88108 6952 88148 6992
rect 87436 6280 87476 6320
rect 87052 3592 87092 3632
rect 87244 3928 87284 3968
rect 87148 3508 87188 3548
rect 87436 4432 87476 4472
rect 87820 6196 87860 6236
rect 87724 4936 87764 4976
rect 88588 7876 88628 7916
rect 89164 8632 89204 8672
rect 89356 8716 89396 8756
rect 89548 8632 89588 8672
rect 92428 10228 92468 10268
rect 90028 9640 90068 9680
rect 89740 9220 89780 9260
rect 89836 9136 89876 9176
rect 89452 8296 89492 8336
rect 89260 8128 89300 8168
rect 88588 7540 88628 7580
rect 89452 7708 89492 7748
rect 88972 7624 89012 7664
rect 89164 7624 89204 7664
rect 88780 7456 88820 7496
rect 88684 7036 88724 7076
rect 88588 6700 88628 6740
rect 88108 4936 88148 4976
rect 88204 4852 88244 4892
rect 87052 3172 87092 3212
rect 86956 2500 86996 2540
rect 87436 3172 87476 3212
rect 86860 1576 86900 1616
rect 86860 1072 86900 1112
rect 86764 736 86804 776
rect 87244 1408 87284 1448
rect 87340 484 87380 524
rect 87820 3508 87860 3548
rect 87724 2668 87764 2708
rect 87628 2500 87668 2540
rect 88204 3928 88244 3968
rect 88108 2668 88148 2708
rect 88492 4936 88532 4976
rect 88396 4096 88436 4136
rect 89356 7540 89396 7580
rect 89068 5104 89108 5144
rect 88780 5020 88820 5060
rect 88684 4852 88724 4892
rect 88972 4684 89012 4724
rect 89644 6868 89684 6908
rect 89548 6280 89588 6320
rect 89740 5020 89780 5060
rect 89644 4768 89684 4808
rect 89740 4264 89780 4304
rect 89932 8212 89972 8252
rect 89932 4264 89972 4304
rect 89836 4096 89876 4136
rect 88012 1576 88052 1616
rect 87916 1324 87956 1364
rect 87820 1240 87860 1280
rect 87532 652 87572 692
rect 88108 988 88148 1028
rect 88396 1492 88436 1532
rect 88588 3424 88628 3464
rect 88588 3004 88628 3044
rect 88588 2668 88628 2708
rect 88588 1912 88628 1952
rect 88492 1408 88532 1448
rect 88396 1324 88436 1364
rect 88684 1240 88724 1280
rect 88876 2416 88916 2456
rect 88876 1660 88916 1700
rect 88972 1492 89012 1532
rect 88780 1072 88820 1112
rect 88780 64 88820 104
rect 89164 3172 89204 3212
rect 89068 1324 89108 1364
rect 89164 1240 89204 1280
rect 89356 2500 89396 2540
rect 89356 2332 89396 2372
rect 89260 148 89300 188
rect 89548 1576 89588 1616
rect 92044 8968 92084 9008
rect 90124 8380 90164 8420
rect 91948 7372 91988 7412
rect 90508 7036 90548 7076
rect 90892 6280 90932 6320
rect 91276 5020 91316 5060
rect 91948 4936 91988 4976
rect 91660 4096 91700 4136
rect 92332 5188 92372 5228
rect 90124 2080 90164 2120
rect 89932 1912 89972 1952
rect 89644 1240 89684 1280
rect 89836 1576 89876 1616
rect 90124 1576 90164 1616
rect 89932 1240 89972 1280
rect 90508 2248 90548 2288
rect 90796 3928 90836 3968
rect 90700 2332 90740 2372
rect 90316 1492 90356 1532
rect 90316 1324 90356 1364
rect 90892 2584 90932 2624
rect 90892 1660 90932 1700
rect 90508 1492 90548 1532
rect 90412 1240 90452 1280
rect 91468 3928 91508 3968
rect 91756 3928 91796 3968
rect 91180 3508 91220 3548
rect 91084 1744 91124 1784
rect 91660 3424 91700 3464
rect 91276 2752 91316 2792
rect 91276 1744 91316 1784
rect 90988 1324 91028 1364
rect 92236 3928 92276 3968
rect 91948 3760 91988 3800
rect 91852 3508 91892 3548
rect 91468 1576 91508 1616
rect 91660 1576 91700 1616
rect 91852 1492 91892 1532
rect 92044 3424 92084 3464
rect 93196 10060 93236 10100
rect 93100 5356 93140 5396
rect 94408 9808 94448 9848
rect 94490 9808 94530 9848
rect 94572 9808 94612 9848
rect 94654 9808 94694 9848
rect 94736 9808 94776 9848
rect 97228 9388 97268 9428
rect 95648 9052 95688 9092
rect 95730 9052 95770 9092
rect 95812 9052 95852 9092
rect 95894 9052 95934 9092
rect 95976 9052 96016 9092
rect 95788 8884 95828 8924
rect 94408 8296 94448 8336
rect 94490 8296 94530 8336
rect 94572 8296 94612 8336
rect 94654 8296 94694 8336
rect 94736 8296 94776 8336
rect 93964 8044 94004 8084
rect 93484 5944 93524 5984
rect 93292 4768 93332 4808
rect 93292 4096 93332 4136
rect 92620 3760 92660 3800
rect 92908 3760 92948 3800
rect 92236 1660 92276 1700
rect 92812 3088 92852 3128
rect 93100 3592 93140 3632
rect 92620 1744 92660 1784
rect 92428 1660 92468 1700
rect 92044 1492 92084 1532
rect 92812 1744 92852 1784
rect 93004 1576 93044 1616
rect 93388 3760 93428 3800
rect 93580 4516 93620 4556
rect 93868 4096 93908 4136
rect 94252 7960 94292 8000
rect 96652 7792 96692 7832
rect 95788 7708 95828 7748
rect 95648 7540 95688 7580
rect 95730 7540 95770 7580
rect 95812 7540 95852 7580
rect 95894 7540 95934 7580
rect 95976 7540 96016 7580
rect 95500 7120 95540 7160
rect 94408 6784 94448 6824
rect 94490 6784 94530 6824
rect 94572 6784 94612 6824
rect 94654 6784 94694 6824
rect 94736 6784 94776 6824
rect 94408 5272 94448 5312
rect 94490 5272 94530 5312
rect 94572 5272 94612 5312
rect 94654 5272 94694 5312
rect 94736 5272 94776 5312
rect 93772 3592 93812 3632
rect 94252 4012 94292 4052
rect 94060 3928 94100 3968
rect 93676 3340 93716 3380
rect 93196 3172 93236 3212
rect 93388 1492 93428 1532
rect 94156 3340 94196 3380
rect 93772 1660 93812 1700
rect 93580 1576 93620 1616
rect 94156 1744 94196 1784
rect 93964 1660 94004 1700
rect 95116 4096 95156 4136
rect 95648 6028 95688 6068
rect 95730 6028 95770 6068
rect 95812 6028 95852 6068
rect 95894 6028 95934 6068
rect 95976 6028 96016 6068
rect 96076 5776 96116 5816
rect 95648 4516 95688 4556
rect 95730 4516 95770 4556
rect 95812 4516 95852 4556
rect 95894 4516 95934 4556
rect 95976 4516 96016 4556
rect 96268 5692 96308 5732
rect 97036 7624 97076 7664
rect 97132 4936 97172 4976
rect 97900 9304 97940 9344
rect 97612 9136 97652 9176
rect 97420 8800 97460 8840
rect 97228 4096 97268 4136
rect 94924 4012 94964 4052
rect 97516 5608 97556 5648
rect 94540 3928 94580 3968
rect 94732 3928 94772 3968
rect 94408 3760 94448 3800
rect 94490 3760 94530 3800
rect 94572 3760 94612 3800
rect 94654 3760 94694 3800
rect 94736 3760 94776 3800
rect 94732 3424 94772 3464
rect 95116 3424 95156 3464
rect 94348 3256 94388 3296
rect 94540 3172 94580 3212
rect 96172 3928 96212 3968
rect 95596 3760 95636 3800
rect 96076 3760 96116 3800
rect 95500 3424 95540 3464
rect 94348 1492 94388 1532
rect 94732 1744 94772 1784
rect 95884 3424 95924 3464
rect 94924 1576 94964 1616
rect 95308 1660 95348 1700
rect 95116 1576 95156 1616
rect 95648 3004 95688 3044
rect 95730 3004 95770 3044
rect 95812 3004 95852 3044
rect 95894 3004 95934 3044
rect 95976 3004 96016 3044
rect 95692 2836 95732 2876
rect 95500 1492 95540 1532
rect 95500 1324 95540 1364
rect 96076 1744 96116 1784
rect 95884 1660 95924 1700
rect 96844 3928 96884 3968
rect 96652 3424 96692 3464
rect 96364 2836 96404 2876
rect 96268 2668 96308 2708
rect 96652 2500 96692 2540
rect 96460 1576 96500 1616
rect 96268 1492 96308 1532
rect 96460 1408 96500 1448
rect 97036 3172 97076 3212
rect 96940 2920 96980 2960
rect 96940 1996 96980 2036
rect 96844 1324 96884 1364
rect 97420 3592 97460 3632
rect 97420 3424 97460 3464
rect 97324 3340 97364 3380
rect 97228 1660 97268 1700
rect 98188 7708 98228 7748
rect 97708 4936 97748 4976
rect 97804 4264 97844 4304
rect 97132 1408 97172 1448
rect 97804 3424 97844 3464
rect 98092 4936 98132 4976
rect 98476 6448 98516 6488
rect 98284 4684 98324 4724
rect 98476 5440 98516 5480
rect 98476 4936 98516 4976
rect 98476 4684 98516 4724
rect 97996 3340 98036 3380
rect 98188 3676 98228 3716
rect 98092 3004 98132 3044
rect 97996 2584 98036 2624
rect 98380 3928 98420 3968
rect 98380 3172 98420 3212
rect 98380 3004 98420 3044
rect 97996 2332 98036 2372
rect 97708 1996 97748 2036
rect 97612 1492 97652 1532
rect 97612 1324 97652 1364
rect 98572 4096 98612 4136
rect 98572 3424 98612 3464
rect 98956 4264 98996 4304
rect 98764 3928 98804 3968
rect 98476 2332 98516 2372
rect 98860 3592 98900 3632
rect 98764 1324 98804 1364
<< metal3 >>
rect 6211 11908 6220 11948
rect 6260 11908 53164 11948
rect 53204 11908 53213 11948
rect 59683 11908 59692 11948
rect 59732 11908 93772 11948
rect 93812 11908 93821 11948
rect 28387 11404 28396 11444
rect 28436 11404 49900 11444
rect 49940 11404 49949 11444
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 18799 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 19185 11360
rect 33919 11320 33928 11360
rect 33968 11320 34010 11360
rect 34050 11320 34092 11360
rect 34132 11320 34174 11360
rect 34214 11320 34256 11360
rect 34296 11320 34305 11360
rect 49039 11320 49048 11360
rect 49088 11320 49130 11360
rect 49170 11320 49212 11360
rect 49252 11320 49294 11360
rect 49334 11320 49376 11360
rect 49416 11320 49425 11360
rect 64159 11320 64168 11360
rect 64208 11320 64250 11360
rect 64290 11320 64332 11360
rect 64372 11320 64414 11360
rect 64454 11320 64496 11360
rect 64536 11320 64545 11360
rect 79279 11320 79288 11360
rect 79328 11320 79370 11360
rect 79410 11320 79452 11360
rect 79492 11320 79534 11360
rect 79574 11320 79616 11360
rect 79656 11320 79665 11360
rect 94399 11320 94408 11360
rect 94448 11320 94490 11360
rect 94530 11320 94572 11360
rect 94612 11320 94654 11360
rect 94694 11320 94736 11360
rect 94776 11320 94785 11360
rect 19555 11068 19564 11108
rect 19604 11068 21196 11108
rect 21236 11068 21245 11108
rect 24355 11068 24364 11108
rect 24404 11068 25420 11108
rect 25460 11068 25469 11108
rect 30595 11068 30604 11108
rect 30644 11068 31372 11108
rect 31412 11068 31421 11108
rect 11971 10984 11980 11024
rect 12020 10984 19276 11024
rect 19316 10984 24460 11024
rect 24500 10984 30988 11024
rect 31028 10984 36172 11024
rect 36212 10984 36221 11024
rect 17443 10940 17501 10941
rect 12163 10900 12172 10940
rect 12212 10900 12748 10940
rect 12788 10900 15860 10940
rect 17358 10900 17452 10940
rect 17492 10900 17501 10940
rect 19939 10900 19948 10940
rect 19988 10900 24748 10940
rect 24788 10900 25228 10940
rect 25268 10900 25277 10940
rect 25411 10900 25420 10940
rect 25460 10900 30508 10940
rect 30548 10900 30557 10940
rect 30787 10900 30796 10940
rect 30836 10900 31180 10940
rect 31220 10900 31229 10940
rect 36067 10900 36076 10940
rect 36116 10900 40780 10940
rect 40820 10900 40829 10940
rect 61315 10900 61324 10940
rect 61364 10900 83116 10940
rect 83156 10900 83165 10940
rect 15820 10856 15860 10900
rect 17443 10899 17501 10900
rect 25228 10856 25268 10900
rect 10723 10816 10732 10856
rect 10772 10816 15724 10856
rect 15764 10816 15773 10856
rect 15820 10816 19564 10856
rect 19604 10816 19613 10856
rect 24067 10816 24076 10856
rect 24116 10816 24364 10856
rect 24404 10816 24413 10856
rect 25228 10816 30604 10856
rect 30644 10816 30653 10856
rect 30700 10816 31084 10856
rect 31124 10816 37036 10856
rect 37076 10816 37420 10856
rect 37460 10816 37820 10856
rect 37987 10816 37996 10856
rect 38036 10816 52108 10856
rect 52148 10816 52157 10856
rect 30700 10772 30740 10816
rect 37780 10772 37820 10816
rect 10819 10732 10828 10772
rect 10868 10732 11500 10772
rect 11540 10732 11788 10772
rect 11828 10732 14572 10772
rect 14612 10732 14621 10772
rect 15139 10732 15148 10772
rect 15188 10732 15628 10772
rect 15668 10732 18604 10772
rect 18644 10732 19660 10772
rect 19700 10732 21292 10772
rect 21332 10732 21341 10772
rect 21475 10732 21484 10772
rect 21524 10732 25132 10772
rect 25172 10732 30740 10772
rect 30796 10732 36652 10772
rect 36692 10732 36701 10772
rect 37780 10732 40588 10772
rect 40628 10732 40637 10772
rect 50275 10732 50284 10772
rect 50324 10732 51244 10772
rect 51284 10732 51293 10772
rect 30796 10688 30836 10732
rect 11587 10648 11596 10688
rect 11636 10648 12364 10688
rect 12404 10648 14956 10688
rect 14996 10648 15532 10688
rect 15572 10648 15581 10688
rect 19075 10648 19084 10688
rect 19124 10648 23404 10688
rect 23444 10648 23453 10688
rect 23875 10648 23884 10688
rect 23924 10648 29260 10688
rect 29300 10648 29309 10688
rect 30787 10648 30796 10688
rect 30836 10648 30845 10688
rect 30979 10648 30988 10688
rect 31028 10648 31372 10688
rect 31412 10648 31421 10688
rect 36451 10648 36460 10688
rect 36500 10648 41260 10688
rect 41300 10648 41309 10688
rect 48643 10648 48652 10688
rect 48692 10648 68428 10688
rect 68468 10648 68477 10688
rect 58531 10604 58589 10605
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 10915 10564 10924 10604
rect 10964 10564 14476 10604
rect 14516 10564 14525 10604
rect 14755 10564 14764 10604
rect 14804 10564 19948 10604
rect 19988 10564 19997 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 23779 10564 23788 10604
rect 23828 10564 31564 10604
rect 31604 10564 31613 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 36643 10564 36652 10604
rect 36692 10564 38092 10604
rect 38132 10564 38141 10604
rect 50279 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 50665 10604
rect 57667 10564 57676 10604
rect 57716 10564 58540 10604
rect 58580 10564 58589 10604
rect 65399 10564 65408 10604
rect 65448 10564 65490 10604
rect 65530 10564 65572 10604
rect 65612 10564 65654 10604
rect 65694 10564 65736 10604
rect 65776 10564 65785 10604
rect 80519 10564 80528 10604
rect 80568 10564 80610 10604
rect 80650 10564 80692 10604
rect 80732 10564 80774 10604
rect 80814 10564 80856 10604
rect 80896 10564 80905 10604
rect 95639 10564 95648 10604
rect 95688 10564 95730 10604
rect 95770 10564 95812 10604
rect 95852 10564 95894 10604
rect 95934 10564 95976 10604
rect 96016 10564 96025 10604
rect 58531 10563 58589 10564
rect 19843 10520 19901 10521
rect 11203 10480 11212 10520
rect 11252 10480 12364 10520
rect 12404 10480 19180 10520
rect 19220 10480 19229 10520
rect 19758 10480 19852 10520
rect 19892 10480 19901 10520
rect 19843 10479 19901 10480
rect 20140 10480 21676 10520
rect 21716 10480 25420 10520
rect 25460 10480 31948 10520
rect 31988 10480 31997 10520
rect 36163 10480 36172 10520
rect 36212 10480 37172 10520
rect 37315 10480 37324 10520
rect 37364 10480 38764 10520
rect 38804 10480 38813 10520
rect 38860 10480 52492 10520
rect 52532 10480 52541 10520
rect 53059 10480 53068 10520
rect 53108 10480 73804 10520
rect 73844 10480 73853 10520
rect 73987 10480 73996 10520
rect 74036 10480 77068 10520
rect 77108 10480 78028 10520
rect 78068 10480 78077 10520
rect 82819 10480 82828 10520
rect 82868 10480 84076 10520
rect 84116 10480 84125 10520
rect 88291 10480 88300 10520
rect 88340 10480 92812 10520
rect 92852 10480 92861 10520
rect 20140 10436 20180 10480
rect 37132 10436 37172 10480
rect 38860 10436 38900 10480
rect 12163 10396 12172 10436
rect 12212 10396 12556 10436
rect 12596 10396 12940 10436
rect 12980 10396 16300 10436
rect 16340 10396 18796 10436
rect 18836 10396 20180 10436
rect 21283 10396 21292 10436
rect 21332 10396 24844 10436
rect 24884 10396 30220 10436
rect 30260 10396 30269 10436
rect 30403 10396 30412 10436
rect 30452 10396 35596 10436
rect 35636 10396 37076 10436
rect 37132 10396 38380 10436
rect 38420 10396 38900 10436
rect 41539 10396 41548 10436
rect 41588 10396 49804 10436
rect 49844 10396 49853 10436
rect 50275 10396 50284 10436
rect 50324 10396 51148 10436
rect 51188 10396 55460 10436
rect 37036 10352 37076 10396
rect 15523 10312 15532 10352
rect 15572 10312 20332 10352
rect 20372 10312 21484 10352
rect 21524 10312 21533 10352
rect 28960 10312 31180 10352
rect 31220 10312 36940 10352
rect 36980 10312 36989 10352
rect 37036 10312 37996 10352
rect 38036 10312 38045 10352
rect 38755 10312 38764 10352
rect 38804 10312 49420 10352
rect 49460 10312 49469 10352
rect 12067 10268 12125 10269
rect 28960 10268 29000 10312
rect 35587 10268 35645 10269
rect 55420 10268 55460 10396
rect 57580 10396 58060 10436
rect 58100 10396 60076 10436
rect 60116 10396 60364 10436
rect 60404 10396 60413 10436
rect 69763 10396 69772 10436
rect 69812 10396 71308 10436
rect 71348 10396 77644 10436
rect 77684 10396 77693 10436
rect 82444 10396 87148 10436
rect 87188 10396 89644 10436
rect 89684 10396 89932 10436
rect 89972 10396 89981 10436
rect 57580 10352 57620 10396
rect 82444 10352 82484 10396
rect 56227 10312 56236 10352
rect 56276 10312 57580 10352
rect 57620 10312 57629 10352
rect 58147 10312 58156 10352
rect 58196 10312 58636 10352
rect 58676 10312 58828 10352
rect 58868 10312 58877 10352
rect 73123 10312 73132 10352
rect 73172 10312 76492 10352
rect 76532 10312 82444 10352
rect 82484 10312 82493 10352
rect 82540 10312 83212 10352
rect 83252 10312 89164 10352
rect 89204 10312 89213 10352
rect 82435 10268 82493 10269
rect 11395 10228 11404 10268
rect 11444 10228 11596 10268
rect 11636 10228 11645 10268
rect 11982 10228 12076 10268
rect 12116 10228 12125 10268
rect 14563 10228 14572 10268
rect 14612 10228 15340 10268
rect 15380 10228 15724 10268
rect 15764 10228 15773 10268
rect 15907 10228 15916 10268
rect 15956 10228 16108 10268
rect 16148 10228 19948 10268
rect 19988 10228 24748 10268
rect 24788 10228 29000 10268
rect 30307 10228 30316 10268
rect 30356 10228 30796 10268
rect 30836 10228 30845 10268
rect 31468 10228 35596 10268
rect 35636 10228 35645 10268
rect 35779 10228 35788 10268
rect 35828 10228 35980 10268
rect 36020 10228 36364 10268
rect 36404 10228 36748 10268
rect 36788 10228 36797 10268
rect 36844 10228 37324 10268
rect 37364 10228 37373 10268
rect 37603 10228 37612 10268
rect 37652 10228 37804 10268
rect 37844 10228 38188 10268
rect 38228 10228 38572 10268
rect 38612 10228 38956 10268
rect 38996 10228 39005 10268
rect 42787 10228 42796 10268
rect 42836 10228 48652 10268
rect 48692 10228 48701 10268
rect 55420 10228 69580 10268
rect 69620 10228 69629 10268
rect 73060 10228 73324 10268
rect 73364 10228 73373 10268
rect 73507 10228 73516 10268
rect 73556 10228 74476 10268
rect 74516 10228 77260 10268
rect 77300 10228 82444 10268
rect 82484 10228 82493 10268
rect 12067 10227 12125 10228
rect 31468 10184 31508 10228
rect 35587 10227 35645 10228
rect 36844 10184 36884 10228
rect 73060 10184 73100 10228
rect 82435 10227 82493 10228
rect 82540 10184 82580 10312
rect 82627 10268 82685 10269
rect 82627 10228 82636 10268
rect 82676 10228 83596 10268
rect 83636 10228 88012 10268
rect 88052 10228 88396 10268
rect 88436 10228 88445 10268
rect 88675 10228 88684 10268
rect 88724 10228 92428 10268
rect 92468 10228 92477 10268
rect 82627 10227 82685 10228
rect 7363 10144 7372 10184
rect 7412 10144 12844 10184
rect 12884 10144 12893 10184
rect 14467 10144 14476 10184
rect 14516 10144 17644 10184
rect 17684 10144 17693 10184
rect 19171 10144 19180 10184
rect 19220 10144 24404 10184
rect 16195 10100 16253 10101
rect 24364 10100 24404 10144
rect 30508 10144 31508 10184
rect 31555 10144 31564 10184
rect 31604 10144 36556 10184
rect 36596 10144 36884 10184
rect 36931 10144 36940 10184
rect 36980 10144 39148 10184
rect 39188 10144 40684 10184
rect 40724 10144 40733 10184
rect 55420 10144 73100 10184
rect 77443 10144 77452 10184
rect 77492 10144 77836 10184
rect 77876 10144 77885 10184
rect 78019 10144 78028 10184
rect 78068 10144 82580 10184
rect 82636 10144 83980 10184
rect 84020 10144 84029 10184
rect 88195 10144 88204 10184
rect 88244 10144 88972 10184
rect 89012 10144 89452 10184
rect 89492 10144 89501 10184
rect 11779 10060 11788 10100
rect 11828 10060 12748 10100
rect 12788 10060 12797 10100
rect 14851 10060 14860 10100
rect 14900 10060 15436 10100
rect 15476 10060 15485 10100
rect 16110 10060 16204 10100
rect 16244 10060 16253 10100
rect 18979 10060 18988 10100
rect 19028 10060 19372 10100
rect 19412 10060 19756 10100
rect 19796 10060 20131 10100
rect 20171 10060 20180 10100
rect 23971 10060 23980 10100
rect 24020 10060 24172 10100
rect 24212 10060 24221 10100
rect 24364 10060 30412 10100
rect 30452 10060 30461 10100
rect 16195 10059 16253 10060
rect 3427 9976 3436 10016
rect 3476 9976 22772 10016
rect 7459 9892 7468 9932
rect 7508 9892 21580 9932
rect 21620 9892 21629 9932
rect 15139 9848 15197 9849
rect 22732 9848 22772 9976
rect 24364 9932 24404 10060
rect 30508 10016 30548 10144
rect 37891 10100 37949 10101
rect 55420 10100 55460 10144
rect 60355 10100 60413 10101
rect 74371 10100 74429 10101
rect 82636 10100 82676 10144
rect 88579 10100 88637 10101
rect 30691 10060 30700 10100
rect 30740 10060 35884 10100
rect 35924 10060 35933 10100
rect 37806 10060 37900 10100
rect 37940 10060 37949 10100
rect 38083 10060 38092 10100
rect 38132 10060 38380 10100
rect 38420 10060 41836 10100
rect 41876 10060 41885 10100
rect 53443 10060 53452 10100
rect 53492 10060 55460 10100
rect 57283 10060 57292 10100
rect 57332 10060 58444 10100
rect 58484 10060 58493 10100
rect 58627 10060 58636 10100
rect 58676 10060 59020 10100
rect 59060 10060 59069 10100
rect 60067 10060 60076 10100
rect 60116 10060 60364 10100
rect 60404 10060 60413 10100
rect 69091 10060 69100 10100
rect 69140 10060 73132 10100
rect 73172 10060 73181 10100
rect 74286 10060 74380 10100
rect 74420 10060 74429 10100
rect 77635 10060 77644 10100
rect 77684 10060 82676 10100
rect 82723 10060 82732 10100
rect 82772 10060 83404 10100
rect 83444 10060 83788 10100
rect 83828 10060 84172 10100
rect 84212 10060 84221 10100
rect 87907 10060 87916 10100
rect 87956 10060 88588 10100
rect 88628 10060 88637 10100
rect 89059 10060 89068 10100
rect 89108 10060 93196 10100
rect 93236 10060 93245 10100
rect 37891 10059 37949 10060
rect 60355 10059 60413 10060
rect 74371 10059 74429 10060
rect 88579 10059 88637 10060
rect 32035 10016 32093 10017
rect 38659 10016 38717 10017
rect 75619 10016 75677 10017
rect 30316 9976 30548 10016
rect 30595 9976 30604 10016
rect 30644 9976 30988 10016
rect 31028 9976 31372 10016
rect 31412 9976 31421 10016
rect 31950 9976 32044 10016
rect 32084 9976 32093 10016
rect 35683 9976 35692 10016
rect 35732 9976 38668 10016
rect 38708 9976 38717 10016
rect 72931 9976 72940 10016
rect 72980 9976 73228 10016
rect 73268 9976 73277 10016
rect 75619 9976 75628 10016
rect 75668 9976 77356 10016
rect 77396 9976 77405 10016
rect 83299 9976 83308 10016
rect 83348 9976 83884 10016
rect 83924 9976 83933 10016
rect 30316 9932 30356 9976
rect 32035 9975 32093 9976
rect 38659 9975 38717 9976
rect 75619 9975 75677 9976
rect 24355 9892 24364 9932
rect 24404 9892 24413 9932
rect 30307 9892 30316 9932
rect 30356 9892 30365 9932
rect 34531 9892 34540 9932
rect 34580 9892 40204 9932
rect 40244 9892 40253 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 15054 9808 15148 9848
rect 15188 9808 15197 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 22732 9808 25324 9848
rect 25364 9808 25373 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 36643 9808 36652 9848
rect 36692 9808 40012 9848
rect 40052 9808 40061 9848
rect 49039 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49425 9848
rect 64159 9808 64168 9848
rect 64208 9808 64250 9848
rect 64290 9808 64332 9848
rect 64372 9808 64414 9848
rect 64454 9808 64496 9848
rect 64536 9808 64545 9848
rect 79279 9808 79288 9848
rect 79328 9808 79370 9848
rect 79410 9808 79452 9848
rect 79492 9808 79534 9848
rect 79574 9808 79616 9848
rect 79656 9808 79665 9848
rect 94399 9808 94408 9848
rect 94448 9808 94490 9848
rect 94530 9808 94572 9848
rect 94612 9808 94654 9848
rect 94694 9808 94736 9848
rect 94776 9808 94785 9848
rect 15139 9807 15197 9808
rect 19555 9724 19564 9764
rect 19604 9724 23788 9764
rect 23828 9724 23837 9764
rect 30883 9724 30892 9764
rect 30932 9724 36844 9764
rect 36884 9724 36893 9764
rect 37780 9724 42316 9764
rect 42356 9724 42365 9764
rect 46243 9724 46252 9764
rect 46292 9724 60460 9764
rect 60500 9724 60509 9764
rect 72163 9724 72172 9764
rect 72212 9724 77932 9764
rect 77972 9724 80620 9764
rect 80660 9724 88108 9764
rect 88148 9724 88157 9764
rect 37780 9680 37820 9724
rect 69475 9680 69533 9681
rect 15139 9640 15148 9680
rect 15188 9640 16300 9680
rect 16340 9640 19180 9680
rect 19220 9640 24076 9680
rect 24116 9640 24125 9680
rect 35107 9640 35116 9680
rect 35156 9640 37820 9680
rect 37891 9640 37900 9680
rect 37940 9640 43660 9680
rect 43700 9640 43709 9680
rect 56611 9640 56620 9680
rect 56660 9640 58636 9680
rect 58676 9640 59404 9680
rect 59444 9640 59884 9680
rect 59924 9640 59933 9680
rect 69475 9640 69484 9680
rect 69524 9640 73804 9680
rect 73844 9640 73853 9680
rect 74179 9640 74188 9680
rect 74228 9640 77452 9680
rect 77492 9640 77501 9680
rect 83203 9640 83212 9680
rect 83252 9640 90028 9680
rect 90068 9640 90077 9680
rect 69475 9639 69533 9640
rect 75235 9596 75293 9597
rect 11395 9556 11404 9596
rect 11444 9556 11692 9596
rect 11732 9556 11741 9596
rect 24259 9556 24268 9596
rect 24308 9556 27724 9596
rect 27764 9556 27773 9596
rect 30499 9556 30508 9596
rect 30548 9556 30557 9596
rect 30892 9556 31084 9596
rect 31124 9556 31133 9596
rect 36355 9556 36364 9596
rect 36404 9556 43084 9596
rect 43124 9556 43133 9596
rect 48451 9556 48460 9596
rect 48500 9556 48940 9596
rect 48980 9556 52108 9596
rect 52148 9556 52157 9596
rect 52291 9556 52300 9596
rect 52340 9556 53068 9596
rect 53108 9556 53117 9596
rect 55843 9556 55852 9596
rect 55892 9556 58732 9596
rect 58772 9556 59212 9596
rect 59252 9556 60844 9596
rect 60884 9556 60893 9596
rect 67939 9556 67948 9596
rect 67988 9556 72076 9596
rect 72116 9556 72125 9596
rect 75235 9556 75244 9596
rect 75284 9556 77740 9596
rect 77780 9556 77789 9596
rect 81859 9556 81868 9596
rect 81908 9556 87532 9596
rect 87572 9556 87581 9596
rect 88579 9556 88588 9596
rect 88628 9556 88637 9596
rect 6211 9472 6220 9512
rect 6260 9472 18700 9512
rect 18740 9472 18749 9512
rect 19459 9472 19468 9512
rect 19508 9472 21964 9512
rect 22004 9472 22013 9512
rect 24643 9472 24652 9512
rect 24692 9472 29644 9512
rect 29684 9472 29693 9512
rect 30508 9428 30548 9556
rect 30892 9512 30932 9556
rect 75235 9555 75293 9556
rect 88588 9512 88628 9556
rect 30883 9472 30892 9512
rect 30932 9472 30941 9512
rect 32236 9472 36460 9512
rect 36500 9472 37460 9512
rect 37507 9472 37516 9512
rect 37556 9472 47596 9512
rect 47636 9472 47645 9512
rect 49795 9472 49804 9512
rect 49844 9472 64280 9512
rect 66883 9472 66892 9512
rect 66932 9472 73036 9512
rect 73076 9472 73085 9512
rect 73219 9472 73228 9512
rect 73268 9472 73708 9512
rect 73748 9472 74284 9512
rect 74324 9472 74333 9512
rect 81004 9472 82060 9512
rect 82100 9472 82732 9512
rect 82772 9472 82781 9512
rect 83971 9472 83980 9512
rect 84020 9472 87916 9512
rect 87956 9472 88204 9512
rect 88244 9472 88628 9512
rect 32236 9428 32276 9472
rect 37420 9428 37460 9472
rect 64240 9428 64280 9472
rect 81004 9428 81044 9472
rect 9187 9388 9196 9428
rect 9236 9388 14668 9428
rect 14708 9388 14717 9428
rect 15907 9388 15916 9428
rect 15956 9388 16108 9428
rect 16148 9388 16157 9428
rect 18979 9388 18988 9428
rect 19028 9388 19372 9428
rect 19412 9388 19948 9428
rect 19988 9388 20620 9428
rect 20660 9388 20669 9428
rect 24163 9388 24172 9428
rect 24212 9388 24556 9428
rect 24596 9388 25228 9428
rect 25268 9388 25277 9428
rect 30508 9388 30796 9428
rect 30836 9388 32236 9428
rect 32276 9388 32285 9428
rect 36259 9388 36268 9428
rect 36308 9388 36652 9428
rect 36692 9388 37324 9428
rect 37364 9388 37373 9428
rect 37420 9388 37900 9428
rect 37940 9388 38188 9428
rect 38228 9388 38237 9428
rect 38284 9388 38956 9428
rect 38996 9388 39340 9428
rect 39380 9388 39389 9428
rect 41560 9388 49652 9428
rect 51427 9388 51436 9428
rect 51476 9388 51820 9428
rect 51860 9388 52012 9428
rect 52052 9388 52061 9428
rect 54787 9388 54796 9428
rect 54836 9388 55660 9428
rect 55700 9388 56140 9428
rect 56180 9388 56189 9428
rect 58147 9388 58156 9428
rect 58196 9388 59116 9428
rect 59156 9388 59165 9428
rect 59587 9388 59596 9428
rect 59636 9388 59884 9428
rect 59924 9388 59933 9428
rect 60355 9388 60364 9428
rect 60404 9388 60844 9428
rect 60884 9388 60893 9428
rect 64240 9388 65164 9428
rect 65204 9388 65213 9428
rect 70723 9388 70732 9428
rect 70772 9388 71788 9428
rect 71828 9388 76972 9428
rect 77012 9388 77021 9428
rect 80227 9388 80236 9428
rect 80276 9388 80812 9428
rect 80852 9388 81004 9428
rect 81044 9388 81053 9428
rect 81196 9388 86860 9428
rect 86900 9388 86909 9428
rect 87811 9388 87820 9428
rect 87860 9388 97228 9428
rect 97268 9388 97277 9428
rect 38284 9344 38324 9388
rect 41560 9344 41600 9388
rect 45283 9344 45341 9345
rect 9571 9304 9580 9344
rect 9620 9304 15436 9344
rect 15476 9304 15485 9344
rect 19459 9304 19468 9344
rect 19508 9304 23500 9344
rect 23540 9304 23549 9344
rect 24259 9304 24268 9344
rect 24308 9304 28108 9344
rect 28148 9304 28157 9344
rect 34915 9304 34924 9344
rect 34964 9304 36404 9344
rect 36835 9304 36844 9344
rect 36884 9304 38324 9344
rect 38467 9304 38476 9344
rect 38516 9304 38525 9344
rect 40291 9304 40300 9344
rect 40340 9304 41600 9344
rect 43267 9304 43276 9344
rect 43316 9304 45292 9344
rect 45332 9304 45341 9344
rect 9763 9220 9772 9260
rect 9812 9220 13036 9260
rect 13076 9220 13085 9260
rect 30595 9220 30604 9260
rect 30644 9220 30988 9260
rect 31028 9220 31037 9260
rect 34819 9220 34828 9260
rect 34868 9220 35116 9260
rect 35156 9220 35165 9260
rect 36364 9176 36404 9304
rect 38476 9260 38516 9304
rect 45283 9303 45341 9304
rect 49612 9260 49652 9388
rect 52012 9344 52052 9388
rect 76972 9344 77012 9388
rect 81196 9344 81236 9388
rect 52012 9304 52396 9344
rect 52436 9304 55948 9344
rect 55988 9304 56332 9344
rect 56372 9304 56716 9344
rect 56756 9304 56765 9344
rect 71587 9304 71596 9344
rect 71636 9304 71980 9344
rect 72020 9304 72940 9344
rect 72980 9304 72989 9344
rect 76972 9304 81196 9344
rect 81236 9304 81245 9344
rect 81475 9304 81484 9344
rect 81524 9304 86764 9344
rect 86804 9304 86813 9344
rect 87043 9304 87052 9344
rect 87092 9304 87724 9344
rect 87764 9304 87773 9344
rect 89059 9304 89068 9344
rect 89108 9304 97900 9344
rect 97940 9304 97949 9344
rect 36931 9220 36940 9260
rect 36980 9220 37804 9260
rect 37844 9220 37853 9260
rect 37987 9220 37996 9260
rect 38036 9220 38380 9260
rect 38420 9220 38429 9260
rect 38476 9220 47020 9260
rect 47060 9220 47069 9260
rect 49603 9220 49612 9260
rect 49652 9220 49661 9260
rect 51427 9220 51436 9260
rect 51476 9220 52012 9260
rect 52052 9220 52588 9260
rect 52628 9220 52637 9260
rect 63715 9220 63724 9260
rect 63764 9220 70060 9260
rect 70100 9220 70109 9260
rect 76675 9220 76684 9260
rect 76724 9220 77164 9260
rect 77204 9220 77548 9260
rect 77588 9220 77597 9260
rect 81667 9220 81676 9260
rect 81716 9220 85996 9260
rect 86036 9220 86045 9260
rect 87724 9176 87764 9304
rect 88195 9220 88204 9260
rect 88244 9220 88396 9260
rect 88436 9220 88780 9260
rect 88820 9220 89548 9260
rect 89588 9220 89597 9260
rect 89731 9220 89740 9260
rect 89780 9220 89789 9260
rect 89740 9176 89780 9220
rect 11683 9136 11692 9176
rect 11732 9136 14476 9176
rect 14516 9136 14525 9176
rect 28675 9136 28684 9176
rect 28724 9136 33388 9176
rect 33428 9136 33437 9176
rect 36364 9136 38036 9176
rect 38083 9136 38092 9176
rect 38132 9136 42700 9176
rect 42740 9136 42749 9176
rect 46600 9136 48172 9176
rect 48212 9136 70540 9176
rect 70580 9136 70589 9176
rect 71203 9136 71212 9176
rect 71252 9136 75436 9176
rect 75476 9136 75485 9176
rect 77356 9136 81868 9176
rect 81908 9136 81917 9176
rect 87724 9136 88972 9176
rect 89012 9136 89780 9176
rect 89827 9136 89836 9176
rect 89876 9136 97612 9176
rect 97652 9136 97661 9176
rect 24451 9092 24509 9093
rect 37996 9092 38036 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 7180 9052 12364 9092
rect 12404 9052 12413 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 24366 9052 24460 9092
rect 24500 9052 24509 9092
rect 7180 8840 7220 9052
rect 24451 9051 24509 9052
rect 24940 9052 25324 9092
rect 25364 9052 25373 9092
rect 30691 9052 30700 9092
rect 30740 9052 35060 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37996 9052 38572 9092
rect 38612 9052 38621 9092
rect 38851 9052 38860 9092
rect 38900 9052 43756 9092
rect 43796 9052 43805 9092
rect 24940 9008 24980 9052
rect 26371 9008 26429 9009
rect 35020 9008 35060 9052
rect 46600 9008 46640 9136
rect 77356 9092 77396 9136
rect 78403 9092 78461 9093
rect 82243 9092 82301 9093
rect 89347 9092 89405 9093
rect 50279 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50665 9092
rect 55459 9052 55468 9092
rect 55508 9052 59596 9092
rect 59636 9052 59645 9092
rect 59875 9052 59884 9092
rect 59924 9052 60172 9092
rect 60212 9052 60364 9092
rect 60404 9052 60413 9092
rect 65399 9052 65408 9092
rect 65448 9052 65490 9092
rect 65530 9052 65572 9092
rect 65612 9052 65654 9092
rect 65694 9052 65736 9092
rect 65776 9052 65785 9092
rect 66115 9052 66124 9092
rect 66164 9052 73324 9092
rect 73364 9052 77356 9092
rect 77396 9052 77405 9092
rect 78318 9052 78412 9092
rect 78452 9052 78461 9092
rect 80519 9052 80528 9092
rect 80568 9052 80610 9092
rect 80650 9052 80692 9092
rect 80732 9052 80774 9092
rect 80814 9052 80856 9092
rect 80896 9052 80905 9092
rect 81091 9052 81100 9092
rect 81140 9052 82252 9092
rect 82292 9052 82301 9092
rect 83587 9052 83596 9092
rect 83636 9052 89356 9092
rect 89396 9052 89405 9092
rect 95639 9052 95648 9092
rect 95688 9052 95730 9092
rect 95770 9052 95812 9092
rect 95852 9052 95894 9092
rect 95934 9052 95976 9092
rect 96016 9052 96025 9092
rect 78403 9051 78461 9052
rect 82243 9051 82301 9052
rect 89347 9051 89405 9052
rect 7555 8968 7564 9008
rect 7604 8968 11980 9008
rect 12020 8968 12029 9008
rect 18403 8968 18412 9008
rect 18452 8968 24980 9008
rect 25027 8968 25036 9008
rect 25076 8968 26380 9008
rect 26420 8968 26429 9008
rect 31075 8968 31084 9008
rect 31124 8968 33484 9008
rect 33524 8968 33533 9008
rect 35020 8968 36844 9008
rect 36884 8968 36893 9008
rect 38371 8968 38380 9008
rect 38420 8968 38764 9008
rect 38804 8968 38813 9008
rect 41539 8968 41548 9008
rect 41588 8968 46640 9008
rect 48835 8968 48844 9008
rect 48884 8968 49324 9008
rect 49364 8968 49373 9008
rect 49603 8968 49612 9008
rect 49652 8968 62092 9008
rect 62132 8968 62141 9008
rect 62947 8968 62956 9008
rect 62996 8968 72172 9008
rect 72212 8968 72221 9008
rect 72931 8968 72940 9008
rect 72980 8968 74668 9008
rect 74708 8968 74717 9008
rect 82051 8968 82060 9008
rect 82100 8968 86092 9008
rect 86132 8968 86141 9008
rect 87715 8968 87724 9008
rect 87764 8968 92044 9008
rect 92084 8968 92093 9008
rect 26371 8967 26429 8968
rect 24931 8924 24989 8925
rect 81091 8924 81149 8925
rect 81571 8924 81629 8925
rect 11299 8884 11308 8924
rect 11348 8884 11788 8924
rect 11828 8884 11837 8924
rect 12451 8884 12460 8924
rect 12500 8884 15532 8924
rect 15572 8884 15581 8924
rect 24846 8884 24940 8924
rect 24980 8884 24989 8924
rect 28291 8884 28300 8924
rect 28340 8884 32620 8924
rect 32660 8884 32669 8924
rect 34819 8884 34828 8924
rect 34868 8884 37996 8924
rect 38036 8884 38045 8924
rect 46600 8884 68716 8924
rect 68756 8884 68765 8924
rect 73027 8884 73036 8924
rect 73076 8884 73100 8924
rect 73699 8884 73708 8924
rect 73748 8884 76588 8924
rect 76628 8884 76637 8924
rect 78211 8884 78220 8924
rect 78260 8884 78932 8924
rect 24931 8883 24989 8884
rect 12547 8840 12605 8841
rect 22147 8840 22205 8841
rect 31651 8840 31709 8841
rect 46600 8840 46640 8884
rect 73060 8841 73100 8884
rect 55075 8840 55133 8841
rect 56803 8840 56861 8841
rect 59683 8840 59741 8841
rect 70531 8840 70589 8841
rect 73027 8840 73100 8841
rect 75043 8840 75101 8841
rect 78892 8840 78932 8884
rect 80716 8884 81100 8924
rect 81140 8884 81149 8924
rect 81283 8884 81292 8924
rect 81332 8884 81580 8924
rect 81620 8884 81629 8924
rect 3043 8800 3052 8840
rect 3092 8800 7220 8840
rect 8803 8800 8812 8840
rect 8852 8800 11596 8840
rect 11636 8800 11645 8840
rect 12462 8800 12556 8840
rect 12596 8800 12605 8840
rect 14563 8800 14572 8840
rect 14612 8800 14956 8840
rect 14996 8800 15436 8840
rect 15476 8800 16300 8840
rect 16340 8800 16349 8840
rect 16771 8800 16780 8840
rect 16820 8800 18700 8840
rect 18740 8800 18749 8840
rect 19075 8800 19084 8840
rect 19124 8800 22156 8840
rect 22196 8800 22205 8840
rect 25027 8800 25036 8840
rect 25076 8800 26860 8840
rect 26900 8800 26909 8840
rect 27907 8800 27916 8840
rect 27956 8800 31660 8840
rect 31700 8800 31709 8840
rect 12547 8799 12605 8800
rect 22147 8799 22205 8800
rect 31651 8799 31709 8800
rect 31756 8800 35692 8840
rect 35732 8800 35741 8840
rect 44131 8800 44140 8840
rect 44180 8800 44908 8840
rect 44948 8800 46640 8840
rect 48451 8800 48460 8840
rect 48500 8800 49420 8840
rect 49460 8800 49708 8840
rect 49748 8800 49757 8840
rect 54986 8800 54995 8840
rect 55035 8800 55084 8840
rect 55124 8800 55133 8840
rect 56718 8800 56812 8840
rect 56852 8800 56861 8840
rect 57187 8800 57196 8840
rect 57236 8800 57245 8840
rect 59598 8800 59692 8840
rect 59732 8800 59741 8840
rect 60451 8800 60460 8840
rect 60500 8800 64012 8840
rect 64052 8800 64061 8840
rect 70531 8800 70540 8840
rect 70580 8800 70924 8840
rect 70964 8800 70973 8840
rect 73020 8800 73036 8840
rect 73076 8800 73100 8840
rect 74958 8800 75052 8840
rect 75092 8800 75101 8840
rect 76003 8800 76012 8840
rect 76052 8800 78796 8840
rect 78836 8800 78845 8840
rect 78892 8800 78988 8840
rect 79028 8800 79400 8840
rect 8995 8756 9053 8757
rect 15139 8756 15197 8757
rect 6115 8716 6124 8756
rect 6164 8716 9004 8756
rect 9044 8716 9053 8756
rect 9667 8716 9676 8756
rect 9716 8716 10060 8756
rect 10100 8716 10109 8756
rect 10627 8716 10636 8756
rect 10676 8716 11116 8756
rect 11156 8716 11500 8756
rect 11540 8716 11884 8756
rect 11924 8716 12268 8756
rect 12308 8716 12317 8756
rect 12451 8716 12460 8756
rect 12500 8716 12652 8756
rect 12692 8716 13324 8756
rect 13364 8716 13373 8756
rect 15139 8716 15148 8756
rect 15188 8716 15244 8756
rect 15284 8716 15293 8756
rect 18595 8716 18604 8756
rect 18644 8716 24076 8756
rect 24116 8716 24125 8756
rect 24355 8716 24364 8756
rect 24404 8716 24556 8756
rect 24596 8716 24940 8756
rect 24980 8716 25420 8756
rect 25460 8716 25469 8756
rect 27619 8716 27628 8756
rect 27668 8716 27820 8756
rect 27860 8716 28204 8756
rect 28244 8716 28588 8756
rect 28628 8716 29356 8756
rect 29396 8716 29405 8756
rect 29539 8716 29548 8756
rect 29588 8716 30028 8756
rect 30068 8716 30220 8756
rect 30260 8716 30269 8756
rect 8995 8715 9053 8716
rect 15139 8715 15197 8716
rect 31756 8672 31796 8800
rect 55075 8799 55133 8800
rect 56803 8799 56861 8800
rect 33763 8756 33821 8757
rect 49987 8756 50045 8757
rect 55084 8756 55124 8799
rect 57196 8756 57236 8800
rect 59683 8799 59741 8800
rect 70531 8799 70589 8800
rect 73027 8799 73085 8800
rect 75043 8799 75101 8800
rect 66979 8756 67037 8757
rect 79360 8756 79400 8800
rect 80716 8756 80756 8884
rect 81091 8883 81149 8884
rect 81571 8883 81629 8884
rect 81859 8924 81917 8925
rect 81859 8884 81868 8924
rect 81908 8884 85036 8924
rect 85076 8884 85085 8924
rect 86947 8884 86956 8924
rect 86996 8884 95788 8924
rect 95828 8884 95837 8924
rect 81859 8883 81917 8884
rect 82051 8840 82109 8841
rect 88867 8840 88925 8841
rect 80899 8800 80908 8840
rect 80948 8800 81484 8840
rect 81524 8800 81533 8840
rect 82020 8800 82060 8840
rect 82100 8800 82109 8840
rect 82339 8800 82348 8840
rect 82388 8800 83980 8840
rect 84020 8800 84029 8840
rect 87427 8800 87436 8840
rect 87476 8800 87916 8840
rect 87956 8800 88220 8840
rect 88836 8800 88876 8840
rect 88916 8800 88925 8840
rect 89059 8800 89068 8840
rect 89108 8800 97420 8840
rect 97460 8800 97469 8840
rect 82051 8799 82109 8800
rect 82060 8756 82100 8799
rect 88180 8756 88220 8800
rect 88867 8799 88925 8800
rect 88876 8756 88916 8799
rect 33763 8716 33772 8756
rect 33812 8716 34156 8756
rect 34196 8716 34205 8756
rect 34339 8716 34348 8756
rect 34388 8716 34732 8756
rect 34772 8716 35116 8756
rect 35156 8716 35500 8756
rect 35540 8716 37036 8756
rect 37076 8716 37085 8756
rect 37315 8716 37324 8756
rect 37364 8716 40588 8756
rect 40628 8716 40637 8756
rect 43363 8716 43372 8756
rect 43412 8716 46252 8756
rect 46292 8716 46301 8756
rect 48355 8716 48364 8756
rect 48404 8716 48748 8756
rect 48788 8716 48797 8756
rect 49902 8716 49996 8756
rect 50036 8716 50045 8756
rect 52867 8716 52876 8756
rect 52916 8716 53452 8756
rect 53492 8716 53501 8756
rect 54892 8716 54910 8756
rect 54950 8716 54972 8756
rect 55084 8716 55948 8756
rect 55988 8716 55997 8756
rect 57196 8716 57676 8756
rect 57716 8716 57725 8756
rect 58915 8716 58924 8756
rect 58964 8716 60076 8756
rect 60116 8716 60844 8756
rect 60884 8716 60893 8756
rect 66894 8716 66988 8756
rect 67028 8716 67037 8756
rect 67171 8716 67180 8756
rect 67220 8716 70156 8756
rect 70196 8716 74708 8756
rect 74755 8716 74764 8756
rect 74804 8716 75148 8756
rect 75188 8716 75532 8756
rect 75572 8716 75581 8756
rect 77923 8716 77932 8756
rect 77972 8716 78220 8756
rect 78260 8716 78892 8756
rect 78932 8716 78941 8756
rect 79360 8716 80756 8756
rect 80803 8716 80812 8756
rect 80852 8716 81196 8756
rect 81236 8716 81580 8756
rect 81620 8716 81964 8756
rect 82004 8716 82013 8756
rect 82060 8716 82156 8756
rect 82196 8716 83692 8756
rect 83732 8716 84364 8756
rect 84404 8716 84413 8756
rect 86851 8716 86860 8756
rect 86900 8716 87628 8756
rect 87668 8716 88012 8756
rect 88052 8716 88061 8756
rect 88180 8716 88396 8756
rect 88436 8716 88445 8756
rect 88876 8716 89356 8756
rect 89396 8716 89405 8756
rect 33763 8715 33821 8716
rect 49987 8715 50045 8716
rect 35203 8672 35261 8673
rect 54892 8672 54932 8716
rect 66979 8715 67037 8716
rect 54979 8672 55037 8673
rect 56803 8672 56861 8673
rect 74668 8672 74708 8716
rect 83683 8672 83741 8673
rect 11320 8632 13708 8672
rect 13748 8632 13757 8672
rect 18787 8632 18796 8672
rect 18836 8632 19372 8672
rect 19412 8632 19421 8672
rect 24739 8632 24748 8672
rect 24788 8632 28396 8672
rect 28436 8632 28445 8672
rect 28675 8632 28684 8672
rect 28724 8632 31756 8672
rect 31796 8632 31805 8672
rect 33667 8632 33676 8672
rect 33716 8632 35212 8672
rect 35252 8632 35308 8672
rect 35348 8632 35357 8672
rect 35683 8632 35692 8672
rect 35732 8632 42508 8672
rect 42548 8632 42557 8672
rect 47107 8632 47116 8672
rect 47156 8632 48268 8672
rect 48308 8632 48317 8672
rect 48931 8632 48940 8672
rect 48980 8632 52396 8672
rect 52436 8632 52684 8672
rect 52724 8632 52733 8672
rect 54307 8632 54316 8672
rect 54356 8632 54988 8672
rect 55028 8632 56812 8672
rect 56852 8632 56861 8672
rect 64963 8632 64972 8672
rect 65012 8632 70636 8672
rect 70676 8632 74612 8672
rect 74668 8632 75340 8672
rect 75380 8632 78700 8672
rect 78740 8632 81388 8672
rect 81428 8632 81920 8672
rect 83011 8632 83020 8672
rect 83060 8632 83500 8672
rect 83540 8632 83549 8672
rect 83683 8632 83692 8672
rect 83732 8632 84268 8672
rect 84308 8632 84317 8672
rect 87235 8632 87244 8672
rect 87284 8632 87532 8672
rect 87572 8632 89164 8672
rect 89204 8632 89548 8672
rect 89588 8632 89597 8672
rect 11320 8588 11360 8632
rect 11299 8548 11308 8588
rect 11348 8548 11360 8588
rect 14371 8548 14380 8588
rect 14420 8548 15724 8588
rect 15764 8548 22348 8588
rect 22388 8548 22397 8588
rect 24748 8504 24788 8632
rect 28099 8588 28157 8589
rect 28014 8548 28108 8588
rect 28148 8548 28157 8588
rect 28396 8588 28436 8632
rect 35203 8631 35261 8632
rect 54979 8631 55037 8632
rect 56803 8631 56861 8632
rect 49507 8588 49565 8589
rect 55843 8588 55901 8589
rect 71011 8588 71069 8589
rect 74572 8588 74612 8632
rect 81880 8588 81920 8632
rect 83683 8631 83741 8632
rect 28396 8548 32524 8588
rect 32564 8548 34540 8588
rect 34580 8548 39916 8588
rect 39956 8548 39965 8588
rect 44899 8548 44908 8588
rect 44948 8548 45196 8588
rect 45236 8548 45245 8588
rect 46531 8548 46540 8588
rect 46580 8548 48076 8588
rect 48116 8548 49516 8588
rect 49556 8548 55852 8588
rect 55892 8548 55988 8588
rect 56035 8548 56044 8588
rect 56084 8548 56428 8588
rect 56468 8548 56716 8588
rect 56756 8548 57004 8588
rect 57044 8548 57196 8588
rect 57236 8548 57245 8588
rect 60556 8548 61228 8588
rect 61268 8548 61277 8588
rect 70926 8548 71020 8588
rect 71060 8548 71069 8588
rect 74563 8548 74572 8588
rect 74612 8548 78507 8588
rect 78547 8548 81772 8588
rect 81812 8548 81821 8588
rect 81880 8548 82444 8588
rect 82484 8548 82493 8588
rect 28099 8547 28157 8548
rect 49507 8547 49565 8548
rect 55843 8547 55901 8548
rect 55948 8504 55988 8548
rect 19555 8464 19564 8504
rect 19604 8464 24788 8504
rect 25603 8464 25612 8504
rect 25652 8464 34060 8504
rect 34100 8464 34109 8504
rect 35587 8464 35596 8504
rect 35636 8464 37324 8504
rect 37364 8464 37373 8504
rect 37780 8464 39764 8504
rect 40867 8464 40876 8504
rect 40916 8464 46924 8504
rect 46964 8464 46973 8504
rect 53827 8464 53836 8504
rect 53876 8464 54700 8504
rect 54740 8464 54749 8504
rect 55948 8464 56140 8504
rect 56180 8464 56189 8504
rect 57379 8464 57388 8504
rect 57428 8464 59308 8504
rect 59348 8464 59357 8504
rect 35203 8420 35261 8421
rect 37780 8420 37820 8464
rect 39724 8420 39764 8464
rect 60556 8420 60596 8548
rect 71011 8547 71069 8548
rect 78787 8504 78845 8505
rect 73060 8464 75148 8504
rect 75188 8464 75197 8504
rect 76771 8464 76780 8504
rect 76820 8464 77164 8504
rect 77204 8464 77213 8504
rect 78403 8464 78412 8504
rect 78452 8464 78796 8504
rect 78836 8464 78845 8504
rect 80899 8464 80908 8504
rect 80948 8464 84268 8504
rect 84308 8464 85132 8504
rect 85172 8464 85181 8504
rect 87427 8464 87436 8504
rect 87476 8464 88108 8504
rect 88148 8464 88157 8504
rect 73060 8420 73100 8464
rect 78787 8463 78845 8464
rect 83779 8420 83837 8421
rect 11011 8380 11020 8420
rect 11060 8380 18604 8420
rect 18644 8380 18653 8420
rect 19267 8380 19276 8420
rect 19316 8380 24172 8420
rect 24212 8380 27436 8420
rect 27476 8380 29000 8420
rect 32131 8380 32140 8420
rect 32180 8380 35020 8420
rect 35060 8380 35069 8420
rect 35203 8380 35212 8420
rect 35252 8380 37820 8420
rect 38092 8380 39628 8420
rect 39668 8380 39677 8420
rect 39724 8380 42412 8420
rect 42452 8380 42461 8420
rect 44611 8380 44620 8420
rect 44660 8380 55460 8420
rect 57763 8380 57772 8420
rect 57812 8380 60556 8420
rect 60596 8380 60605 8420
rect 61219 8380 61228 8420
rect 61268 8380 73100 8420
rect 73411 8380 73420 8420
rect 73460 8380 76876 8420
rect 76916 8380 79796 8420
rect 80995 8380 81004 8420
rect 81044 8380 83404 8420
rect 83444 8380 83453 8420
rect 83779 8380 83788 8420
rect 83828 8380 90124 8420
rect 90164 8380 90173 8420
rect 28960 8336 29000 8380
rect 35203 8379 35261 8380
rect 37027 8336 37085 8337
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 9475 8296 9484 8336
rect 9524 8296 10156 8336
rect 10196 8296 10924 8336
rect 10964 8296 17836 8336
rect 17876 8296 17885 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 25315 8296 25324 8336
rect 25364 8296 28588 8336
rect 28628 8296 28637 8336
rect 28960 8296 32908 8336
rect 32948 8296 32957 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 34435 8296 34444 8336
rect 34484 8296 37036 8336
rect 37076 8296 37085 8336
rect 37027 8295 37085 8296
rect 38092 8252 38132 8380
rect 55075 8336 55133 8337
rect 38659 8296 38668 8336
rect 38708 8296 44660 8336
rect 49039 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49425 8336
rect 54595 8296 54604 8336
rect 54644 8296 55084 8336
rect 55124 8296 55133 8336
rect 55420 8336 55460 8380
rect 70627 8336 70685 8337
rect 79756 8336 79796 8380
rect 83779 8379 83837 8380
rect 55420 8296 62092 8336
rect 62132 8296 62141 8336
rect 64159 8296 64168 8336
rect 64208 8296 64250 8336
rect 64290 8296 64332 8336
rect 64372 8296 64414 8336
rect 64454 8296 64496 8336
rect 64536 8296 64545 8336
rect 70627 8296 70636 8336
rect 70676 8296 73324 8336
rect 73364 8296 73373 8336
rect 74371 8296 74380 8336
rect 74420 8296 78988 8336
rect 79028 8296 79037 8336
rect 79279 8296 79288 8336
rect 79328 8296 79370 8336
rect 79410 8296 79452 8336
rect 79492 8296 79534 8336
rect 79574 8296 79616 8336
rect 79656 8296 79665 8336
rect 79756 8296 81140 8336
rect 81571 8296 81580 8336
rect 81620 8296 85900 8336
rect 85940 8296 85949 8336
rect 87811 8296 87820 8336
rect 87860 8296 88204 8336
rect 88244 8296 89452 8336
rect 89492 8296 89501 8336
rect 94399 8296 94408 8336
rect 94448 8296 94490 8336
rect 94530 8296 94572 8336
rect 94612 8296 94654 8336
rect 94694 8296 94736 8336
rect 94776 8296 94785 8336
rect 44620 8252 44660 8296
rect 55075 8295 55133 8296
rect 70627 8295 70685 8296
rect 81100 8252 81140 8296
rect 83683 8252 83741 8253
rect 8419 8212 8428 8252
rect 8468 8212 9140 8252
rect 12931 8212 12940 8252
rect 12980 8212 25132 8252
rect 25172 8212 28012 8252
rect 28052 8212 28684 8252
rect 28724 8212 28733 8252
rect 30787 8212 30796 8252
rect 30836 8212 34828 8252
rect 34868 8212 34877 8252
rect 35011 8212 35020 8252
rect 35060 8212 35444 8252
rect 36739 8212 36748 8252
rect 36788 8212 38132 8252
rect 38179 8212 38188 8252
rect 38228 8212 44140 8252
rect 44180 8212 44189 8252
rect 44611 8212 44620 8252
rect 44660 8212 44669 8252
rect 49507 8212 49516 8252
rect 49556 8212 50764 8252
rect 50804 8212 51148 8252
rect 51188 8212 51340 8252
rect 51380 8212 51389 8252
rect 52675 8212 52684 8252
rect 52724 8212 59828 8252
rect 63619 8212 63628 8252
rect 63668 8212 71116 8252
rect 71156 8212 74956 8252
rect 74996 8212 78124 8252
rect 78164 8212 81004 8252
rect 81044 8212 81053 8252
rect 81100 8212 83692 8252
rect 83732 8212 83741 8252
rect 1987 8128 1996 8168
rect 2036 8128 8812 8168
rect 8852 8128 8861 8168
rect 9100 8084 9140 8212
rect 19180 8168 19220 8212
rect 35404 8168 35444 8212
rect 57955 8168 58013 8169
rect 59788 8168 59828 8212
rect 83683 8211 83741 8212
rect 83788 8212 89932 8252
rect 89972 8212 89981 8252
rect 83788 8168 83828 8212
rect 88675 8168 88733 8169
rect 89251 8168 89309 8169
rect 9283 8128 9292 8168
rect 9332 8128 10060 8168
rect 10100 8128 11980 8168
rect 12020 8128 12748 8168
rect 12788 8128 13132 8168
rect 13172 8128 13516 8168
rect 13556 8128 14188 8168
rect 14228 8128 14237 8168
rect 14284 8128 18796 8168
rect 18836 8128 18845 8168
rect 19171 8128 19180 8168
rect 19220 8128 19229 8168
rect 24547 8128 24556 8168
rect 24596 8128 28204 8168
rect 28244 8128 28253 8168
rect 32899 8128 32908 8168
rect 32948 8128 34636 8168
rect 34676 8128 35308 8168
rect 35348 8128 35357 8168
rect 35404 8128 38420 8168
rect 39043 8128 39052 8168
rect 39092 8128 47500 8168
rect 47540 8128 47549 8168
rect 48259 8128 48268 8168
rect 48308 8128 49420 8168
rect 49460 8128 49469 8168
rect 49804 8128 57772 8168
rect 57812 8128 57821 8168
rect 57955 8128 57964 8168
rect 58004 8128 58732 8168
rect 58772 8128 58781 8168
rect 59788 8128 66412 8168
rect 66452 8128 66461 8168
rect 72067 8128 72076 8168
rect 72116 8128 72556 8168
rect 72596 8128 72605 8168
rect 75043 8128 75052 8168
rect 75092 8128 75244 8168
rect 75284 8128 75916 8168
rect 75956 8128 75965 8168
rect 76867 8128 76876 8168
rect 76916 8128 80908 8168
rect 80948 8128 80957 8168
rect 81763 8128 81772 8168
rect 81812 8128 83596 8168
rect 83636 8128 83645 8168
rect 83779 8128 83788 8168
rect 83828 8128 83837 8168
rect 87523 8128 87532 8168
rect 87572 8128 88204 8168
rect 88244 8128 88253 8168
rect 88590 8128 88684 8168
rect 88724 8128 88733 8168
rect 89166 8128 89260 8168
rect 89300 8128 89309 8168
rect 14284 8084 14324 8128
rect 31939 8084 31997 8085
rect 9100 8044 12460 8084
rect 12500 8044 12509 8084
rect 13315 8044 13324 8084
rect 13364 8044 14324 8084
rect 17827 8044 17836 8084
rect 17876 8044 25900 8084
rect 25940 8044 28972 8084
rect 29012 8044 29021 8084
rect 31267 8044 31276 8084
rect 31316 8044 31948 8084
rect 31988 8044 31997 8084
rect 33763 8044 33772 8084
rect 33812 8044 37708 8084
rect 37748 8044 38284 8084
rect 38324 8044 38333 8084
rect 31939 8043 31997 8044
rect 32419 8000 32477 8001
rect 37219 8000 37277 8001
rect 9859 7960 9868 8000
rect 9908 7960 10252 8000
rect 10292 7960 10636 8000
rect 10676 7960 10685 8000
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 15052 7960 19564 8000
rect 19604 7960 19613 8000
rect 20035 7960 20044 8000
rect 20084 7960 25132 8000
rect 25172 7960 28876 8000
rect 28916 7960 32140 8000
rect 32180 7960 32189 8000
rect 32334 7960 32428 8000
rect 32468 7960 32477 8000
rect 34915 7960 34924 8000
rect 34964 7960 37228 8000
rect 37268 7960 37277 8000
rect 38380 8000 38420 8128
rect 49804 8084 49844 8128
rect 57955 8127 58013 8128
rect 88675 8127 88733 8128
rect 89251 8127 89309 8128
rect 56803 8084 56861 8085
rect 59971 8084 60029 8085
rect 74851 8084 74909 8085
rect 81667 8084 81725 8085
rect 39715 8044 39724 8084
rect 39764 8044 49844 8084
rect 56611 8044 56620 8084
rect 56660 8044 56812 8084
rect 56852 8044 58444 8084
rect 58484 8044 59212 8084
rect 59252 8044 59261 8084
rect 59491 8044 59500 8084
rect 59540 8044 59980 8084
rect 60020 8044 60029 8084
rect 64675 8044 64684 8084
rect 64724 8044 70732 8084
rect 70772 8044 74380 8084
rect 74420 8044 74429 8084
rect 74851 8044 74860 8084
rect 74900 8044 78988 8084
rect 79028 8044 81676 8084
rect 81716 8044 81725 8084
rect 82147 8044 82156 8084
rect 82196 8044 82828 8084
rect 82868 8044 82877 8084
rect 83011 8044 83020 8084
rect 83060 8044 83252 8084
rect 85219 8044 85228 8084
rect 85268 8044 93964 8084
rect 94004 8044 94013 8084
rect 56803 8043 56861 8044
rect 59971 8043 60029 8044
rect 74851 8043 74909 8044
rect 81667 8043 81725 8044
rect 45283 8000 45341 8001
rect 45571 8000 45629 8001
rect 83212 8000 83252 8044
rect 38380 7960 40396 8000
rect 40436 7960 40445 8000
rect 45283 7960 45292 8000
rect 45332 7960 45388 8000
rect 45428 7960 45437 8000
rect 45486 7960 45580 8000
rect 45620 7960 45629 8000
rect 47299 7960 47308 8000
rect 47348 7960 51340 8000
rect 51380 7960 54412 8000
rect 54452 7960 54461 8000
rect 54691 7960 54700 8000
rect 54740 7960 58348 8000
rect 58388 7960 58397 8000
rect 62083 7960 62092 8000
rect 62132 7960 64280 8000
rect 67843 7960 67852 8000
rect 67892 7960 70348 8000
rect 70388 7960 73100 8000
rect 73987 7960 73996 8000
rect 74036 7960 77548 8000
rect 77588 7960 82060 8000
rect 82100 7960 83116 8000
rect 83156 7960 83165 8000
rect 83212 7960 83788 8000
rect 83828 7960 83837 8000
rect 84835 7960 84844 8000
rect 84884 7960 94252 8000
rect 94292 7960 94301 8000
rect 12076 7916 12116 7960
rect 8899 7876 8908 7916
rect 8948 7876 9292 7916
rect 9332 7876 9341 7916
rect 9667 7876 9676 7916
rect 9716 7876 11020 7916
rect 11060 7876 11069 7916
rect 12076 7876 12364 7916
rect 12404 7876 12940 7916
rect 12980 7876 12989 7916
rect 9676 7832 9716 7876
rect 9091 7792 9100 7832
rect 9140 7792 9716 7832
rect 11320 7792 11692 7832
rect 11732 7792 11741 7832
rect 12067 7792 12076 7832
rect 12116 7792 14284 7832
rect 14324 7792 14333 7832
rect 11320 7748 11360 7792
rect 15052 7748 15092 7960
rect 32419 7959 32477 7960
rect 37219 7959 37277 7960
rect 45283 7959 45341 7960
rect 45571 7959 45629 7960
rect 32995 7916 33053 7917
rect 33187 7916 33245 7917
rect 36163 7916 36221 7917
rect 42115 7916 42173 7917
rect 44035 7916 44093 7917
rect 46915 7916 46973 7917
rect 62659 7916 62717 7917
rect 18019 7876 18028 7916
rect 18068 7876 18220 7916
rect 18260 7876 18604 7916
rect 18644 7876 18988 7916
rect 19028 7876 19372 7916
rect 19412 7876 20428 7916
rect 20468 7876 20477 7916
rect 22627 7876 22636 7916
rect 22676 7876 23308 7916
rect 23348 7876 23596 7916
rect 23636 7876 23645 7916
rect 24067 7876 24076 7916
rect 24116 7876 24556 7916
rect 24596 7876 24605 7916
rect 24739 7876 24748 7916
rect 24788 7876 24940 7916
rect 24980 7876 25516 7916
rect 25556 7876 25708 7916
rect 25748 7876 25757 7916
rect 27619 7876 27628 7916
rect 27668 7876 28012 7916
rect 28052 7876 28396 7916
rect 28436 7876 28780 7916
rect 28820 7876 28829 7916
rect 28963 7876 28972 7916
rect 29012 7876 30796 7916
rect 30836 7876 30845 7916
rect 30979 7876 30988 7916
rect 31028 7876 31180 7916
rect 31220 7876 31564 7916
rect 31604 7876 31948 7916
rect 31988 7876 32372 7916
rect 32803 7876 32812 7916
rect 32852 7876 33004 7916
rect 33044 7876 33053 7916
rect 33102 7876 33196 7916
rect 33236 7876 33245 7916
rect 33571 7876 33580 7916
rect 33620 7876 33629 7916
rect 34435 7876 34444 7916
rect 34484 7876 34828 7916
rect 34868 7876 34877 7916
rect 36078 7876 36172 7916
rect 36212 7876 36221 7916
rect 36739 7876 36748 7916
rect 36788 7876 37420 7916
rect 37460 7876 37469 7916
rect 37780 7876 41164 7916
rect 41204 7876 41213 7916
rect 42030 7876 42124 7916
rect 42164 7876 42173 7916
rect 43363 7876 43372 7916
rect 43412 7876 44044 7916
rect 44084 7876 44093 7916
rect 44995 7876 45004 7916
rect 45044 7876 45868 7916
rect 45908 7876 46156 7916
rect 46196 7876 46205 7916
rect 46531 7876 46540 7916
rect 46580 7876 46589 7916
rect 46830 7876 46924 7916
rect 46964 7876 46973 7916
rect 49603 7876 49612 7916
rect 49652 7876 50092 7916
rect 50132 7876 50141 7916
rect 54787 7876 54796 7916
rect 54836 7876 55372 7916
rect 55412 7876 55421 7916
rect 56131 7876 56140 7916
rect 56180 7876 57868 7916
rect 57908 7876 58252 7916
rect 58292 7876 58828 7916
rect 58868 7876 58877 7916
rect 62574 7876 62668 7916
rect 62708 7876 62717 7916
rect 64240 7916 64280 7960
rect 66787 7916 66845 7917
rect 67651 7916 67709 7917
rect 72067 7916 72125 7917
rect 64240 7876 65260 7916
rect 65300 7876 65309 7916
rect 66787 7876 66796 7916
rect 66836 7876 67180 7916
rect 67220 7876 67229 7916
rect 67566 7876 67660 7916
rect 67700 7876 67709 7916
rect 68899 7876 68908 7916
rect 68948 7876 69772 7916
rect 69812 7876 69821 7916
rect 69955 7876 69964 7916
rect 70004 7876 70156 7916
rect 70196 7876 70540 7916
rect 70580 7876 70924 7916
rect 70964 7876 71692 7916
rect 71732 7876 71741 7916
rect 72067 7876 72076 7916
rect 72116 7876 72748 7916
rect 72788 7876 72797 7916
rect 17443 7832 17501 7833
rect 19948 7832 19988 7876
rect 24643 7832 24701 7833
rect 30883 7832 30941 7833
rect 31267 7832 31325 7833
rect 31843 7832 31901 7833
rect 32035 7832 32093 7833
rect 32332 7832 32372 7876
rect 32995 7875 33053 7876
rect 33187 7875 33245 7876
rect 33580 7832 33620 7876
rect 36163 7875 36221 7876
rect 37780 7832 37820 7876
rect 42115 7875 42173 7876
rect 44035 7875 44093 7876
rect 45091 7832 45149 7833
rect 46540 7832 46580 7876
rect 46915 7875 46973 7876
rect 62659 7875 62717 7876
rect 66787 7875 66845 7876
rect 67651 7875 67709 7876
rect 72067 7875 72125 7876
rect 73060 7832 73100 7960
rect 83212 7916 83252 7960
rect 85603 7916 85661 7917
rect 74179 7876 74188 7916
rect 74228 7876 74572 7916
rect 74612 7876 74621 7916
rect 77731 7876 77740 7916
rect 77780 7876 78412 7916
rect 78452 7876 78796 7916
rect 78836 7876 78845 7916
rect 80707 7876 80716 7916
rect 80756 7876 81099 7916
rect 81139 7876 81484 7916
rect 81524 7876 81868 7916
rect 81908 7876 81917 7916
rect 82435 7876 82444 7916
rect 82484 7876 82828 7916
rect 82868 7876 82877 7916
rect 82924 7876 83212 7916
rect 83252 7876 83261 7916
rect 83395 7876 83404 7916
rect 83444 7876 83980 7916
rect 84020 7876 84029 7916
rect 84163 7876 84172 7916
rect 84212 7876 84556 7916
rect 84596 7876 84940 7916
rect 84980 7876 84989 7916
rect 85603 7876 85612 7916
rect 85652 7876 88396 7916
rect 88436 7876 88588 7916
rect 88628 7876 88637 7916
rect 82924 7832 82964 7876
rect 84172 7832 84212 7876
rect 85603 7875 85661 7876
rect 17443 7792 17452 7832
rect 17492 7792 17932 7832
rect 17972 7792 17981 7832
rect 18787 7792 18796 7832
rect 18836 7792 19276 7832
rect 19316 7792 19325 7832
rect 19939 7792 19948 7832
rect 19988 7792 19997 7832
rect 20611 7792 20620 7832
rect 20660 7792 20812 7832
rect 20852 7792 23020 7832
rect 23060 7792 23069 7832
rect 23203 7792 23212 7832
rect 23252 7792 24652 7832
rect 24692 7792 24701 7832
rect 25027 7792 25036 7832
rect 25076 7792 26476 7832
rect 26516 7792 26525 7832
rect 30798 7792 30892 7832
rect 30932 7792 30941 7832
rect 31182 7792 31276 7832
rect 31316 7792 31325 7832
rect 31651 7792 31660 7832
rect 31700 7792 31852 7832
rect 31892 7792 31901 7832
rect 31950 7792 32044 7832
rect 32084 7792 32093 7832
rect 32323 7792 32332 7832
rect 32372 7792 32716 7832
rect 32756 7792 33100 7832
rect 33140 7792 33620 7832
rect 33859 7792 33868 7832
rect 33908 7792 34772 7832
rect 35011 7792 35020 7832
rect 35060 7792 37820 7832
rect 44227 7792 44236 7832
rect 44276 7792 45100 7832
rect 45140 7792 46580 7832
rect 48739 7792 48748 7832
rect 48788 7792 49996 7832
rect 50036 7792 50045 7832
rect 65827 7792 65836 7832
rect 65876 7792 70252 7832
rect 70292 7792 70301 7832
rect 73060 7792 75916 7832
rect 75956 7792 75965 7832
rect 76291 7792 76300 7832
rect 76340 7792 78028 7832
rect 78068 7792 78077 7832
rect 80803 7792 80812 7832
rect 80852 7792 81388 7832
rect 81428 7792 81437 7832
rect 82627 7792 82636 7832
rect 82676 7792 82964 7832
rect 83011 7792 83020 7832
rect 83060 7792 84212 7832
rect 84451 7792 84460 7832
rect 84500 7792 87628 7832
rect 87668 7792 87677 7832
rect 88291 7792 88300 7832
rect 88340 7792 96652 7832
rect 96692 7792 96701 7832
rect 17443 7791 17501 7792
rect 24643 7791 24701 7792
rect 30883 7791 30941 7792
rect 31267 7791 31325 7792
rect 31843 7791 31901 7792
rect 32035 7791 32093 7792
rect 34732 7748 34772 7792
rect 45091 7791 45149 7792
rect 54883 7748 54941 7749
rect 59683 7748 59741 7749
rect 75916 7748 75956 7792
rect 88867 7748 88925 7749
rect 2371 7708 2380 7748
rect 2420 7708 7564 7748
rect 7604 7708 7613 7748
rect 8035 7708 8044 7748
rect 8084 7708 11360 7748
rect 11587 7708 11596 7748
rect 11636 7708 12172 7748
rect 12212 7708 15092 7748
rect 18883 7708 18892 7748
rect 18932 7708 25228 7748
rect 25268 7708 27820 7748
rect 27860 7708 27869 7748
rect 28579 7708 28588 7748
rect 28628 7708 31372 7748
rect 31412 7708 34636 7748
rect 34676 7708 34685 7748
rect 34732 7708 39724 7748
rect 39764 7708 39773 7748
rect 41347 7708 41356 7748
rect 41396 7708 45580 7748
rect 45620 7708 45629 7748
rect 45859 7708 45868 7748
rect 45908 7708 46540 7748
rect 46580 7708 47212 7748
rect 47252 7708 47261 7748
rect 49123 7708 49132 7748
rect 49172 7708 49516 7748
rect 49556 7708 49565 7748
rect 54798 7708 54892 7748
rect 54932 7708 54941 7748
rect 56899 7708 56908 7748
rect 56948 7708 58828 7748
rect 58868 7708 58877 7748
rect 59683 7708 59692 7748
rect 59732 7708 59884 7748
rect 59924 7708 59933 7748
rect 67363 7708 67372 7748
rect 67412 7708 70732 7748
rect 70772 7708 73996 7748
rect 74036 7708 74045 7748
rect 75916 7708 77932 7748
rect 77972 7708 81292 7748
rect 81332 7708 84748 7748
rect 84788 7708 84797 7748
rect 84931 7708 84940 7748
rect 84980 7708 85324 7748
rect 85364 7708 86860 7748
rect 86900 7708 86909 7748
rect 87811 7708 87820 7748
rect 87860 7708 88876 7748
rect 88916 7708 89452 7748
rect 89492 7708 89501 7748
rect 95779 7708 95788 7748
rect 95828 7708 98188 7748
rect 98228 7708 98237 7748
rect 22819 7664 22877 7665
rect 10339 7624 10348 7664
rect 10388 7624 13324 7664
rect 13364 7624 13373 7664
rect 13699 7624 13708 7664
rect 13748 7624 19756 7664
rect 19796 7624 19805 7664
rect 22531 7624 22540 7664
rect 22580 7624 22828 7664
rect 22868 7624 22877 7664
rect 27820 7664 27860 7708
rect 54883 7707 54941 7708
rect 59683 7707 59741 7708
rect 36835 7664 36893 7665
rect 44323 7664 44381 7665
rect 75811 7664 75869 7665
rect 78403 7664 78461 7665
rect 83779 7664 83837 7665
rect 83980 7664 84020 7708
rect 88867 7707 88925 7708
rect 27820 7624 33292 7664
rect 33332 7624 35020 7664
rect 35060 7624 35069 7664
rect 36750 7624 36844 7664
rect 36884 7624 36893 7664
rect 42019 7624 42028 7664
rect 42068 7624 44332 7664
rect 44372 7624 44381 7664
rect 55363 7624 55372 7664
rect 55412 7624 56812 7664
rect 56852 7624 57676 7664
rect 57716 7624 58348 7664
rect 58388 7624 59500 7664
rect 59540 7624 59549 7664
rect 66211 7624 66220 7664
rect 66260 7624 73420 7664
rect 73460 7624 73469 7664
rect 74668 7624 75244 7664
rect 75284 7624 75293 7664
rect 75726 7624 75820 7664
rect 75860 7624 75869 7664
rect 76771 7624 76780 7664
rect 76820 7624 77452 7664
rect 77492 7624 77501 7664
rect 78307 7624 78316 7664
rect 78356 7624 78412 7664
rect 78452 7624 78461 7664
rect 83299 7624 83308 7664
rect 83348 7624 83788 7664
rect 83828 7624 83837 7664
rect 83971 7624 83980 7664
rect 84020 7624 84029 7664
rect 84163 7624 84172 7664
rect 84212 7624 88972 7664
rect 89012 7624 89021 7664
rect 89155 7624 89164 7664
rect 89204 7624 97036 7664
rect 97076 7624 97085 7664
rect 22819 7623 22877 7624
rect 36835 7623 36893 7624
rect 44323 7623 44381 7624
rect 19363 7580 19421 7581
rect 74668 7580 74708 7624
rect 75811 7623 75869 7624
rect 78403 7623 78461 7624
rect 83779 7623 83837 7624
rect 74851 7580 74909 7581
rect 77059 7580 77117 7581
rect 82915 7580 82973 7581
rect 88387 7580 88445 7581
rect 88579 7580 88637 7581
rect 89347 7580 89405 7581
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 10435 7540 10444 7580
rect 10484 7540 10636 7580
rect 10676 7540 11360 7580
rect 11320 7496 11360 7540
rect 11404 7540 18892 7580
rect 18932 7540 18941 7580
rect 19363 7540 19372 7580
rect 19412 7540 19852 7580
rect 19892 7540 19901 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 24259 7540 24268 7580
rect 24308 7540 25708 7580
rect 25748 7540 25757 7580
rect 28195 7540 28204 7580
rect 28244 7540 32812 7580
rect 32852 7540 33676 7580
rect 33716 7540 33725 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 36739 7540 36748 7580
rect 36788 7540 37420 7580
rect 37460 7540 37612 7580
rect 37652 7540 37661 7580
rect 44611 7540 44620 7580
rect 44660 7540 45292 7580
rect 45332 7540 45341 7580
rect 45763 7540 45772 7580
rect 45812 7540 46444 7580
rect 46484 7540 47116 7580
rect 47156 7540 47165 7580
rect 49219 7540 49228 7580
rect 49268 7540 49900 7580
rect 49940 7540 49949 7580
rect 50279 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50665 7580
rect 52867 7540 52876 7580
rect 52916 7540 56524 7580
rect 56564 7540 56573 7580
rect 57763 7540 57772 7580
rect 57812 7540 60500 7580
rect 60643 7540 60652 7580
rect 60692 7540 62380 7580
rect 62420 7540 62429 7580
rect 65399 7540 65408 7580
rect 65448 7540 65490 7580
rect 65530 7540 65572 7580
rect 65612 7540 65654 7580
rect 65694 7540 65736 7580
rect 65776 7540 65785 7580
rect 69763 7540 69772 7580
rect 69812 7540 74708 7580
rect 74766 7540 74860 7580
rect 74900 7540 74909 7580
rect 75043 7540 75052 7580
rect 75092 7540 75436 7580
rect 75476 7540 75485 7580
rect 76974 7540 77068 7580
rect 77108 7540 77117 7580
rect 80519 7540 80528 7580
rect 80568 7540 80610 7580
rect 80650 7540 80692 7580
rect 80732 7540 80774 7580
rect 80814 7540 80856 7580
rect 80896 7540 80905 7580
rect 82830 7540 82924 7580
rect 82964 7540 82973 7580
rect 83779 7540 83788 7580
rect 83828 7540 84020 7580
rect 84067 7540 84076 7580
rect 84116 7540 88396 7580
rect 88436 7540 88445 7580
rect 88494 7540 88588 7580
rect 88628 7540 88637 7580
rect 89262 7540 89356 7580
rect 89396 7540 89405 7580
rect 95639 7540 95648 7580
rect 95688 7540 95730 7580
rect 95770 7540 95812 7580
rect 95852 7540 95894 7580
rect 95934 7540 95976 7580
rect 96016 7540 96025 7580
rect 11404 7496 11444 7540
rect 19363 7539 19421 7540
rect 30115 7496 30173 7497
rect 33763 7496 33821 7497
rect 37891 7496 37949 7497
rect 11320 7456 11444 7496
rect 11683 7456 11692 7496
rect 11732 7456 11884 7496
rect 11924 7456 11933 7496
rect 12547 7456 12556 7496
rect 12596 7456 12748 7496
rect 12788 7456 12797 7496
rect 13516 7456 18412 7496
rect 18452 7456 18461 7496
rect 19267 7456 19276 7496
rect 19316 7456 24172 7496
rect 24212 7456 24221 7496
rect 30019 7456 30028 7496
rect 30068 7456 30124 7496
rect 30164 7456 30173 7496
rect 30979 7456 30988 7496
rect 31028 7456 33772 7496
rect 33812 7456 37228 7496
rect 37268 7456 37277 7496
rect 37507 7456 37516 7496
rect 37556 7456 37900 7496
rect 37940 7456 37949 7496
rect 39235 7456 39244 7496
rect 39284 7456 50764 7496
rect 50804 7456 50813 7496
rect 50947 7456 50956 7496
rect 50996 7456 54356 7496
rect 55843 7456 55852 7496
rect 55892 7456 59828 7496
rect 13516 7412 13556 7456
rect 30115 7455 30173 7456
rect 33763 7455 33821 7456
rect 37891 7455 37949 7456
rect 19267 7412 19325 7413
rect 54316 7412 54356 7456
rect 10051 7372 10060 7412
rect 10100 7372 13556 7412
rect 13603 7372 13612 7412
rect 13652 7372 14188 7412
rect 14228 7372 14237 7412
rect 18691 7372 18700 7412
rect 18740 7372 19276 7412
rect 19316 7372 19325 7412
rect 22627 7372 22636 7412
rect 22676 7372 22828 7412
rect 22868 7372 23020 7412
rect 23060 7372 23069 7412
rect 24451 7372 24460 7412
rect 24500 7372 29548 7412
rect 29588 7372 29597 7412
rect 33283 7372 33292 7412
rect 33332 7372 33868 7412
rect 33908 7372 33917 7412
rect 34627 7372 34636 7412
rect 34676 7372 42988 7412
rect 43028 7372 43037 7412
rect 45955 7372 45964 7412
rect 46004 7372 46636 7412
rect 46676 7372 46685 7412
rect 50563 7372 50572 7412
rect 50612 7372 51244 7412
rect 51284 7372 51532 7412
rect 51572 7372 51581 7412
rect 51907 7372 51916 7412
rect 51956 7372 52204 7412
rect 52244 7372 52253 7412
rect 54307 7372 54316 7412
rect 54356 7372 55756 7412
rect 55796 7372 56140 7412
rect 56180 7372 56189 7412
rect 59395 7372 59404 7412
rect 59444 7372 59692 7412
rect 59732 7372 59741 7412
rect 10060 7328 10100 7372
rect 19267 7371 19325 7372
rect 34435 7328 34493 7329
rect 56227 7328 56285 7329
rect 59683 7328 59741 7329
rect 9676 7288 10100 7328
rect 10147 7288 10156 7328
rect 10196 7288 10348 7328
rect 10388 7288 10397 7328
rect 10819 7288 10828 7328
rect 10868 7288 10908 7328
rect 11875 7288 11884 7328
rect 11924 7288 13708 7328
rect 13748 7288 13757 7328
rect 23116 7288 23596 7328
rect 23636 7288 24748 7328
rect 24788 7288 24797 7328
rect 34435 7288 34444 7328
rect 34484 7288 37708 7328
rect 37748 7288 37757 7328
rect 39523 7288 39532 7328
rect 39572 7288 55460 7328
rect 56142 7288 56236 7328
rect 56276 7288 56285 7328
rect 9676 7244 9716 7288
rect 10828 7244 10868 7288
rect 22915 7244 22973 7245
rect 23116 7244 23156 7288
rect 34435 7287 34493 7288
rect 25699 7244 25757 7245
rect 30019 7244 30077 7245
rect 33763 7244 33821 7245
rect 40099 7244 40157 7245
rect 55420 7244 55460 7288
rect 56227 7287 56285 7288
rect 57868 7288 59692 7328
rect 59732 7288 59741 7328
rect 57868 7244 57908 7288
rect 59683 7287 59741 7288
rect 59788 7328 59828 7456
rect 59875 7412 59933 7413
rect 59875 7372 59884 7412
rect 59924 7372 60364 7412
rect 60404 7372 60413 7412
rect 59875 7371 59933 7372
rect 60259 7328 60317 7329
rect 59788 7288 60268 7328
rect 60308 7288 60409 7328
rect 59788 7244 59828 7288
rect 60259 7287 60317 7288
rect 60369 7244 60409 7288
rect 60460 7244 60500 7540
rect 74851 7539 74909 7540
rect 77059 7539 77117 7540
rect 82915 7539 82973 7540
rect 64003 7496 64061 7497
rect 83980 7496 84020 7540
rect 88387 7539 88445 7540
rect 88579 7539 88637 7540
rect 89347 7539 89405 7540
rect 88195 7496 88253 7497
rect 88675 7496 88733 7497
rect 60739 7456 60748 7496
rect 60788 7456 64012 7496
rect 64052 7456 64061 7496
rect 72835 7456 72844 7496
rect 72884 7456 74764 7496
rect 74804 7456 74813 7496
rect 80419 7456 80428 7496
rect 80468 7456 83884 7496
rect 83924 7456 83933 7496
rect 83980 7456 84172 7496
rect 84212 7456 84221 7496
rect 88195 7456 88204 7496
rect 88244 7456 88338 7496
rect 88675 7456 88684 7496
rect 88724 7456 88780 7496
rect 88820 7456 88829 7496
rect 64003 7455 64061 7456
rect 88195 7455 88253 7456
rect 88675 7455 88733 7456
rect 74947 7412 75005 7413
rect 78883 7412 78941 7413
rect 60547 7372 60556 7412
rect 60596 7372 61708 7412
rect 61748 7372 71500 7412
rect 71540 7372 71549 7412
rect 71875 7372 71884 7412
rect 71924 7372 74476 7412
rect 74516 7372 74525 7412
rect 74862 7372 74956 7412
rect 74996 7372 75005 7412
rect 78798 7372 78892 7412
rect 78932 7372 78941 7412
rect 79171 7372 79180 7412
rect 79220 7372 85516 7412
rect 85556 7372 85565 7412
rect 85699 7372 85708 7412
rect 85748 7372 91948 7412
rect 91988 7372 91997 7412
rect 74947 7371 75005 7372
rect 78883 7371 78941 7372
rect 71011 7328 71069 7329
rect 88195 7328 88253 7329
rect 64003 7288 64012 7328
rect 64052 7288 71020 7328
rect 71060 7288 71069 7328
rect 77731 7288 77740 7328
rect 77780 7288 78508 7328
rect 78548 7288 78557 7328
rect 78691 7288 78700 7328
rect 78740 7288 80812 7328
rect 80852 7288 87572 7328
rect 87715 7288 87724 7328
rect 87764 7288 88204 7328
rect 88244 7288 88253 7328
rect 71011 7287 71069 7288
rect 63043 7244 63101 7245
rect 64483 7244 64541 7245
rect 66787 7244 66845 7245
rect 81859 7244 81917 7245
rect 83683 7244 83741 7245
rect 87532 7244 87572 7288
rect 88195 7287 88253 7288
rect 9667 7204 9676 7244
rect 9716 7204 9725 7244
rect 9859 7204 9868 7244
rect 9908 7204 10540 7244
rect 10580 7204 11212 7244
rect 11252 7204 11261 7244
rect 13603 7204 13612 7244
rect 13652 7204 17164 7244
rect 17204 7204 22732 7244
rect 22772 7204 22781 7244
rect 22915 7204 22924 7244
rect 22964 7204 23058 7244
rect 23107 7204 23116 7244
rect 23156 7204 23165 7244
rect 24067 7204 24076 7244
rect 24116 7204 24364 7244
rect 24404 7204 24413 7244
rect 25123 7204 25132 7244
rect 25172 7204 25708 7244
rect 25748 7204 25757 7244
rect 26947 7204 26956 7244
rect 26996 7204 27005 7244
rect 29934 7204 30028 7244
rect 30068 7204 30077 7244
rect 31939 7204 31948 7244
rect 31988 7204 32140 7244
rect 32180 7204 32189 7244
rect 32323 7204 32332 7244
rect 32372 7204 32381 7244
rect 33763 7204 33772 7244
rect 33812 7204 33868 7244
rect 33908 7204 33917 7244
rect 34051 7204 34060 7244
rect 34100 7204 34348 7244
rect 34388 7204 34397 7244
rect 34627 7204 34636 7244
rect 34676 7204 37324 7244
rect 37364 7204 37373 7244
rect 37507 7204 37516 7244
rect 37556 7204 37900 7244
rect 37940 7204 38284 7244
rect 38324 7204 38333 7244
rect 40014 7204 40108 7244
rect 40148 7204 40157 7244
rect 43459 7204 43468 7244
rect 43508 7204 43948 7244
rect 43988 7204 43997 7244
rect 44419 7204 44428 7244
rect 44468 7204 44908 7244
rect 44948 7204 45196 7244
rect 45236 7204 45245 7244
rect 48163 7204 48172 7244
rect 48212 7204 48364 7244
rect 48404 7204 49324 7244
rect 49364 7204 49373 7244
rect 50755 7204 50764 7244
rect 50804 7204 51244 7244
rect 51284 7204 51436 7244
rect 51476 7204 51628 7244
rect 51668 7204 51677 7244
rect 51907 7204 51916 7244
rect 51956 7204 52300 7244
rect 52340 7204 53068 7244
rect 53108 7204 53117 7244
rect 55420 7204 57908 7244
rect 59779 7204 59788 7244
rect 59828 7204 59837 7244
rect 59971 7204 59980 7244
rect 60020 7204 60268 7244
rect 60308 7204 60317 7244
rect 60360 7204 60369 7244
rect 60409 7204 60418 7244
rect 60460 7204 60652 7244
rect 60692 7204 60701 7244
rect 61891 7204 61900 7244
rect 61940 7204 62188 7244
rect 62228 7204 62237 7244
rect 62958 7204 63052 7244
rect 63092 7204 63101 7244
rect 64398 7204 64492 7244
rect 64532 7204 64541 7244
rect 66702 7204 66796 7244
rect 66836 7204 66845 7244
rect 68035 7204 68044 7244
rect 68084 7204 68716 7244
rect 68756 7204 69196 7244
rect 69236 7204 69245 7244
rect 72355 7204 72364 7244
rect 72404 7204 77260 7244
rect 77300 7204 77309 7244
rect 77539 7204 77548 7244
rect 77588 7204 78604 7244
rect 78644 7204 78653 7244
rect 81859 7204 81868 7244
rect 81908 7204 82636 7244
rect 82676 7204 82685 7244
rect 83011 7204 83020 7244
rect 83060 7204 83404 7244
rect 83444 7204 83453 7244
rect 83683 7204 83692 7244
rect 83732 7204 85556 7244
rect 85603 7204 85612 7244
rect 85652 7204 86380 7244
rect 86420 7204 86429 7244
rect 87523 7204 87532 7244
rect 87572 7204 87581 7244
rect 22915 7203 22973 7204
rect 25699 7203 25757 7204
rect 26956 7160 26996 7204
rect 30019 7203 30077 7204
rect 32332 7160 32372 7204
rect 33763 7203 33821 7204
rect 36451 7160 36509 7161
rect 5347 7120 5356 7160
rect 5396 7120 12268 7160
rect 12308 7120 12317 7160
rect 12835 7120 12844 7160
rect 12884 7120 13132 7160
rect 13172 7120 13181 7160
rect 23203 7120 23212 7160
rect 23252 7120 29000 7160
rect 29827 7120 29836 7160
rect 29876 7120 31660 7160
rect 31700 7120 33196 7160
rect 33236 7120 33245 7160
rect 34243 7120 34252 7160
rect 34292 7120 34732 7160
rect 34772 7120 34781 7160
rect 36366 7120 36460 7160
rect 36500 7120 36509 7160
rect 28960 7076 29000 7120
rect 36451 7119 36509 7120
rect 34531 7076 34589 7077
rect 9475 7036 9484 7076
rect 9524 7036 9964 7076
rect 10004 7036 10013 7076
rect 19075 7036 19084 7076
rect 19124 7036 21004 7076
rect 21044 7036 21053 7076
rect 23299 7036 23308 7076
rect 23348 7036 24460 7076
rect 24500 7036 25036 7076
rect 25076 7036 25085 7076
rect 28960 7036 32276 7076
rect 32323 7036 32332 7076
rect 32372 7036 33292 7076
rect 33332 7036 33341 7076
rect 34446 7036 34540 7076
rect 34580 7036 34589 7076
rect 37324 7076 37364 7204
rect 40099 7203 40157 7204
rect 63043 7203 63101 7204
rect 64483 7203 64541 7204
rect 66787 7203 66845 7204
rect 81859 7203 81917 7204
rect 83683 7203 83741 7204
rect 46339 7160 46397 7161
rect 37699 7120 37708 7160
rect 37748 7120 41932 7160
rect 41972 7120 41981 7160
rect 46254 7120 46348 7160
rect 46388 7120 46397 7160
rect 46627 7120 46636 7160
rect 46676 7120 48652 7160
rect 48692 7120 48701 7160
rect 51715 7120 51724 7160
rect 51764 7120 52108 7160
rect 52148 7120 52780 7160
rect 52820 7120 52829 7160
rect 56227 7120 56236 7160
rect 56276 7120 62476 7160
rect 62516 7120 62525 7160
rect 66211 7120 66220 7160
rect 66260 7120 68236 7160
rect 68276 7120 74565 7160
rect 74605 7120 74614 7160
rect 75235 7120 75244 7160
rect 75284 7120 76876 7160
rect 76916 7120 78028 7160
rect 78068 7120 78077 7160
rect 82819 7120 82828 7160
rect 82868 7120 84076 7160
rect 84116 7120 84125 7160
rect 46339 7119 46397 7120
rect 51811 7076 51869 7077
rect 85516 7076 85556 7204
rect 85699 7120 85708 7160
rect 85748 7120 85996 7160
rect 86036 7120 86045 7160
rect 86275 7120 86284 7160
rect 86324 7120 87340 7160
rect 87380 7120 87389 7160
rect 87619 7120 87628 7160
rect 87668 7120 95500 7160
rect 95540 7120 95549 7160
rect 88195 7076 88253 7077
rect 37324 7036 39340 7076
rect 39380 7036 39389 7076
rect 42883 7036 42892 7076
rect 42932 7036 51668 7076
rect 51726 7036 51820 7076
rect 51860 7036 64012 7076
rect 64052 7036 64061 7076
rect 66979 7036 66988 7076
rect 67028 7036 67948 7076
rect 67988 7036 73100 7076
rect 74275 7036 74284 7076
rect 74324 7036 78508 7076
rect 78548 7036 78557 7076
rect 78988 7036 84652 7076
rect 84692 7036 84701 7076
rect 85516 7036 85804 7076
rect 85844 7036 86860 7076
rect 86900 7036 88012 7076
rect 88052 7036 88061 7076
rect 88195 7036 88204 7076
rect 88244 7036 88338 7076
rect 88675 7036 88684 7076
rect 88724 7036 90508 7076
rect 90548 7036 90557 7076
rect 23491 6992 23549 6993
rect 6499 6952 6508 6992
rect 6548 6952 9772 6992
rect 9812 6952 9821 6992
rect 11203 6952 11212 6992
rect 11252 6952 11788 6992
rect 11828 6952 12076 6992
rect 12116 6952 12748 6992
rect 12788 6952 13420 6992
rect 13460 6952 13469 6992
rect 18787 6952 18796 6992
rect 18836 6952 20716 6992
rect 20756 6952 20765 6992
rect 23491 6952 23500 6992
rect 23540 6952 24364 6992
rect 24404 6952 24413 6992
rect 24739 6952 24748 6992
rect 24788 6952 30988 6992
rect 31028 6952 31037 6992
rect 31171 6952 31180 6992
rect 31220 6952 32140 6992
rect 32180 6952 32189 6992
rect 23491 6951 23549 6952
rect 12547 6908 12605 6909
rect 32236 6908 32276 7036
rect 34531 7035 34589 7036
rect 34819 6992 34877 6993
rect 37507 6992 37565 6993
rect 48931 6992 48989 6993
rect 51628 6992 51668 7036
rect 51811 7035 51869 7036
rect 59971 6992 60029 6993
rect 33955 6952 33964 6992
rect 34004 6952 34828 6992
rect 34868 6952 34877 6992
rect 36163 6952 36172 6992
rect 36212 6952 36652 6992
rect 36692 6952 36701 6992
rect 37422 6952 37516 6992
rect 37556 6952 37565 6992
rect 44515 6952 44524 6992
rect 44564 6952 46636 6992
rect 46676 6952 46685 6992
rect 48931 6952 48940 6992
rect 48980 6952 49036 6992
rect 49076 6952 49085 6992
rect 49315 6952 49324 6992
rect 49364 6952 50804 6992
rect 51628 6952 52108 6992
rect 52148 6952 57868 6992
rect 57908 6952 57917 6992
rect 58531 6952 58540 6992
rect 58580 6952 59788 6992
rect 59828 6952 59837 6992
rect 59971 6952 59980 6992
rect 60020 6952 60114 6992
rect 60547 6952 60556 6992
rect 60596 6952 61036 6992
rect 61076 6952 61085 6992
rect 34819 6951 34877 6952
rect 37507 6951 37565 6952
rect 48931 6951 48989 6952
rect 36451 6908 36509 6909
rect 50764 6908 50804 6952
rect 59971 6951 60029 6952
rect 55747 6908 55805 6909
rect 56131 6908 56189 6909
rect 73060 6908 73100 7036
rect 74083 6992 74141 6993
rect 78988 6992 79028 7036
rect 88195 7035 88253 7036
rect 74083 6952 74092 6992
rect 74132 6952 74188 6992
rect 74228 6952 74237 6992
rect 74467 6952 74476 6992
rect 74516 6952 75628 6992
rect 75668 6952 75677 6992
rect 77740 6952 78988 6992
rect 79028 6952 79037 6992
rect 79171 6952 79180 6992
rect 79220 6952 82868 6992
rect 82915 6952 82924 6992
rect 82964 6952 82973 6992
rect 83491 6952 83500 6992
rect 83540 6952 86572 6992
rect 86612 6952 86621 6992
rect 87331 6952 87340 6992
rect 87380 6952 88108 6992
rect 88148 6952 88157 6992
rect 74083 6951 74141 6952
rect 75043 6908 75101 6909
rect 77740 6908 77780 6952
rect 5731 6868 5740 6908
rect 5780 6868 12556 6908
rect 12596 6868 12605 6908
rect 15523 6868 15532 6908
rect 15572 6868 16588 6908
rect 16628 6868 17740 6908
rect 17780 6868 24268 6908
rect 24308 6868 27340 6908
rect 27380 6868 31604 6908
rect 32035 6868 32044 6908
rect 32084 6868 34828 6908
rect 34868 6868 34877 6908
rect 36451 6868 36460 6908
rect 36500 6868 39436 6908
rect 39476 6868 46004 6908
rect 47971 6868 47980 6908
rect 48020 6868 48556 6908
rect 48596 6868 50708 6908
rect 50764 6868 52588 6908
rect 52628 6868 55756 6908
rect 55796 6868 56084 6908
rect 12547 6867 12605 6868
rect 26947 6824 27005 6825
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 24163 6784 24172 6824
rect 24212 6784 26956 6824
rect 26996 6784 27005 6824
rect 27907 6784 27916 6824
rect 27956 6784 28396 6824
rect 28436 6784 28445 6824
rect 28960 6784 29740 6824
rect 29780 6784 29789 6824
rect 26947 6783 27005 6784
rect 16195 6740 16253 6741
rect 23395 6740 23453 6741
rect 24547 6740 24605 6741
rect 28960 6740 29000 6784
rect 31564 6740 31604 6868
rect 34723 6824 34781 6825
rect 31651 6784 31660 6824
rect 31700 6784 32236 6824
rect 32276 6784 32285 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 34435 6784 34444 6824
rect 34484 6784 34732 6824
rect 34772 6784 34781 6824
rect 34828 6824 34868 6868
rect 36451 6867 36509 6868
rect 34828 6784 36844 6824
rect 36884 6784 36893 6824
rect 38659 6784 38668 6824
rect 38708 6784 41740 6824
rect 41780 6784 41789 6824
rect 34723 6783 34781 6784
rect 45964 6740 46004 6868
rect 46723 6784 46732 6824
rect 46772 6784 47212 6824
rect 47252 6784 48460 6824
rect 48500 6784 48748 6824
rect 48788 6784 48797 6824
rect 49039 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49425 6824
rect 50668 6740 50708 6868
rect 55747 6867 55805 6868
rect 55555 6824 55613 6825
rect 56044 6824 56084 6868
rect 56131 6868 56140 6908
rect 56180 6868 57196 6908
rect 57236 6868 57245 6908
rect 57667 6868 57676 6908
rect 57716 6868 64972 6908
rect 65012 6868 65021 6908
rect 67075 6868 67084 6908
rect 67124 6868 72844 6908
rect 72884 6868 72893 6908
rect 73060 6868 74996 6908
rect 56131 6867 56189 6868
rect 74956 6824 74996 6868
rect 75043 6868 75052 6908
rect 75092 6868 75148 6908
rect 75188 6868 77356 6908
rect 77396 6868 77740 6908
rect 77780 6868 77789 6908
rect 78691 6868 78700 6908
rect 78740 6868 82156 6908
rect 82196 6868 82205 6908
rect 75043 6867 75101 6868
rect 82828 6824 82868 6952
rect 82924 6908 82964 6952
rect 82924 6868 89644 6908
rect 89684 6868 89693 6908
rect 51427 6784 51436 6824
rect 51476 6784 55460 6824
rect 55420 6740 55460 6784
rect 55555 6784 55564 6824
rect 55604 6784 55660 6824
rect 55700 6784 55709 6824
rect 56035 6784 56044 6824
rect 56084 6784 56093 6824
rect 56515 6784 56524 6824
rect 56564 6784 59212 6824
rect 59252 6784 59261 6824
rect 64159 6784 64168 6824
rect 64208 6784 64250 6824
rect 64290 6784 64332 6824
rect 64372 6784 64414 6824
rect 64454 6784 64496 6824
rect 64536 6784 64545 6824
rect 65155 6784 65164 6824
rect 65204 6784 68044 6824
rect 68084 6784 74284 6824
rect 74324 6784 74333 6824
rect 74947 6784 74956 6824
rect 74996 6784 79180 6824
rect 79220 6784 79229 6824
rect 79279 6784 79288 6824
rect 79328 6784 79370 6824
rect 79410 6784 79452 6824
rect 79492 6784 79534 6824
rect 79574 6784 79616 6824
rect 79656 6784 79665 6824
rect 82819 6784 82828 6824
rect 82868 6784 82877 6824
rect 83107 6784 83116 6824
rect 83156 6784 83788 6824
rect 83828 6784 83837 6824
rect 94399 6784 94408 6824
rect 94448 6784 94490 6824
rect 94530 6784 94572 6824
rect 94612 6784 94654 6824
rect 94694 6784 94736 6824
rect 94776 6784 94785 6824
rect 55555 6783 55613 6784
rect 10051 6700 10060 6740
rect 10100 6700 15244 6740
rect 15284 6700 15293 6740
rect 16110 6700 16204 6740
rect 16244 6700 16253 6740
rect 19459 6700 19468 6740
rect 19508 6700 21100 6740
rect 21140 6700 21149 6740
rect 23310 6700 23404 6740
rect 23444 6700 23453 6740
rect 24462 6700 24556 6740
rect 24596 6700 24605 6740
rect 25027 6700 25036 6740
rect 25076 6700 29000 6740
rect 31555 6700 31564 6740
rect 31604 6700 33676 6740
rect 33716 6700 38092 6740
rect 38132 6700 38141 6740
rect 45964 6700 49844 6740
rect 50659 6700 50668 6740
rect 50708 6700 53356 6740
rect 53396 6700 53405 6740
rect 55420 6700 64280 6740
rect 70051 6700 70060 6740
rect 70100 6700 75340 6740
rect 75380 6700 75389 6740
rect 81283 6700 81292 6740
rect 81332 6700 83156 6740
rect 83875 6700 83884 6740
rect 83924 6700 88588 6740
rect 88628 6700 88637 6740
rect 16195 6699 16253 6700
rect 23395 6699 23453 6700
rect 24547 6699 24605 6700
rect 48931 6656 48989 6657
rect 3139 6616 3148 6656
rect 3188 6616 15820 6656
rect 15860 6616 15869 6656
rect 15916 6616 18220 6656
rect 18260 6616 23788 6656
rect 23828 6616 23837 6656
rect 25123 6616 25132 6656
rect 25172 6616 27148 6656
rect 27188 6616 31660 6656
rect 31700 6616 31709 6656
rect 31843 6616 31852 6656
rect 31892 6616 34060 6656
rect 34100 6616 38668 6656
rect 38708 6616 38717 6656
rect 40195 6616 40204 6656
rect 40244 6616 48940 6656
rect 48980 6616 48989 6656
rect 49804 6656 49844 6700
rect 64240 6656 64280 6700
rect 71971 6656 72029 6657
rect 76291 6656 76349 6657
rect 77539 6656 77597 6657
rect 80419 6656 80477 6657
rect 83116 6656 83156 6700
rect 84259 6656 84317 6657
rect 49804 6616 59308 6656
rect 59348 6616 60268 6656
rect 60308 6616 61036 6656
rect 61076 6616 61085 6656
rect 64240 6616 68620 6656
rect 68660 6616 68669 6656
rect 71491 6616 71500 6656
rect 71540 6616 71788 6656
rect 71828 6616 71837 6656
rect 71886 6616 71980 6656
rect 72020 6616 72652 6656
rect 72692 6616 72701 6656
rect 73987 6616 73996 6656
rect 74036 6616 74045 6656
rect 74179 6616 74188 6656
rect 74228 6616 76300 6656
rect 76340 6616 76349 6656
rect 77454 6616 77548 6656
rect 77588 6616 77597 6656
rect 78595 6616 78604 6656
rect 78644 6616 79468 6656
rect 79508 6616 79517 6656
rect 80419 6616 80428 6656
rect 80468 6616 82252 6656
rect 82292 6616 82301 6656
rect 83116 6616 84268 6656
rect 84308 6616 84317 6656
rect 15916 6572 15956 6616
rect 25132 6572 25172 6616
rect 31852 6572 31892 6616
rect 48931 6615 48989 6616
rect 71971 6615 72029 6616
rect 35683 6572 35741 6573
rect 38467 6572 38525 6573
rect 56899 6572 56957 6573
rect 57379 6572 57437 6573
rect 60739 6572 60797 6573
rect 66979 6572 67037 6573
rect 67171 6572 67229 6573
rect 73996 6572 74036 6616
rect 76291 6615 76349 6616
rect 77539 6615 77597 6616
rect 80419 6615 80477 6616
rect 84259 6615 84317 6616
rect 79843 6572 79901 6573
rect 82339 6572 82397 6573
rect 10243 6532 10252 6572
rect 10292 6532 10444 6572
rect 10484 6532 10493 6572
rect 12259 6532 12268 6572
rect 12308 6532 15148 6572
rect 15188 6532 15197 6572
rect 15619 6532 15628 6572
rect 15668 6532 15956 6572
rect 16387 6532 16396 6572
rect 16436 6532 16445 6572
rect 18307 6532 18316 6572
rect 18356 6532 19468 6572
rect 19508 6532 19517 6572
rect 19852 6532 25172 6572
rect 26572 6532 31892 6572
rect 32227 6532 32236 6572
rect 32276 6532 34636 6572
rect 34676 6532 34685 6572
rect 35491 6532 35500 6572
rect 35540 6532 35692 6572
rect 35732 6532 35741 6572
rect 37891 6532 37900 6572
rect 37940 6532 38476 6572
rect 38516 6532 38525 6572
rect 16396 6488 16436 6532
rect 19852 6488 19892 6532
rect 26572 6488 26612 6532
rect 35683 6531 35741 6532
rect 38467 6531 38525 6532
rect 38572 6532 43468 6572
rect 43508 6532 43517 6572
rect 44620 6532 47884 6572
rect 47924 6532 47933 6572
rect 51235 6532 51244 6572
rect 51284 6532 52300 6572
rect 52340 6532 52349 6572
rect 55171 6532 55180 6572
rect 55220 6532 56620 6572
rect 56660 6532 56669 6572
rect 56899 6532 56908 6572
rect 56948 6532 57100 6572
rect 57140 6532 57149 6572
rect 57283 6532 57292 6572
rect 57332 6532 57388 6572
rect 57428 6532 57437 6572
rect 60654 6532 60748 6572
rect 60788 6532 61324 6572
rect 61364 6532 61373 6572
rect 61891 6532 61900 6572
rect 61940 6532 66988 6572
rect 67028 6532 67037 6572
rect 67086 6532 67180 6572
rect 67220 6532 67229 6572
rect 68803 6532 68812 6572
rect 68852 6532 69676 6572
rect 69716 6532 74036 6572
rect 74083 6532 74092 6572
rect 74132 6532 76780 6572
rect 76820 6532 77068 6572
rect 77108 6532 77492 6572
rect 77635 6532 77644 6572
rect 77684 6532 78220 6572
rect 78260 6532 78269 6572
rect 79267 6532 79276 6572
rect 79316 6532 79325 6572
rect 79758 6532 79852 6572
rect 79892 6532 79901 6572
rect 82254 6532 82348 6572
rect 82388 6532 82397 6572
rect 83299 6532 83308 6572
rect 83348 6532 85420 6572
rect 85460 6532 85469 6572
rect 86467 6532 86476 6572
rect 86516 6532 87436 6572
rect 87476 6532 87485 6572
rect 38572 6488 38612 6532
rect 1411 6448 1420 6488
rect 1460 6448 10156 6488
rect 10196 6448 10205 6488
rect 10348 6448 11156 6488
rect 12547 6448 12556 6488
rect 12596 6448 16436 6488
rect 17620 6448 18700 6488
rect 18740 6448 19892 6488
rect 23779 6448 23788 6488
rect 23828 6448 26572 6488
rect 26612 6448 26621 6488
rect 27907 6448 27916 6488
rect 27956 6448 27996 6488
rect 28960 6448 29164 6488
rect 29204 6448 33004 6488
rect 33044 6448 33053 6488
rect 33187 6448 33196 6488
rect 33236 6448 36020 6488
rect 37315 6448 37324 6488
rect 37364 6448 37804 6488
rect 37844 6448 37853 6488
rect 37900 6448 38612 6488
rect 38755 6448 38764 6488
rect 38804 6448 44428 6488
rect 44468 6448 44477 6488
rect 10348 6404 10388 6448
rect 11116 6404 11156 6448
rect 17620 6404 17660 6448
rect 19939 6404 19997 6405
rect 27916 6404 27956 6448
rect 28960 6404 29000 6448
rect 30115 6404 30173 6405
rect 35779 6404 35837 6405
rect 35980 6404 36020 6448
rect 37900 6404 37940 6448
rect 44620 6404 44660 6532
rect 56899 6531 56957 6532
rect 57379 6531 57437 6532
rect 60739 6531 60797 6532
rect 66979 6531 67037 6532
rect 67171 6531 67229 6532
rect 55651 6488 55709 6489
rect 77452 6488 77492 6532
rect 79276 6488 79316 6532
rect 79843 6531 79901 6532
rect 82339 6531 82397 6532
rect 81955 6488 82013 6489
rect 82243 6488 82301 6489
rect 44803 6448 44812 6488
rect 44852 6448 45100 6488
rect 45140 6448 47404 6488
rect 47444 6448 47692 6488
rect 47732 6448 50324 6488
rect 50851 6448 50860 6488
rect 50900 6448 51436 6488
rect 51476 6448 52012 6488
rect 52052 6448 52588 6488
rect 52628 6448 52637 6488
rect 53347 6448 53356 6488
rect 53396 6448 55604 6488
rect 45667 6404 45725 6405
rect 2755 6364 2764 6404
rect 2804 6364 10388 6404
rect 10435 6364 10444 6404
rect 10484 6364 10924 6404
rect 10964 6364 10973 6404
rect 11116 6364 11360 6404
rect 13219 6364 13228 6404
rect 13268 6364 15052 6404
rect 15092 6364 15101 6404
rect 15811 6364 15820 6404
rect 15860 6364 16012 6404
rect 16052 6364 16244 6404
rect 16291 6364 16300 6404
rect 16340 6364 17660 6404
rect 19564 6364 19660 6404
rect 19700 6364 19948 6404
rect 19988 6364 19997 6404
rect 22915 6364 22924 6404
rect 22964 6364 23212 6404
rect 23252 6364 23261 6404
rect 23395 6364 23404 6404
rect 23444 6364 23596 6404
rect 23636 6364 24076 6404
rect 24116 6364 25036 6404
rect 25076 6364 25324 6404
rect 25364 6364 25373 6404
rect 25507 6364 25516 6404
rect 25556 6364 26188 6404
rect 26228 6364 26237 6404
rect 26371 6364 26380 6404
rect 26420 6364 26764 6404
rect 26804 6364 26956 6404
rect 26996 6364 27532 6404
rect 27572 6364 28492 6404
rect 28532 6364 28541 6404
rect 28675 6364 28684 6404
rect 28724 6364 29000 6404
rect 30019 6364 30028 6404
rect 30068 6364 30124 6404
rect 30164 6364 30173 6404
rect 32035 6364 32044 6404
rect 32084 6364 32093 6404
rect 32611 6364 32620 6404
rect 32660 6364 33100 6404
rect 33140 6364 33149 6404
rect 33859 6364 33868 6404
rect 33908 6364 34348 6404
rect 34388 6364 35020 6404
rect 35060 6364 35069 6404
rect 35779 6364 35788 6404
rect 35828 6364 35878 6404
rect 35918 6364 35927 6404
rect 35971 6364 35980 6404
rect 36020 6364 36364 6404
rect 36404 6364 36413 6404
rect 36835 6364 36844 6404
rect 36884 6364 37940 6404
rect 38083 6364 38092 6404
rect 38132 6364 39148 6404
rect 39188 6364 39197 6404
rect 41635 6364 41644 6404
rect 41684 6364 44660 6404
rect 44707 6364 44716 6404
rect 44756 6364 44765 6404
rect 45582 6364 45676 6404
rect 45716 6364 45725 6404
rect 48067 6364 48076 6404
rect 48116 6364 49324 6404
rect 49364 6364 49373 6404
rect 11320 6320 11360 6364
rect 16204 6320 16244 6364
rect 19564 6320 19604 6364
rect 19939 6363 19997 6364
rect 19747 6320 19805 6321
rect 25516 6320 25556 6364
rect 30115 6363 30173 6364
rect 32044 6320 32084 6364
rect 35779 6363 35837 6364
rect 32899 6320 32957 6321
rect 33763 6320 33821 6321
rect 34339 6320 34397 6321
rect 36163 6320 36221 6321
rect 37891 6320 37949 6321
rect 6883 6280 6892 6320
rect 6932 6280 11116 6320
rect 11156 6280 11165 6320
rect 11320 6280 16108 6320
rect 16148 6280 16157 6320
rect 16204 6280 16397 6320
rect 16437 6280 17260 6320
rect 17300 6280 19604 6320
rect 19662 6280 19756 6320
rect 19796 6280 19805 6320
rect 19747 6279 19805 6280
rect 20145 6280 25556 6320
rect 26380 6280 27052 6320
rect 27092 6280 27101 6320
rect 27427 6280 27436 6320
rect 27476 6280 29836 6320
rect 29876 6280 29885 6320
rect 31651 6280 31660 6320
rect 31700 6280 32084 6320
rect 32323 6280 32332 6320
rect 32372 6280 32908 6320
rect 32948 6280 32957 6320
rect 20145 6236 20185 6280
rect 26380 6236 26420 6280
rect 32899 6279 32957 6280
rect 33004 6280 33772 6320
rect 33812 6280 33821 6320
rect 34147 6280 34156 6320
rect 34196 6280 34348 6320
rect 34388 6280 34397 6320
rect 33004 6236 33044 6280
rect 33763 6279 33821 6280
rect 34339 6279 34397 6280
rect 34540 6280 36172 6320
rect 36212 6280 36221 6320
rect 37806 6280 37900 6320
rect 37940 6280 37949 6320
rect 38275 6280 38284 6320
rect 38324 6280 38860 6320
rect 38900 6280 38909 6320
rect 34243 6236 34301 6237
rect 34540 6236 34580 6280
rect 36163 6279 36221 6280
rect 37891 6279 37949 6280
rect 37315 6236 37373 6237
rect 44716 6236 44756 6364
rect 45667 6363 45725 6364
rect 50284 6320 50324 6448
rect 54979 6404 55037 6405
rect 55564 6404 55604 6448
rect 55651 6448 55660 6488
rect 55700 6448 57484 6488
rect 57524 6448 57533 6488
rect 57859 6448 57868 6488
rect 57908 6448 64280 6488
rect 64771 6448 64780 6488
rect 64820 6448 66548 6488
rect 66595 6448 66604 6488
rect 66644 6448 69100 6488
rect 69140 6448 74612 6488
rect 74659 6448 74668 6488
rect 74708 6448 75340 6488
rect 75380 6448 75389 6488
rect 77443 6448 77452 6488
rect 77492 6448 77501 6488
rect 77731 6448 77740 6488
rect 77780 6448 78028 6488
rect 78068 6448 78077 6488
rect 78787 6448 78796 6488
rect 78836 6448 78845 6488
rect 79276 6448 80140 6488
rect 80180 6448 80189 6488
rect 80323 6448 80332 6488
rect 80372 6448 81140 6488
rect 55651 6447 55709 6448
rect 60067 6404 60125 6405
rect 64240 6404 64280 6448
rect 66508 6404 66548 6448
rect 69379 6404 69437 6405
rect 74572 6404 74612 6448
rect 78796 6404 78836 6448
rect 50371 6364 50380 6404
rect 50420 6364 50764 6404
rect 50804 6364 50813 6404
rect 51523 6364 51532 6404
rect 51572 6364 51916 6404
rect 51956 6364 51965 6404
rect 52675 6364 52684 6404
rect 52724 6364 54796 6404
rect 54836 6364 54845 6404
rect 54979 6364 54988 6404
rect 55028 6364 55122 6404
rect 55555 6364 55564 6404
rect 55604 6364 55613 6404
rect 56515 6364 56524 6404
rect 56564 6364 57004 6404
rect 57044 6364 57053 6404
rect 57571 6364 57580 6404
rect 57620 6364 58252 6404
rect 58292 6364 58301 6404
rect 58435 6364 58444 6404
rect 58484 6364 58924 6404
rect 58964 6364 58973 6404
rect 59982 6364 60076 6404
rect 60116 6364 60125 6404
rect 60451 6364 60460 6404
rect 60500 6364 61900 6404
rect 61940 6364 61949 6404
rect 62275 6364 62284 6404
rect 62324 6364 62668 6404
rect 62708 6364 63148 6404
rect 63188 6364 63197 6404
rect 64240 6364 65260 6404
rect 65300 6364 65309 6404
rect 66508 6364 67084 6404
rect 67124 6364 67372 6404
rect 67412 6364 67421 6404
rect 67747 6364 67756 6404
rect 67796 6364 68140 6404
rect 68180 6364 68524 6404
rect 68564 6364 68573 6404
rect 69379 6364 69388 6404
rect 69428 6364 71404 6404
rect 71444 6364 71453 6404
rect 71779 6364 71788 6404
rect 71828 6364 74092 6404
rect 74132 6364 74141 6404
rect 74563 6364 74572 6404
rect 74612 6364 78700 6404
rect 78740 6364 78749 6404
rect 78796 6364 80468 6404
rect 54979 6363 55037 6364
rect 60067 6363 60125 6364
rect 69379 6363 69437 6364
rect 57283 6320 57341 6321
rect 57571 6320 57629 6321
rect 60076 6320 60116 6363
rect 71011 6320 71069 6321
rect 71299 6320 71357 6321
rect 71971 6320 72029 6321
rect 73027 6320 73085 6321
rect 77827 6320 77885 6321
rect 79939 6320 79997 6321
rect 80428 6320 80468 6364
rect 81100 6320 81140 6448
rect 81955 6448 81964 6488
rect 82004 6448 82098 6488
rect 82243 6448 82252 6488
rect 82292 6448 82386 6488
rect 83107 6448 83116 6488
rect 83156 6448 83404 6488
rect 83444 6448 83453 6488
rect 83587 6448 83596 6488
rect 83636 6448 83645 6488
rect 85315 6448 85324 6488
rect 85364 6448 98476 6488
rect 98516 6448 98525 6488
rect 81955 6447 82013 6448
rect 82243 6447 82301 6448
rect 82147 6404 82205 6405
rect 83596 6404 83636 6448
rect 82147 6364 82156 6404
rect 82196 6364 82348 6404
rect 82388 6364 82924 6404
rect 82964 6364 82973 6404
rect 83596 6364 87860 6404
rect 82147 6363 82205 6364
rect 82819 6320 82877 6321
rect 83779 6320 83837 6321
rect 5443 6196 5452 6236
rect 5492 6196 12556 6236
rect 12596 6196 12605 6236
rect 15139 6196 15148 6236
rect 15188 6196 15724 6236
rect 15764 6196 15773 6236
rect 18211 6196 18220 6236
rect 18260 6196 18269 6236
rect 18595 6196 18604 6236
rect 18644 6196 18892 6236
rect 18932 6196 19372 6236
rect 19412 6196 19421 6236
rect 19843 6196 19852 6236
rect 19892 6196 20185 6236
rect 20419 6196 20428 6236
rect 20468 6196 21484 6236
rect 21524 6196 21533 6236
rect 24259 6196 24268 6236
rect 24308 6196 24460 6236
rect 24500 6196 24788 6236
rect 26371 6196 26380 6236
rect 26420 6196 26429 6236
rect 26563 6196 26572 6236
rect 26612 6196 31468 6236
rect 31508 6196 33044 6236
rect 33763 6196 33772 6236
rect 33812 6196 34252 6236
rect 34292 6196 34301 6236
rect 34531 6196 34540 6236
rect 34580 6196 34589 6236
rect 37230 6196 37324 6236
rect 37364 6196 37373 6236
rect 14467 6152 14525 6153
rect 18220 6152 18260 6196
rect 19852 6152 19892 6196
rect 24643 6152 24701 6153
rect 4771 6112 4780 6152
rect 4820 6112 7372 6152
rect 7412 6112 7421 6152
rect 8995 6112 9004 6152
rect 9044 6112 13708 6152
rect 13748 6112 13757 6152
rect 14382 6112 14476 6152
rect 14516 6112 14525 6152
rect 14755 6112 14764 6152
rect 14804 6112 18260 6152
rect 19171 6112 19180 6152
rect 19220 6112 19892 6152
rect 24558 6112 24652 6152
rect 24692 6112 24701 6152
rect 14467 6111 14525 6112
rect 24643 6111 24701 6112
rect 23011 6068 23069 6069
rect 24748 6068 24788 6196
rect 34243 6195 34301 6196
rect 37315 6195 37373 6196
rect 37420 6196 44756 6236
rect 46600 6280 50188 6320
rect 50228 6280 50237 6320
rect 50284 6280 51052 6320
rect 51092 6280 51572 6320
rect 52483 6280 52492 6320
rect 52532 6280 52876 6320
rect 52916 6280 53260 6320
rect 53300 6280 53309 6320
rect 54124 6280 54412 6320
rect 54452 6280 54700 6320
rect 54740 6280 54749 6320
rect 56131 6280 56140 6320
rect 56180 6280 56716 6320
rect 56756 6280 57292 6320
rect 57332 6280 57388 6320
rect 57428 6280 57437 6320
rect 57571 6280 57580 6320
rect 57620 6280 59116 6320
rect 59156 6280 59165 6320
rect 60076 6280 60308 6320
rect 60355 6280 60364 6320
rect 60404 6280 60556 6320
rect 60596 6280 61420 6320
rect 61460 6280 62092 6320
rect 62132 6280 64780 6320
rect 64820 6280 64829 6320
rect 64963 6280 64972 6320
rect 65012 6280 68908 6320
rect 68948 6280 68957 6320
rect 70926 6280 71020 6320
rect 71060 6280 71069 6320
rect 71214 6280 71308 6320
rect 71348 6280 71980 6320
rect 72020 6280 72029 6320
rect 72942 6280 73036 6320
rect 73076 6280 73085 6320
rect 74371 6280 74380 6320
rect 74420 6280 74668 6320
rect 74708 6280 75148 6320
rect 75188 6280 75197 6320
rect 77827 6280 77836 6320
rect 77876 6280 78412 6320
rect 78452 6280 78461 6320
rect 79939 6280 79948 6320
rect 79988 6280 80236 6320
rect 80276 6280 80285 6320
rect 80419 6280 80428 6320
rect 80468 6280 80477 6320
rect 81100 6280 82636 6320
rect 82676 6280 82685 6320
rect 82734 6280 82828 6320
rect 82868 6280 82877 6320
rect 83011 6280 83020 6320
rect 83060 6280 83308 6320
rect 83348 6280 83692 6320
rect 83732 6280 83788 6320
rect 83828 6280 83837 6320
rect 83971 6280 83980 6320
rect 84020 6280 84788 6320
rect 84835 6280 84844 6320
rect 84884 6280 86668 6320
rect 86708 6280 87436 6320
rect 87476 6280 87485 6320
rect 32131 6152 32189 6153
rect 34915 6152 34973 6153
rect 37420 6152 37460 6196
rect 30307 6112 30316 6152
rect 30356 6112 32140 6152
rect 32180 6112 32189 6152
rect 32707 6112 32716 6152
rect 32756 6112 34924 6152
rect 34964 6112 34973 6152
rect 37219 6112 37228 6152
rect 37268 6112 37460 6152
rect 37699 6152 37757 6153
rect 41539 6152 41597 6153
rect 45091 6152 45149 6153
rect 46600 6152 46640 6280
rect 51532 6236 51572 6280
rect 54124 6236 54164 6280
rect 57283 6279 57341 6280
rect 57571 6279 57629 6280
rect 56995 6236 57053 6237
rect 57187 6236 57245 6237
rect 58051 6236 58109 6237
rect 51523 6196 51532 6236
rect 51572 6196 51581 6236
rect 54115 6196 54124 6236
rect 54164 6196 54173 6236
rect 54307 6196 54316 6236
rect 54356 6196 54892 6236
rect 54932 6196 54941 6236
rect 55459 6196 55468 6236
rect 55508 6196 56332 6236
rect 56372 6196 56381 6236
rect 56428 6196 57004 6236
rect 57044 6196 57053 6236
rect 57102 6196 57196 6236
rect 57236 6196 57245 6236
rect 57955 6196 57964 6236
rect 58004 6196 58060 6236
rect 58100 6196 58109 6236
rect 60268 6236 60308 6280
rect 71011 6279 71069 6280
rect 71299 6279 71357 6280
rect 71971 6279 72029 6280
rect 73027 6279 73085 6280
rect 77827 6279 77885 6280
rect 79939 6279 79997 6280
rect 82819 6279 82877 6280
rect 83779 6279 83837 6280
rect 71020 6236 71060 6279
rect 72739 6236 72797 6237
rect 74947 6236 75005 6237
rect 60268 6196 61228 6236
rect 61268 6196 61277 6236
rect 68227 6196 68236 6236
rect 68276 6196 69196 6236
rect 69236 6196 69245 6236
rect 69379 6196 69388 6236
rect 69428 6196 70156 6236
rect 70196 6196 70205 6236
rect 71020 6196 71980 6236
rect 72020 6196 72364 6236
rect 72404 6196 72413 6236
rect 72739 6196 72748 6236
rect 72788 6196 72940 6236
rect 72980 6196 72989 6236
rect 73507 6196 73516 6236
rect 73556 6196 73900 6236
rect 73940 6196 73949 6236
rect 74862 6196 74956 6236
rect 74996 6196 75005 6236
rect 55747 6152 55805 6153
rect 56428 6152 56468 6196
rect 56995 6195 57053 6196
rect 57187 6195 57245 6196
rect 58051 6195 58109 6196
rect 72739 6195 72797 6196
rect 74947 6195 75005 6196
rect 76867 6236 76925 6237
rect 76867 6196 76876 6236
rect 76916 6196 77068 6236
rect 77108 6196 77117 6236
rect 78412 6196 79660 6236
rect 79700 6196 81920 6236
rect 81962 6196 81971 6236
rect 82011 6196 84308 6236
rect 76867 6195 76925 6196
rect 57859 6152 57917 6153
rect 78412 6152 78452 6196
rect 81880 6152 81920 6196
rect 37699 6112 37708 6152
rect 37748 6112 41548 6152
rect 41588 6112 41597 6152
rect 45006 6112 45100 6152
rect 45140 6112 45149 6152
rect 46339 6112 46348 6152
rect 46388 6112 46640 6152
rect 50188 6112 52588 6152
rect 52628 6112 52637 6152
rect 53443 6112 53452 6152
rect 53492 6112 55372 6152
rect 55412 6112 55421 6152
rect 55651 6112 55660 6152
rect 55700 6112 55756 6152
rect 55796 6112 55805 6152
rect 32131 6111 32189 6112
rect 34915 6111 34973 6112
rect 37699 6111 37757 6112
rect 41539 6111 41597 6112
rect 45091 6111 45149 6112
rect 38179 6068 38237 6069
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 16003 6028 16012 6068
rect 16052 6028 16684 6068
rect 16724 6028 19084 6068
rect 19124 6028 19133 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 22926 6028 23020 6068
rect 23060 6028 23069 6068
rect 23011 6027 23069 6028
rect 23116 6028 23308 6068
rect 23348 6028 23357 6068
rect 24739 6028 24748 6068
rect 24788 6028 24797 6068
rect 27715 6028 27724 6068
rect 27764 6028 31852 6068
rect 31892 6028 31901 6068
rect 32332 6028 34732 6068
rect 34772 6028 34781 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 35596 6028 37900 6068
rect 37940 6028 37949 6068
rect 38094 6028 38188 6068
rect 38228 6028 38237 6068
rect 23116 5984 23156 6028
rect 24547 5984 24605 5985
rect 32332 5984 32372 6028
rect 34732 5984 34772 6028
rect 35596 5984 35636 6028
rect 38179 6027 38237 6028
rect 38467 6068 38525 6069
rect 50188 6068 50228 6112
rect 55747 6111 55805 6112
rect 56044 6112 56468 6152
rect 56611 6112 56620 6152
rect 56660 6112 57868 6152
rect 57908 6112 57917 6152
rect 59587 6112 59596 6152
rect 59636 6112 60364 6152
rect 60404 6112 60413 6152
rect 65059 6112 65068 6152
rect 65108 6112 68716 6152
rect 68756 6112 68765 6152
rect 68899 6112 68908 6152
rect 68948 6112 73652 6152
rect 75331 6112 75340 6152
rect 75380 6112 78452 6152
rect 78499 6112 78508 6152
rect 78548 6112 78796 6152
rect 78836 6112 78845 6152
rect 81880 6112 83308 6152
rect 83348 6112 83500 6152
rect 83540 6112 83884 6152
rect 83924 6112 83933 6152
rect 56044 6068 56084 6112
rect 57859 6111 57917 6112
rect 38467 6028 38476 6068
rect 38516 6028 38956 6068
rect 38996 6028 39005 6068
rect 44323 6028 44332 6068
rect 44372 6028 50228 6068
rect 50279 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50665 6068
rect 55267 6028 55276 6068
rect 55316 6028 56084 6068
rect 56131 6028 56140 6068
rect 56180 6028 57676 6068
rect 57716 6028 57725 6068
rect 65399 6028 65408 6068
rect 65448 6028 65490 6068
rect 65530 6028 65572 6068
rect 65612 6028 65654 6068
rect 65694 6028 65736 6068
rect 65776 6028 65785 6068
rect 65836 6028 70636 6068
rect 70676 6028 70685 6068
rect 72748 6028 73228 6068
rect 73268 6028 73277 6068
rect 38467 6027 38525 6028
rect 15907 5944 15916 5984
rect 15956 5944 16396 5984
rect 16436 5944 16445 5984
rect 17059 5944 17068 5984
rect 17108 5944 17452 5984
rect 17492 5944 18316 5984
rect 18356 5944 22924 5984
rect 22964 5944 22973 5984
rect 23107 5944 23116 5984
rect 23156 5944 23165 5984
rect 23308 5944 24556 5984
rect 24596 5944 24605 5984
rect 26179 5944 26188 5984
rect 26228 5944 32332 5984
rect 32372 5944 32381 5984
rect 33379 5944 33388 5984
rect 33428 5944 33772 5984
rect 33812 5944 33821 5984
rect 34732 5944 35636 5984
rect 36163 5984 36221 5985
rect 60259 5984 60317 5985
rect 65836 5984 65876 6028
rect 68323 5984 68381 5985
rect 72748 5984 72788 6028
rect 72931 5984 72989 5985
rect 73612 5984 73652 6112
rect 73795 6068 73853 6069
rect 73795 6028 73804 6068
rect 73844 6028 73938 6068
rect 73987 6028 73996 6068
rect 74036 6028 78412 6068
rect 78452 6028 78461 6068
rect 78883 6028 78892 6068
rect 78932 6028 79084 6068
rect 79124 6028 79133 6068
rect 79363 6028 79372 6068
rect 79412 6028 80044 6068
rect 80084 6028 80093 6068
rect 80519 6028 80528 6068
rect 80568 6028 80610 6068
rect 80650 6028 80692 6068
rect 80732 6028 80774 6068
rect 80814 6028 80856 6068
rect 80896 6028 80905 6068
rect 81091 6028 81100 6068
rect 81140 6028 81964 6068
rect 82004 6028 82013 6068
rect 82156 6028 84172 6068
rect 84212 6028 84221 6068
rect 73795 6027 73853 6028
rect 81667 5984 81725 5985
rect 82156 5984 82196 6028
rect 82531 5984 82589 5985
rect 36163 5944 36172 5984
rect 36212 5944 41260 5984
rect 41300 5944 41309 5984
rect 41356 5944 45676 5984
rect 45716 5944 45725 5984
rect 45955 5944 45964 5984
rect 46004 5944 46828 5984
rect 46868 5944 47020 5984
rect 47060 5944 47069 5984
rect 47875 5944 47884 5984
rect 47924 5944 48404 5984
rect 53731 5944 53740 5984
rect 53780 5944 53932 5984
rect 53972 5944 53981 5984
rect 54595 5944 54604 5984
rect 54644 5944 59116 5984
rect 59156 5944 59165 5984
rect 60259 5944 60268 5984
rect 60308 5944 61324 5984
rect 61364 5944 61804 5984
rect 61844 5944 61996 5984
rect 62036 5944 62045 5984
rect 65251 5944 65260 5984
rect 65300 5944 65876 5984
rect 68238 5944 68332 5984
rect 68372 5944 68381 5984
rect 68707 5944 68716 5984
rect 68756 5944 70100 5984
rect 71491 5944 71500 5984
rect 71540 5944 72748 5984
rect 72788 5944 72797 5984
rect 72931 5944 72940 5984
rect 72980 5944 73516 5984
rect 73556 5944 73565 5984
rect 73612 5944 73900 5984
rect 73940 5944 78508 5984
rect 78548 5944 81676 5984
rect 81716 5944 81725 5984
rect 19171 5900 19229 5901
rect 23308 5900 23348 5944
rect 24547 5943 24605 5944
rect 36163 5943 36221 5944
rect 23875 5900 23933 5901
rect 24556 5900 24596 5943
rect 26947 5900 27005 5901
rect 30019 5900 30077 5901
rect 33091 5900 33149 5901
rect 34435 5900 34493 5901
rect 36067 5900 36125 5901
rect 9667 5860 9676 5900
rect 9716 5860 16972 5900
rect 17012 5860 17021 5900
rect 17155 5860 17164 5900
rect 17204 5860 19180 5900
rect 19220 5860 19229 5900
rect 19555 5860 19564 5900
rect 19604 5860 19948 5900
rect 19988 5860 23348 5900
rect 23395 5860 23404 5900
rect 23444 5860 23692 5900
rect 23732 5860 23741 5900
rect 23875 5860 23884 5900
rect 23924 5860 23980 5900
rect 24020 5860 24029 5900
rect 24556 5860 26572 5900
rect 26612 5860 26621 5900
rect 26862 5860 26956 5900
rect 26996 5860 27005 5900
rect 28099 5860 28108 5900
rect 28148 5860 30028 5900
rect 30068 5860 30077 5900
rect 30307 5860 30316 5900
rect 30356 5860 30892 5900
rect 30932 5860 31084 5900
rect 31124 5860 31133 5900
rect 33006 5860 33100 5900
rect 33140 5860 34156 5900
rect 34196 5860 34444 5900
rect 34484 5860 34493 5900
rect 35587 5860 35596 5900
rect 35636 5860 36076 5900
rect 36116 5860 36125 5900
rect 19171 5859 19229 5860
rect 23875 5859 23933 5860
rect 26947 5859 27005 5860
rect 30019 5859 30077 5860
rect 33091 5859 33149 5860
rect 34435 5859 34493 5860
rect 36067 5859 36125 5860
rect 36172 5860 39148 5900
rect 39188 5860 39197 5900
rect 31267 5816 31325 5817
rect 36172 5816 36212 5860
rect 41356 5816 41396 5944
rect 48364 5900 48404 5944
rect 60259 5943 60317 5944
rect 68323 5943 68381 5944
rect 61987 5900 62045 5901
rect 70060 5900 70100 5944
rect 72931 5943 72989 5944
rect 81667 5943 81725 5944
rect 82060 5944 82196 5984
rect 82446 5944 82540 5984
rect 82580 5944 82589 5984
rect 83107 5944 83116 5984
rect 83156 5944 84076 5984
rect 84116 5944 84125 5984
rect 82060 5900 82100 5944
rect 82531 5943 82589 5944
rect 83875 5900 83933 5901
rect 84268 5900 84308 6196
rect 84748 5984 84788 6280
rect 87820 6236 87860 6364
rect 89539 6280 89548 6320
rect 89588 6280 90892 6320
rect 90932 6280 90941 6320
rect 87811 6196 87820 6236
rect 87860 6196 87869 6236
rect 95639 6028 95648 6068
rect 95688 6028 95730 6068
rect 95770 6028 95812 6068
rect 95852 6028 95894 6068
rect 95934 6028 95976 6068
rect 96016 6028 96025 6068
rect 84748 5944 93484 5984
rect 93524 5944 93533 5984
rect 44131 5860 44140 5900
rect 44180 5860 48268 5900
rect 48308 5860 48317 5900
rect 48364 5860 56140 5900
rect 56180 5860 56189 5900
rect 56323 5860 56332 5900
rect 56372 5860 56524 5900
rect 56564 5860 56573 5900
rect 56803 5860 56812 5900
rect 56852 5860 61996 5900
rect 62036 5860 62045 5900
rect 63907 5860 63916 5900
rect 63956 5860 69964 5900
rect 70004 5860 70013 5900
rect 70060 5860 71692 5900
rect 71732 5860 71741 5900
rect 72067 5860 72076 5900
rect 72116 5860 76684 5900
rect 76724 5860 76733 5900
rect 78883 5860 78892 5900
rect 78932 5860 80908 5900
rect 80948 5860 80957 5900
rect 81379 5860 81388 5900
rect 81428 5860 82100 5900
rect 82147 5860 82156 5900
rect 82196 5860 82924 5900
rect 82964 5860 83692 5900
rect 83732 5860 83741 5900
rect 83875 5860 83884 5900
rect 83924 5860 83964 5900
rect 84268 5860 85132 5900
rect 85172 5860 85181 5900
rect 55843 5816 55901 5817
rect 56524 5816 56564 5860
rect 61987 5859 62045 5860
rect 83875 5859 83933 5860
rect 57475 5816 57533 5817
rect 67843 5816 67901 5817
rect 72931 5816 72989 5817
rect 83884 5816 83924 5859
rect 15331 5776 15340 5816
rect 15380 5776 16108 5816
rect 16148 5776 16876 5816
rect 16916 5776 19084 5816
rect 19124 5776 19756 5816
rect 19796 5776 20276 5816
rect 20323 5776 20332 5816
rect 20372 5776 20716 5816
rect 20756 5776 24020 5816
rect 15619 5732 15677 5733
rect 4099 5692 4108 5732
rect 4148 5692 15628 5732
rect 15668 5692 15677 5732
rect 15619 5691 15677 5692
rect 1699 5648 1757 5649
rect 15724 5648 15764 5776
rect 15811 5732 15869 5733
rect 20236 5732 20276 5776
rect 23299 5732 23357 5733
rect 23980 5732 24020 5776
rect 30028 5776 30740 5816
rect 31182 5776 31276 5816
rect 31316 5776 31325 5816
rect 31843 5776 31852 5816
rect 31892 5776 34540 5816
rect 34580 5776 36212 5816
rect 37027 5776 37036 5816
rect 37076 5776 37085 5816
rect 37507 5776 37516 5816
rect 37556 5776 41396 5816
rect 44323 5776 44332 5816
rect 44372 5776 44716 5816
rect 44756 5776 45196 5816
rect 45236 5776 46060 5816
rect 46100 5776 46109 5816
rect 50947 5776 50956 5816
rect 50996 5776 55700 5816
rect 15811 5692 15820 5732
rect 15860 5692 15869 5732
rect 16483 5692 16492 5732
rect 16532 5692 17260 5732
rect 17300 5692 17309 5732
rect 18115 5692 18124 5732
rect 18164 5692 18604 5732
rect 18644 5692 18653 5732
rect 18787 5692 18796 5732
rect 18836 5692 19180 5732
rect 19220 5692 19229 5732
rect 20236 5692 20524 5732
rect 20564 5692 20573 5732
rect 23214 5692 23308 5732
rect 23348 5692 23357 5732
rect 23971 5692 23980 5732
rect 24020 5692 27724 5732
rect 27764 5692 27773 5732
rect 28483 5692 28492 5732
rect 28532 5692 28780 5732
rect 28820 5692 28972 5732
rect 29012 5692 29021 5732
rect 15811 5691 15869 5692
rect 23299 5691 23357 5692
rect 15820 5648 15860 5691
rect 30028 5648 30068 5776
rect 30115 5692 30124 5732
rect 30164 5692 30604 5732
rect 30644 5692 30653 5732
rect 30700 5648 30740 5776
rect 31267 5775 31325 5776
rect 30787 5692 30796 5732
rect 30836 5692 31660 5732
rect 31700 5692 32044 5732
rect 32084 5692 32428 5732
rect 32468 5692 32812 5732
rect 32852 5692 32861 5732
rect 34339 5692 34348 5732
rect 34388 5692 34732 5732
rect 34772 5692 35404 5732
rect 35444 5692 35453 5732
rect 36259 5692 36268 5732
rect 36308 5692 36556 5732
rect 36596 5692 36605 5732
rect 34915 5648 34973 5649
rect 1614 5608 1708 5648
rect 1748 5608 1757 5648
rect 2083 5608 2092 5648
rect 2132 5608 9580 5648
rect 9620 5608 9629 5648
rect 15715 5608 15724 5648
rect 15764 5608 15773 5648
rect 15820 5608 20236 5648
rect 20276 5608 20285 5648
rect 27619 5608 27628 5648
rect 27668 5608 30068 5648
rect 30403 5608 30412 5648
rect 30452 5608 30461 5648
rect 30700 5608 32524 5648
rect 32564 5608 32573 5648
rect 34830 5608 34924 5648
rect 34964 5608 34973 5648
rect 1699 5607 1757 5608
rect 19939 5564 19997 5565
rect 30412 5564 30452 5608
rect 34915 5607 34973 5608
rect 35971 5648 36029 5649
rect 37036 5648 37076 5776
rect 37699 5692 37708 5732
rect 37748 5692 38572 5732
rect 38612 5692 38621 5732
rect 38755 5692 38764 5732
rect 38804 5692 38813 5732
rect 39139 5692 39148 5732
rect 39188 5692 40780 5732
rect 40820 5692 40829 5732
rect 41560 5692 48652 5732
rect 48692 5692 48701 5732
rect 49603 5692 49612 5732
rect 49652 5692 51436 5732
rect 51476 5692 51485 5732
rect 53923 5692 53932 5732
rect 53972 5692 54316 5732
rect 54356 5692 54365 5732
rect 54499 5692 54508 5732
rect 54548 5692 54988 5732
rect 55028 5692 55037 5732
rect 38764 5648 38804 5692
rect 35971 5608 35980 5648
rect 36020 5608 36460 5648
rect 36500 5608 36509 5648
rect 37036 5608 38092 5648
rect 38132 5608 39052 5648
rect 39092 5608 39340 5648
rect 39380 5608 39389 5648
rect 35971 5607 36029 5608
rect 33763 5564 33821 5565
rect 41560 5564 41600 5692
rect 43651 5648 43709 5649
rect 55660 5648 55700 5776
rect 55843 5776 55852 5816
rect 55892 5776 55986 5816
rect 56524 5776 57484 5816
rect 57524 5776 57676 5816
rect 57716 5776 57725 5816
rect 67758 5776 67852 5816
rect 67892 5776 67901 5816
rect 55843 5775 55901 5776
rect 57475 5775 57533 5776
rect 67843 5775 67901 5776
rect 67948 5776 69388 5816
rect 69428 5776 69437 5816
rect 70147 5776 70156 5816
rect 70196 5776 72940 5816
rect 72980 5776 72989 5816
rect 58243 5732 58301 5733
rect 61219 5732 61277 5733
rect 64579 5732 64637 5733
rect 67948 5732 67988 5776
rect 72931 5775 72989 5776
rect 73420 5776 74284 5816
rect 74324 5776 80236 5816
rect 80276 5776 80812 5816
rect 80852 5776 80861 5816
rect 81484 5776 82348 5816
rect 82388 5776 82828 5816
rect 82868 5776 82877 5816
rect 82924 5776 83828 5816
rect 83875 5776 83884 5816
rect 83924 5776 85516 5816
rect 85556 5776 85565 5816
rect 86563 5776 86572 5816
rect 86612 5776 96076 5816
rect 96116 5776 96125 5816
rect 73420 5732 73460 5776
rect 76579 5732 76637 5733
rect 81484 5732 81524 5776
rect 81859 5732 81917 5733
rect 82924 5732 82964 5776
rect 83788 5732 83828 5776
rect 84355 5732 84413 5733
rect 55747 5692 55756 5732
rect 55796 5692 56908 5732
rect 56948 5692 57388 5732
rect 57428 5692 58252 5732
rect 58292 5692 58301 5732
rect 61134 5692 61228 5732
rect 61268 5692 61277 5732
rect 64494 5692 64588 5732
rect 64628 5692 64637 5732
rect 66403 5692 66412 5732
rect 66452 5692 67988 5732
rect 68035 5692 68044 5732
rect 68084 5692 68332 5732
rect 68372 5692 68381 5732
rect 69763 5692 69772 5732
rect 69812 5692 71308 5732
rect 71348 5692 71357 5732
rect 71404 5692 73420 5732
rect 73460 5692 73469 5732
rect 73603 5692 73612 5732
rect 73652 5692 73996 5732
rect 74036 5692 74045 5732
rect 74467 5692 74476 5732
rect 74516 5692 74668 5732
rect 74708 5692 74956 5732
rect 74996 5692 75005 5732
rect 75235 5692 75244 5732
rect 75284 5692 76588 5732
rect 76628 5692 76637 5732
rect 78403 5692 78412 5732
rect 78452 5692 78461 5732
rect 78787 5692 78796 5732
rect 78836 5692 79084 5732
rect 79124 5692 79468 5732
rect 79508 5692 79852 5732
rect 79892 5692 80044 5732
rect 80084 5692 80093 5732
rect 80419 5692 80428 5732
rect 80468 5692 80908 5732
rect 80948 5692 81292 5732
rect 81332 5692 81341 5732
rect 81475 5692 81484 5732
rect 81524 5692 81533 5732
rect 81859 5692 81868 5732
rect 81908 5692 82964 5732
rect 83779 5692 83788 5732
rect 83828 5692 83837 5732
rect 84270 5692 84364 5732
rect 84404 5692 84413 5732
rect 58243 5691 58301 5692
rect 61219 5691 61277 5692
rect 64579 5691 64637 5692
rect 56707 5648 56765 5649
rect 66787 5648 66845 5649
rect 71404 5648 71444 5692
rect 76579 5691 76637 5692
rect 78412 5648 78452 5692
rect 81859 5691 81917 5692
rect 84355 5691 84413 5692
rect 88387 5732 88445 5733
rect 88387 5692 88396 5732
rect 88436 5692 96268 5732
rect 96308 5692 96317 5732
rect 88387 5691 88445 5692
rect 81763 5648 81821 5649
rect 82147 5648 82205 5649
rect 97507 5648 97565 5649
rect 14284 5524 17260 5564
rect 17300 5524 17309 5564
rect 17356 5524 19756 5564
rect 19796 5524 19805 5564
rect 19939 5524 19948 5564
rect 19988 5524 20140 5564
rect 20180 5524 22732 5564
rect 22772 5524 30452 5564
rect 30499 5524 30508 5564
rect 30548 5524 32276 5564
rect 32323 5524 32332 5564
rect 32372 5524 32620 5564
rect 32660 5524 32669 5564
rect 33763 5524 33772 5564
rect 33812 5524 37516 5564
rect 37556 5524 37565 5564
rect 38476 5524 41600 5564
rect 41644 5608 43276 5648
rect 43316 5608 43325 5648
rect 43566 5608 43660 5648
rect 43700 5608 43709 5648
rect 45283 5608 45292 5648
rect 45332 5608 47884 5648
rect 47924 5608 47933 5648
rect 54883 5608 54892 5648
rect 54932 5608 55460 5648
rect 55660 5608 56660 5648
rect 14284 5480 14324 5524
rect 17356 5480 17396 5524
rect 19939 5523 19997 5524
rect 1123 5440 1132 5480
rect 1172 5440 1900 5480
rect 1940 5440 1949 5480
rect 3331 5440 3340 5480
rect 3380 5440 14324 5480
rect 16483 5440 16492 5480
rect 16532 5440 16541 5480
rect 16588 5440 17396 5480
rect 18691 5480 18749 5481
rect 20611 5480 20669 5481
rect 18691 5440 18700 5480
rect 18740 5440 18892 5480
rect 18932 5440 18941 5480
rect 19075 5440 19084 5480
rect 19124 5440 19508 5480
rect 19555 5440 19564 5480
rect 19604 5440 20332 5480
rect 20372 5440 20381 5480
rect 20515 5440 20524 5480
rect 20564 5440 20620 5480
rect 20660 5440 20669 5480
rect 16492 5396 16532 5440
rect 7363 5356 7372 5396
rect 7412 5356 16532 5396
rect 16588 5312 16628 5440
rect 18691 5439 18749 5440
rect 19468 5397 19508 5440
rect 20611 5439 20669 5440
rect 21571 5480 21629 5481
rect 32236 5480 32276 5524
rect 33763 5523 33821 5524
rect 33667 5480 33725 5481
rect 36547 5480 36605 5481
rect 37315 5480 37373 5481
rect 37699 5480 37757 5481
rect 38476 5480 38516 5524
rect 41644 5480 41684 5608
rect 43651 5607 43709 5608
rect 21571 5440 21580 5480
rect 21620 5440 23788 5480
rect 23828 5440 23837 5480
rect 27235 5440 27244 5480
rect 27284 5440 28492 5480
rect 28532 5440 28541 5480
rect 30403 5440 30412 5480
rect 30452 5440 31084 5480
rect 31124 5440 31133 5480
rect 31651 5440 31660 5480
rect 31700 5440 31948 5480
rect 31988 5440 31997 5480
rect 32227 5440 32236 5480
rect 32276 5440 32285 5480
rect 32419 5440 32428 5480
rect 32468 5440 33292 5480
rect 33332 5440 33341 5480
rect 33667 5440 33676 5480
rect 33716 5440 33964 5480
rect 34004 5440 34013 5480
rect 34339 5440 34348 5480
rect 34388 5440 36556 5480
rect 36596 5440 36605 5480
rect 37230 5440 37324 5480
rect 37364 5440 37373 5480
rect 37614 5440 37708 5480
rect 37748 5440 37757 5480
rect 37891 5440 37900 5480
rect 37940 5440 38516 5480
rect 38563 5440 38572 5480
rect 38612 5440 41684 5480
rect 41731 5480 41789 5481
rect 55420 5480 55460 5608
rect 55651 5564 55709 5565
rect 56515 5564 56573 5565
rect 55566 5524 55660 5564
rect 55700 5524 55709 5564
rect 56430 5524 56524 5564
rect 56564 5524 56573 5564
rect 56620 5564 56660 5608
rect 56707 5608 56716 5648
rect 56756 5608 60652 5648
rect 60692 5608 60701 5648
rect 61123 5608 61132 5648
rect 61172 5608 63532 5648
rect 63572 5608 63581 5648
rect 64003 5608 64012 5648
rect 64052 5608 66796 5648
rect 66836 5608 66845 5648
rect 66979 5608 66988 5648
rect 67028 5608 68140 5648
rect 68180 5608 68189 5648
rect 68899 5608 68908 5648
rect 68948 5608 71444 5648
rect 71683 5608 71692 5648
rect 71732 5608 73228 5648
rect 73268 5608 73277 5648
rect 73507 5608 73516 5648
rect 73556 5608 75532 5648
rect 75572 5608 75581 5648
rect 75628 5608 76876 5648
rect 76916 5608 76925 5648
rect 77059 5608 77068 5648
rect 77108 5608 78316 5648
rect 78356 5608 78365 5648
rect 78412 5608 79276 5648
rect 79316 5608 80564 5648
rect 80611 5608 80620 5648
rect 80660 5608 81388 5648
rect 81428 5608 81772 5648
rect 81812 5608 81868 5648
rect 81908 5608 82156 5648
rect 82196 5608 82205 5648
rect 82627 5608 82636 5648
rect 82676 5608 86188 5648
rect 86228 5608 86237 5648
rect 97422 5608 97516 5648
rect 97556 5608 97565 5648
rect 56707 5607 56765 5608
rect 66787 5607 66845 5608
rect 57667 5564 57725 5565
rect 60451 5564 60509 5565
rect 68908 5564 68948 5608
rect 74467 5564 74525 5565
rect 75043 5564 75101 5565
rect 56620 5524 57676 5564
rect 57716 5524 57725 5564
rect 57859 5524 57868 5564
rect 57908 5524 60268 5564
rect 60308 5524 60317 5564
rect 60451 5524 60460 5564
rect 60500 5524 61900 5564
rect 61940 5524 62956 5564
rect 62996 5524 63005 5564
rect 63244 5524 65396 5564
rect 65443 5524 65452 5564
rect 65492 5524 68948 5564
rect 69571 5524 69580 5564
rect 69620 5524 72748 5564
rect 72788 5524 73100 5564
rect 74382 5524 74476 5564
rect 74516 5524 74525 5564
rect 74958 5524 75052 5564
rect 75092 5524 75101 5564
rect 55651 5523 55709 5524
rect 56515 5523 56573 5524
rect 57667 5523 57725 5524
rect 60451 5523 60509 5524
rect 58243 5480 58301 5481
rect 61891 5480 61949 5481
rect 63244 5480 63284 5524
rect 41731 5440 41740 5480
rect 41780 5440 41874 5480
rect 44035 5440 44044 5480
rect 44084 5440 44620 5480
rect 44660 5440 45388 5480
rect 45428 5440 45868 5480
rect 45908 5440 45917 5480
rect 55420 5440 57620 5480
rect 58158 5440 58252 5480
rect 58292 5440 58301 5480
rect 59779 5440 59788 5480
rect 59828 5440 60076 5480
rect 60116 5440 60125 5480
rect 61891 5440 61900 5480
rect 61940 5440 62668 5480
rect 62708 5440 62717 5480
rect 63235 5440 63244 5480
rect 63284 5440 63293 5480
rect 21571 5439 21629 5440
rect 33667 5439 33725 5440
rect 36547 5439 36605 5440
rect 37315 5439 37373 5440
rect 37699 5439 37757 5440
rect 41731 5439 41789 5440
rect 17347 5396 17405 5397
rect 19459 5396 19517 5397
rect 17155 5356 17164 5396
rect 17204 5356 17356 5396
rect 17396 5356 17740 5396
rect 17780 5356 18508 5396
rect 18548 5356 19412 5396
rect 17347 5355 17405 5356
rect 19372 5312 19412 5356
rect 19459 5356 19468 5396
rect 19508 5356 19517 5396
rect 19459 5355 19517 5356
rect 20707 5396 20765 5397
rect 39907 5396 39965 5397
rect 41059 5396 41117 5397
rect 52195 5396 52253 5397
rect 56131 5396 56189 5397
rect 20707 5356 20716 5396
rect 20756 5356 25036 5396
rect 25076 5356 25085 5396
rect 31843 5356 31852 5396
rect 31892 5356 34964 5396
rect 35299 5356 35308 5396
rect 35348 5356 39724 5396
rect 39764 5356 39773 5396
rect 39907 5356 39916 5396
rect 39956 5356 41068 5396
rect 41108 5356 41117 5396
rect 42595 5356 42604 5396
rect 42644 5356 52204 5396
rect 52244 5356 52253 5396
rect 20707 5355 20765 5356
rect 22915 5312 22973 5313
rect 28387 5312 28445 5313
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 8899 5272 8908 5312
rect 8948 5272 16108 5312
rect 16148 5272 16157 5312
rect 16204 5272 16628 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19372 5272 20716 5312
rect 20756 5272 20765 5312
rect 22830 5272 22924 5312
rect 22964 5272 22973 5312
rect 27811 5272 27820 5312
rect 27860 5272 28108 5312
rect 28148 5272 28157 5312
rect 28302 5272 28396 5312
rect 28436 5272 28445 5312
rect 16204 5228 16244 5272
rect 22915 5271 22973 5272
rect 28387 5271 28445 5272
rect 28579 5312 28637 5313
rect 31852 5312 31892 5356
rect 34924 5312 34964 5356
rect 39907 5355 39965 5356
rect 41059 5355 41117 5356
rect 52195 5355 52253 5356
rect 52300 5356 56140 5396
rect 56180 5356 56189 5396
rect 49891 5312 49949 5313
rect 52300 5312 52340 5356
rect 56131 5355 56189 5356
rect 57283 5312 57341 5313
rect 57580 5312 57620 5440
rect 58243 5439 58301 5440
rect 61891 5439 61949 5440
rect 57667 5396 57725 5397
rect 61699 5396 61757 5397
rect 57667 5356 57676 5396
rect 57716 5356 61708 5396
rect 61748 5356 61996 5396
rect 62036 5356 62764 5396
rect 62804 5356 62813 5396
rect 57667 5355 57725 5356
rect 61699 5355 61757 5356
rect 58147 5312 58205 5313
rect 65356 5312 65396 5524
rect 71971 5480 72029 5481
rect 72547 5480 72605 5481
rect 72931 5480 72989 5481
rect 66499 5440 66508 5480
rect 66548 5440 68332 5480
rect 68372 5440 68381 5480
rect 69379 5440 69388 5480
rect 69428 5440 69964 5480
rect 70004 5440 70013 5480
rect 70531 5440 70540 5480
rect 70580 5440 70924 5480
rect 70964 5440 70973 5480
rect 71971 5440 71980 5480
rect 72020 5440 72364 5480
rect 72404 5440 72413 5480
rect 72462 5440 72556 5480
rect 72596 5440 72605 5480
rect 72846 5440 72940 5480
rect 72980 5440 72989 5480
rect 73060 5480 73100 5524
rect 74467 5523 74525 5524
rect 75043 5523 75101 5524
rect 73060 5440 74516 5480
rect 71971 5439 72029 5440
rect 72547 5439 72605 5440
rect 72931 5439 72989 5440
rect 70339 5396 70397 5397
rect 70819 5396 70877 5397
rect 72643 5396 72701 5397
rect 69283 5356 69292 5396
rect 69332 5356 70060 5396
rect 70100 5356 70109 5396
rect 70339 5356 70348 5396
rect 70388 5356 70636 5396
rect 70676 5356 70685 5396
rect 70734 5356 70828 5396
rect 70868 5356 70877 5396
rect 71491 5356 71500 5396
rect 71540 5356 71980 5396
rect 72020 5356 72029 5396
rect 72558 5356 72652 5396
rect 72692 5356 72701 5396
rect 73219 5356 73228 5396
rect 73268 5356 74188 5396
rect 74228 5356 74237 5396
rect 70339 5355 70397 5356
rect 70819 5355 70877 5356
rect 72643 5355 72701 5356
rect 74476 5312 74516 5440
rect 75628 5312 75668 5608
rect 80131 5564 80189 5565
rect 75907 5524 75916 5564
rect 75956 5524 80140 5564
rect 80180 5524 80189 5564
rect 80524 5564 80564 5608
rect 81763 5607 81821 5608
rect 82147 5607 82205 5608
rect 97507 5607 97565 5608
rect 80524 5524 81236 5564
rect 80131 5523 80189 5524
rect 75907 5480 75965 5481
rect 77827 5480 77885 5481
rect 79747 5480 79805 5481
rect 80611 5480 80669 5481
rect 75907 5440 75916 5480
rect 75956 5440 76108 5480
rect 76148 5440 76157 5480
rect 77443 5440 77452 5480
rect 77492 5440 77501 5480
rect 77742 5440 77836 5480
rect 77876 5440 77885 5480
rect 78019 5440 78028 5480
rect 78068 5440 78412 5480
rect 78452 5440 78461 5480
rect 78691 5440 78700 5480
rect 78740 5440 78749 5480
rect 79662 5440 79756 5480
rect 79796 5440 79805 5480
rect 80526 5440 80620 5480
rect 80660 5440 80669 5480
rect 81196 5480 81236 5524
rect 81676 5524 82156 5564
rect 82196 5524 82540 5564
rect 82580 5524 82589 5564
rect 83875 5524 83884 5564
rect 83924 5524 85804 5564
rect 85844 5524 85853 5564
rect 81676 5480 81716 5524
rect 81859 5480 81917 5481
rect 81196 5440 81676 5480
rect 81716 5440 81725 5480
rect 81774 5440 81868 5480
rect 81908 5440 81917 5480
rect 82339 5440 82348 5480
rect 82388 5440 82397 5480
rect 83491 5440 83500 5480
rect 83540 5440 98476 5480
rect 98516 5440 98525 5480
rect 75907 5439 75965 5440
rect 76387 5356 76396 5396
rect 76436 5356 77356 5396
rect 77396 5356 77405 5396
rect 28579 5272 28588 5312
rect 28628 5272 28684 5312
rect 28724 5272 28733 5312
rect 29443 5272 29452 5312
rect 29492 5272 31892 5312
rect 32803 5272 32812 5312
rect 32852 5272 33484 5312
rect 33524 5272 33533 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 34915 5272 34924 5312
rect 34964 5272 35636 5312
rect 38083 5272 38092 5312
rect 38132 5272 45676 5312
rect 45716 5272 45725 5312
rect 49039 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49425 5312
rect 49891 5272 49900 5312
rect 49940 5272 52340 5312
rect 55363 5272 55372 5312
rect 55412 5272 57236 5312
rect 28579 5271 28637 5272
rect 20803 5228 20861 5229
rect 23971 5228 24029 5229
rect 24355 5228 24413 5229
rect 35596 5228 35636 5272
rect 49891 5271 49949 5272
rect 40291 5228 40349 5229
rect 41635 5228 41693 5229
rect 56611 5228 56669 5229
rect 57091 5228 57149 5229
rect 9187 5188 9196 5228
rect 9236 5188 9580 5228
rect 9620 5188 9629 5228
rect 11587 5188 11596 5228
rect 11636 5188 16244 5228
rect 16291 5188 16300 5228
rect 16340 5188 19372 5228
rect 19412 5188 19421 5228
rect 20803 5188 20812 5228
rect 20852 5188 20908 5228
rect 20948 5188 20957 5228
rect 21379 5188 21388 5228
rect 21428 5188 23980 5228
rect 24020 5188 24029 5228
rect 24270 5188 24364 5228
rect 24404 5188 24413 5228
rect 25123 5188 25132 5228
rect 25172 5188 28972 5228
rect 29012 5188 30604 5228
rect 30644 5188 35404 5228
rect 35444 5188 35453 5228
rect 35596 5188 39820 5228
rect 39860 5188 39869 5228
rect 40291 5188 40300 5228
rect 40340 5188 40876 5228
rect 40916 5188 40925 5228
rect 41635 5188 41644 5228
rect 41684 5188 44140 5228
rect 44180 5188 44189 5228
rect 46627 5188 46636 5228
rect 46676 5188 56620 5228
rect 56660 5188 56669 5228
rect 57006 5188 57100 5228
rect 57140 5188 57149 5228
rect 57196 5228 57236 5272
rect 57283 5272 57292 5312
rect 57332 5272 57426 5312
rect 57580 5272 57868 5312
rect 57908 5272 57917 5312
rect 58062 5272 58156 5312
rect 58196 5272 58205 5312
rect 59491 5272 59500 5312
rect 59540 5272 63860 5312
rect 64159 5272 64168 5312
rect 64208 5272 64250 5312
rect 64290 5272 64332 5312
rect 64372 5272 64414 5312
rect 64454 5272 64496 5312
rect 64536 5272 64545 5312
rect 65356 5272 67564 5312
rect 67604 5272 67613 5312
rect 69763 5272 69772 5312
rect 69812 5272 73900 5312
rect 73940 5272 73949 5312
rect 74467 5272 74476 5312
rect 74516 5272 74525 5312
rect 75043 5272 75052 5312
rect 75092 5272 75668 5312
rect 76099 5312 76157 5313
rect 77452 5312 77492 5440
rect 77827 5439 77885 5440
rect 78700 5396 78740 5440
rect 79747 5439 79805 5440
rect 80611 5439 80669 5440
rect 81859 5439 81917 5440
rect 81475 5396 81533 5397
rect 78700 5356 81484 5396
rect 81524 5356 81533 5396
rect 82348 5396 82388 5440
rect 82348 5356 93100 5396
rect 93140 5356 93149 5396
rect 81475 5355 81533 5356
rect 81667 5312 81725 5313
rect 76099 5272 76108 5312
rect 76148 5272 76876 5312
rect 76916 5272 76925 5312
rect 77452 5272 79084 5312
rect 79124 5272 79133 5312
rect 79279 5272 79288 5312
rect 79328 5272 79370 5312
rect 79410 5272 79452 5312
rect 79492 5272 79534 5312
rect 79574 5272 79616 5312
rect 79656 5272 79665 5312
rect 81091 5272 81100 5312
rect 81140 5272 81484 5312
rect 81524 5272 81533 5312
rect 81667 5272 81676 5312
rect 81716 5272 81810 5312
rect 83971 5272 83980 5312
rect 84020 5272 84364 5312
rect 84404 5272 84413 5312
rect 94399 5272 94408 5312
rect 94448 5272 94490 5312
rect 94530 5272 94572 5312
rect 94612 5272 94654 5312
rect 94694 5272 94736 5312
rect 94776 5272 94785 5312
rect 57283 5271 57341 5272
rect 58147 5271 58205 5272
rect 57196 5188 60940 5228
rect 60980 5188 60989 5228
rect 61795 5188 61804 5228
rect 61844 5188 62860 5228
rect 62900 5188 62909 5228
rect 20803 5187 20861 5188
rect 23971 5187 24029 5188
rect 24355 5187 24413 5188
rect 40291 5187 40349 5188
rect 41635 5187 41693 5188
rect 56611 5187 56669 5188
rect 57091 5187 57149 5188
rect 38083 5144 38141 5145
rect 63820 5144 63860 5272
rect 76099 5271 76157 5272
rect 81667 5271 81725 5272
rect 64003 5228 64061 5229
rect 67843 5228 67901 5229
rect 63918 5188 64012 5228
rect 64052 5188 64061 5228
rect 67747 5188 67756 5228
rect 67796 5188 67852 5228
rect 67892 5188 67901 5228
rect 64003 5187 64061 5188
rect 67843 5187 67901 5188
rect 68995 5228 69053 5229
rect 68995 5188 69004 5228
rect 69044 5188 71596 5228
rect 71636 5188 71645 5228
rect 72643 5188 72652 5228
rect 72692 5188 77548 5228
rect 77588 5188 77597 5228
rect 77731 5188 77740 5228
rect 77780 5188 79604 5228
rect 79843 5188 79852 5228
rect 79892 5188 82636 5228
rect 82676 5188 82685 5228
rect 83107 5188 83116 5228
rect 83156 5188 92332 5228
rect 92372 5188 92381 5228
rect 68995 5187 69053 5188
rect 68611 5144 68669 5145
rect 73699 5144 73757 5145
rect 76675 5144 76733 5145
rect 79564 5144 79604 5188
rect 3811 5104 3820 5144
rect 3860 5104 7468 5144
rect 7508 5104 7517 5144
rect 9283 5104 9292 5144
rect 9332 5104 15724 5144
rect 15764 5104 15773 5144
rect 16483 5104 16492 5144
rect 16532 5104 17836 5144
rect 17876 5104 17885 5144
rect 18211 5104 18220 5144
rect 18260 5104 18892 5144
rect 18932 5104 22828 5144
rect 22868 5104 22877 5144
rect 23011 5104 23020 5144
rect 23060 5104 25420 5144
rect 25460 5104 25469 5144
rect 27139 5104 27148 5144
rect 27188 5104 29548 5144
rect 29588 5104 29597 5144
rect 30691 5104 30700 5144
rect 30740 5104 34156 5144
rect 34196 5104 34205 5144
rect 34819 5104 34828 5144
rect 34868 5104 34877 5144
rect 35107 5104 35116 5144
rect 35156 5104 38092 5144
rect 38132 5104 38141 5144
rect 42691 5104 42700 5144
rect 42740 5104 44372 5144
rect 45571 5104 45580 5144
rect 45620 5104 52780 5144
rect 52820 5104 52829 5144
rect 53155 5104 53164 5144
rect 53204 5104 58732 5144
rect 58772 5104 58781 5144
rect 63820 5104 68044 5144
rect 68084 5104 68093 5144
rect 68611 5104 68620 5144
rect 68660 5104 69580 5144
rect 69620 5104 69629 5144
rect 70348 5104 73172 5144
rect 73507 5104 73516 5144
rect 73556 5104 73708 5144
rect 73748 5104 73757 5144
rect 73987 5104 73996 5144
rect 74036 5104 76108 5144
rect 76148 5104 76157 5144
rect 76675 5104 76684 5144
rect 76724 5104 76780 5144
rect 76820 5104 76829 5144
rect 77155 5104 77164 5144
rect 77204 5104 77452 5144
rect 77492 5104 77501 5144
rect 78019 5104 78028 5144
rect 78068 5104 78796 5144
rect 78836 5104 79372 5144
rect 79412 5104 79421 5144
rect 79555 5104 79564 5144
rect 79604 5104 79613 5144
rect 80803 5104 80812 5144
rect 80852 5104 81580 5144
rect 81620 5104 81629 5144
rect 81955 5104 81964 5144
rect 82004 5104 82732 5144
rect 82772 5104 82781 5144
rect 84259 5104 84268 5144
rect 84308 5104 89068 5144
rect 89108 5104 89117 5144
rect 19651 5060 19709 5061
rect 21379 5060 21437 5061
rect 21955 5060 22013 5061
rect 28579 5060 28637 5061
rect 34828 5060 34868 5104
rect 38083 5103 38141 5104
rect 44227 5060 44285 5061
rect 4195 5020 4204 5060
rect 4244 5020 6220 5060
rect 6260 5020 6269 5060
rect 11203 5020 11212 5060
rect 11252 5020 15340 5060
rect 15380 5020 15389 5060
rect 15526 5020 15535 5060
rect 15575 5020 16108 5060
rect 16148 5020 16157 5060
rect 16771 5020 16780 5060
rect 16820 5020 18604 5060
rect 18644 5020 18653 5060
rect 19651 5020 19660 5060
rect 19700 5020 19948 5060
rect 19988 5020 19997 5060
rect 20140 5020 21388 5060
rect 21428 5020 21437 5060
rect 21870 5020 21964 5060
rect 22004 5020 22013 5060
rect 22435 5020 22444 5060
rect 22484 5020 23596 5060
rect 23636 5020 25132 5060
rect 25172 5020 25181 5060
rect 25891 5020 25900 5060
rect 25940 5020 28396 5060
rect 28436 5020 28445 5060
rect 28579 5020 28588 5060
rect 28628 5020 29000 5060
rect 31651 5020 31660 5060
rect 31700 5020 31709 5060
rect 34828 5020 40972 5060
rect 41012 5020 41021 5060
rect 41539 5020 41548 5060
rect 41588 5020 42508 5060
rect 42548 5020 42557 5060
rect 42979 5020 42988 5060
rect 43028 5020 44236 5060
rect 44276 5020 44285 5060
rect 44332 5060 44372 5104
rect 68611 5103 68669 5104
rect 57475 5060 57533 5061
rect 44332 5020 49036 5060
rect 49076 5020 49085 5060
rect 49132 5020 52108 5060
rect 52148 5020 52157 5060
rect 57390 5020 57484 5060
rect 57524 5020 57533 5060
rect 19651 5019 19709 5020
rect 2083 4976 2141 4977
rect 2467 4976 2525 4977
rect 20140 4976 20180 5020
rect 21379 5019 21437 5020
rect 21955 5019 22013 5020
rect 28579 5019 28637 5020
rect 24835 4976 24893 4977
rect 28771 4976 28829 4977
rect 1998 4936 2092 4976
rect 2132 4936 2141 4976
rect 2382 4936 2476 4976
rect 2516 4936 2525 4976
rect 8803 4936 8812 4976
rect 8852 4936 11980 4976
rect 12020 4936 12029 4976
rect 13891 4936 13900 4976
rect 13940 4936 13949 4976
rect 14659 4936 14668 4976
rect 14708 4936 16916 4976
rect 19176 4936 19185 4976
rect 19225 4936 20180 4976
rect 20323 4936 20332 4976
rect 20372 4936 24652 4976
rect 24692 4936 24701 4976
rect 24835 4936 24844 4976
rect 24884 4936 28780 4976
rect 28820 4936 28829 4976
rect 28960 4976 29000 5020
rect 31660 4976 31700 5020
rect 44227 5019 44285 5020
rect 34531 4976 34589 4977
rect 38179 4976 38237 4977
rect 47299 4976 47357 4977
rect 48355 4976 48413 4977
rect 49132 4976 49172 5020
rect 57475 5019 57533 5020
rect 57859 5060 57917 5061
rect 68707 5060 68765 5061
rect 70348 5060 70388 5104
rect 71875 5060 71933 5061
rect 73132 5060 73172 5104
rect 73699 5103 73757 5104
rect 76675 5103 76733 5104
rect 57859 5020 57868 5060
rect 57908 5020 59348 5060
rect 60163 5020 60172 5060
rect 60212 5020 62764 5060
rect 62804 5020 62813 5060
rect 62947 5020 62956 5060
rect 62996 5020 64780 5060
rect 64820 5020 64829 5060
rect 67651 5020 67660 5060
rect 67700 5020 68428 5060
rect 68468 5020 68477 5060
rect 68707 5020 68716 5060
rect 68756 5020 70348 5060
rect 70388 5020 70397 5060
rect 71683 5020 71692 5060
rect 71732 5020 71884 5060
rect 71924 5020 71933 5060
rect 72163 5020 72172 5060
rect 72212 5020 72556 5060
rect 72596 5020 72844 5060
rect 72884 5020 72893 5060
rect 73132 5020 75820 5060
rect 75860 5020 75869 5060
rect 75919 5020 75928 5060
rect 75968 5020 78508 5060
rect 78548 5020 78557 5060
rect 79459 5020 79468 5060
rect 79508 5020 79852 5060
rect 79892 5020 79901 5060
rect 80035 5020 80044 5060
rect 80084 5020 83020 5060
rect 83060 5020 83069 5060
rect 84067 5020 84076 5060
rect 84116 5020 85324 5060
rect 85364 5020 85373 5060
rect 86947 5020 86956 5060
rect 86996 5020 88780 5060
rect 88820 5020 88829 5060
rect 89731 5020 89740 5060
rect 89780 5020 91276 5060
rect 91316 5020 91325 5060
rect 57859 5019 57917 5020
rect 56611 4976 56669 4977
rect 58243 4976 58301 4977
rect 28960 4936 30700 4976
rect 30740 4936 30749 4976
rect 31660 4936 33004 4976
rect 33044 4936 33053 4976
rect 33379 4936 33388 4976
rect 33428 4936 33437 4976
rect 33571 4936 33580 4976
rect 33620 4936 33772 4976
rect 33812 4936 33821 4976
rect 34531 4936 34540 4976
rect 34580 4936 36460 4976
rect 36500 4936 36509 4976
rect 36643 4936 36652 4976
rect 36692 4936 37516 4976
rect 37556 4936 37565 4976
rect 38179 4936 38188 4976
rect 38228 4936 41600 4976
rect 46147 4936 46156 4976
rect 46196 4936 46636 4976
rect 46676 4936 46685 4976
rect 46819 4936 46828 4976
rect 46868 4936 47308 4976
rect 47348 4936 47788 4976
rect 47828 4936 47837 4976
rect 48270 4936 48364 4976
rect 48404 4936 48413 4976
rect 48739 4936 48748 4976
rect 48788 4936 48797 4976
rect 48931 4936 48940 4976
rect 48980 4936 49172 4976
rect 50467 4936 50476 4976
rect 50516 4936 50956 4976
rect 50996 4936 51005 4976
rect 52387 4936 52396 4976
rect 52436 4936 52876 4976
rect 52916 4936 52925 4976
rect 55420 4936 56468 4976
rect 2083 4935 2141 4936
rect 2467 4935 2525 4936
rect 1603 4852 1612 4892
rect 1652 4852 10252 4892
rect 10292 4852 10301 4892
rect 13900 4808 13940 4936
rect 15427 4852 15436 4892
rect 15476 4852 16532 4892
rect 1699 4768 1708 4808
rect 1748 4768 10348 4808
rect 10388 4768 10397 4808
rect 13900 4768 15052 4808
rect 15092 4768 15101 4808
rect 15619 4724 15677 4725
rect 9187 4684 9196 4724
rect 9236 4684 12652 4724
rect 12692 4684 12701 4724
rect 15534 4684 15628 4724
rect 15668 4684 15677 4724
rect 16492 4724 16532 4852
rect 16876 4808 16916 4936
rect 24835 4935 24893 4936
rect 28771 4935 28829 4936
rect 17539 4892 17597 4893
rect 19939 4892 19997 4893
rect 21283 4892 21341 4893
rect 27619 4892 27677 4893
rect 17347 4852 17356 4892
rect 17396 4852 17548 4892
rect 17588 4852 17597 4892
rect 18787 4852 18796 4892
rect 18836 4852 19948 4892
rect 19988 4852 20121 4892
rect 20161 4852 20170 4892
rect 20899 4852 20908 4892
rect 20948 4852 21292 4892
rect 21332 4852 21341 4892
rect 17539 4851 17597 4852
rect 19939 4851 19997 4852
rect 21283 4851 21341 4852
rect 21484 4852 21868 4892
rect 21908 4852 22252 4892
rect 22292 4852 22301 4892
rect 23212 4852 23636 4892
rect 24163 4852 24172 4892
rect 24212 4852 24556 4892
rect 24596 4852 24940 4892
rect 24980 4852 25324 4892
rect 25364 4852 25373 4892
rect 26659 4852 26668 4892
rect 26708 4852 26956 4892
rect 26996 4852 27005 4892
rect 27534 4852 27628 4892
rect 27668 4852 27677 4892
rect 27811 4852 27820 4892
rect 27860 4852 28012 4892
rect 28052 4852 28436 4892
rect 28867 4852 28876 4892
rect 28916 4852 29000 4892
rect 30499 4852 30508 4892
rect 30548 4852 30892 4892
rect 30932 4852 30941 4892
rect 31555 4852 31564 4892
rect 31604 4852 31613 4892
rect 21484 4808 21524 4852
rect 23212 4808 23252 4852
rect 16876 4768 19084 4808
rect 19124 4768 19133 4808
rect 19948 4768 21428 4808
rect 21475 4768 21484 4808
rect 21524 4768 21533 4808
rect 21580 4768 22540 4808
rect 22580 4768 23252 4808
rect 23299 4808 23357 4809
rect 23299 4768 23308 4808
rect 23348 4768 23404 4808
rect 23444 4768 23453 4808
rect 18499 4724 18557 4725
rect 19363 4724 19421 4725
rect 19948 4724 19988 4768
rect 21187 4724 21245 4725
rect 16492 4684 18316 4724
rect 18356 4684 18365 4724
rect 18414 4684 18508 4724
rect 18548 4684 18557 4724
rect 19278 4684 19372 4724
rect 19412 4684 19421 4724
rect 19939 4684 19948 4724
rect 19988 4684 19997 4724
rect 20707 4684 20716 4724
rect 20756 4684 21196 4724
rect 21236 4684 21245 4724
rect 21388 4724 21428 4768
rect 21580 4724 21620 4768
rect 23299 4767 23357 4768
rect 22339 4724 22397 4725
rect 23596 4724 23636 4852
rect 27619 4851 27677 4852
rect 25507 4808 25565 4809
rect 28396 4808 28436 4852
rect 28960 4808 29000 4852
rect 31459 4808 31517 4809
rect 23779 4768 23788 4808
rect 23828 4768 25228 4808
rect 25268 4768 25277 4808
rect 25422 4768 25516 4808
rect 25556 4768 25565 4808
rect 26467 4768 26476 4808
rect 26516 4768 28244 4808
rect 28387 4768 28396 4808
rect 28436 4768 28780 4808
rect 28820 4768 28829 4808
rect 28960 4768 31468 4808
rect 31508 4768 31517 4808
rect 31564 4808 31604 4852
rect 31564 4768 32716 4808
rect 32756 4768 32765 4808
rect 25507 4767 25565 4768
rect 24835 4724 24893 4725
rect 25027 4724 25085 4725
rect 28204 4724 28244 4768
rect 31459 4767 31517 4768
rect 30595 4724 30653 4725
rect 21388 4684 21620 4724
rect 22254 4684 22348 4724
rect 22388 4684 22397 4724
rect 22819 4684 22828 4724
rect 22868 4684 23212 4724
rect 23252 4684 23261 4724
rect 23596 4684 24844 4724
rect 24884 4684 24893 4724
rect 24942 4684 25036 4724
rect 25076 4684 25085 4724
rect 25315 4684 25324 4724
rect 25364 4684 28108 4724
rect 28148 4684 28157 4724
rect 28204 4684 28972 4724
rect 29012 4684 29021 4724
rect 29347 4684 29356 4724
rect 29396 4684 29836 4724
rect 29876 4684 29885 4724
rect 30124 4684 30316 4724
rect 30356 4684 30604 4724
rect 30644 4684 30653 4724
rect 30787 4684 30796 4724
rect 30836 4684 31564 4724
rect 31604 4684 31613 4724
rect 15619 4683 15677 4684
rect 18499 4683 18557 4684
rect 19363 4683 19421 4684
rect 21187 4683 21245 4684
rect 22339 4683 22397 4684
rect 24835 4683 24893 4684
rect 25027 4683 25085 4684
rect 17155 4640 17213 4641
rect 9379 4600 9388 4640
rect 9428 4600 12364 4640
rect 12404 4600 12413 4640
rect 17070 4600 17164 4640
rect 17204 4600 17213 4640
rect 17155 4599 17213 4600
rect 17347 4640 17405 4641
rect 23203 4640 23261 4641
rect 30124 4640 30164 4684
rect 30595 4683 30653 4684
rect 33388 4640 33428 4936
rect 34531 4935 34589 4936
rect 38179 4935 38237 4936
rect 35491 4892 35549 4893
rect 37027 4892 37085 4893
rect 34243 4852 34252 4892
rect 34292 4852 34540 4892
rect 34580 4852 34589 4892
rect 34723 4852 34732 4892
rect 34772 4852 35116 4892
rect 35156 4852 35500 4892
rect 35540 4852 35884 4892
rect 35924 4852 36268 4892
rect 36308 4852 36556 4892
rect 36596 4852 36605 4892
rect 36942 4852 37036 4892
rect 37076 4852 37085 4892
rect 35491 4851 35549 4852
rect 37027 4851 37085 4852
rect 37219 4892 37277 4893
rect 41560 4892 41600 4936
rect 47299 4935 47357 4936
rect 48355 4935 48413 4936
rect 48748 4892 48788 4936
rect 37219 4852 37228 4892
rect 37268 4852 37362 4892
rect 39331 4852 39340 4892
rect 39380 4852 39628 4892
rect 39668 4852 39677 4892
rect 41560 4852 48788 4892
rect 37219 4851 37277 4852
rect 38851 4808 38909 4809
rect 34540 4768 35308 4808
rect 35348 4768 37612 4808
rect 37652 4768 37661 4808
rect 37804 4768 38668 4808
rect 38708 4768 38860 4808
rect 38900 4768 38909 4808
rect 33571 4684 33580 4724
rect 33620 4684 33772 4724
rect 33812 4684 33821 4724
rect 17347 4600 17356 4640
rect 17396 4600 17490 4640
rect 17731 4600 17740 4640
rect 17780 4600 18988 4640
rect 19028 4600 19852 4640
rect 19892 4600 21100 4640
rect 21140 4600 22252 4640
rect 22292 4600 23212 4640
rect 23252 4600 23261 4640
rect 24355 4600 24364 4640
rect 24404 4600 27820 4640
rect 27860 4600 30164 4640
rect 30211 4600 30220 4640
rect 30260 4600 33428 4640
rect 33475 4640 33533 4641
rect 33475 4600 33484 4640
rect 33524 4600 34060 4640
rect 34100 4600 34109 4640
rect 17347 4599 17405 4600
rect 23203 4599 23261 4600
rect 20707 4556 20765 4557
rect 24364 4556 24404 4600
rect 33475 4599 33533 4600
rect 28771 4556 28829 4557
rect 34243 4556 34301 4557
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 14659 4516 14668 4556
rect 14708 4516 18124 4556
rect 18164 4516 18173 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20622 4516 20716 4556
rect 20756 4516 20765 4556
rect 21283 4516 21292 4556
rect 21332 4516 22156 4556
rect 22196 4516 24404 4556
rect 24739 4516 24748 4556
rect 24788 4516 28204 4556
rect 28244 4516 28588 4556
rect 28628 4516 28637 4556
rect 28771 4516 28780 4556
rect 28820 4516 29164 4556
rect 29204 4516 33868 4556
rect 33908 4516 33917 4556
rect 34243 4516 34252 4556
rect 34292 4516 34348 4556
rect 34388 4516 34397 4556
rect 20707 4515 20765 4516
rect 17347 4472 17405 4473
rect 19363 4472 19421 4473
rect 21187 4472 21245 4473
rect 24748 4472 24788 4516
rect 28771 4515 28829 4516
rect 34243 4515 34301 4516
rect 34540 4472 34580 4768
rect 35491 4724 35549 4725
rect 35971 4724 36029 4725
rect 37804 4724 37844 4768
rect 38851 4767 38909 4768
rect 39043 4808 39101 4809
rect 48940 4808 48980 4936
rect 49507 4892 49565 4893
rect 49422 4852 49516 4892
rect 49556 4852 49565 4892
rect 49699 4852 49708 4892
rect 49748 4852 49900 4892
rect 49940 4852 51724 4892
rect 51764 4852 51773 4892
rect 54787 4852 54796 4892
rect 54836 4852 55180 4892
rect 55220 4852 55229 4892
rect 49507 4851 49565 4852
rect 55420 4808 55460 4936
rect 56428 4892 56468 4936
rect 56611 4936 56620 4976
rect 56660 4936 56715 4976
rect 56755 4936 56764 4976
rect 56899 4936 56908 4976
rect 56948 4936 57964 4976
rect 58004 4936 58013 4976
rect 58243 4936 58252 4976
rect 58292 4936 59212 4976
rect 59252 4936 59261 4976
rect 56611 4935 56669 4936
rect 58243 4935 58301 4936
rect 57475 4892 57533 4893
rect 55939 4852 55948 4892
rect 55988 4852 56332 4892
rect 56372 4852 56381 4892
rect 56428 4852 57484 4892
rect 57524 4852 57533 4892
rect 57667 4852 57676 4892
rect 57716 4852 58252 4892
rect 58292 4852 58301 4892
rect 58435 4852 58444 4892
rect 58484 4852 58493 4892
rect 59011 4852 59020 4892
rect 59060 4852 59069 4892
rect 39043 4768 39052 4808
rect 39092 4768 42220 4808
rect 42260 4768 42269 4808
rect 46531 4768 46540 4808
rect 46580 4768 47020 4808
rect 47060 4768 47500 4808
rect 47540 4768 47549 4808
rect 47596 4768 48980 4808
rect 49987 4768 49996 4808
rect 50036 4768 50572 4808
rect 50612 4768 50621 4808
rect 53923 4768 53932 4808
rect 53972 4768 55460 4808
rect 39043 4767 39101 4768
rect 47596 4724 47636 4768
rect 55948 4724 55988 4852
rect 57475 4851 57533 4852
rect 58444 4808 58484 4852
rect 56611 4768 56620 4808
rect 56660 4768 57868 4808
rect 57908 4768 57917 4808
rect 58060 4768 58484 4808
rect 35011 4684 35020 4724
rect 35060 4684 35069 4724
rect 35406 4684 35500 4724
rect 35540 4684 35549 4724
rect 35683 4684 35692 4724
rect 35732 4684 35980 4724
rect 36020 4684 36029 4724
rect 36163 4684 36172 4724
rect 36212 4684 37844 4724
rect 38371 4684 38380 4724
rect 38420 4684 41836 4724
rect 41876 4684 41885 4724
rect 45571 4684 45580 4724
rect 45620 4684 45868 4724
rect 45908 4684 45917 4724
rect 47107 4684 47116 4724
rect 47156 4684 47636 4724
rect 47779 4684 47788 4724
rect 47828 4684 48460 4724
rect 48500 4684 48509 4724
rect 49219 4684 49228 4724
rect 49268 4684 49612 4724
rect 49652 4684 49804 4724
rect 49844 4684 50188 4724
rect 50228 4684 50237 4724
rect 50371 4684 50380 4724
rect 50420 4684 50860 4724
rect 50900 4684 50909 4724
rect 53251 4684 53260 4724
rect 53300 4684 55988 4724
rect 56227 4724 56285 4725
rect 56803 4724 56861 4725
rect 58060 4724 58100 4768
rect 59020 4724 59060 4852
rect 59308 4808 59348 5020
rect 68707 5019 68765 5020
rect 71875 5019 71933 5020
rect 67939 4976 67997 4977
rect 73132 4976 73172 5020
rect 76003 4976 76061 4977
rect 76771 4976 76829 4977
rect 87043 4976 87101 4977
rect 87715 4976 87773 4977
rect 88483 4976 88541 4977
rect 97699 4976 97757 4977
rect 98083 4976 98141 4977
rect 59395 4936 59404 4976
rect 59444 4936 59692 4976
rect 59732 4936 64396 4976
rect 64436 4936 64445 4976
rect 64579 4936 64588 4976
rect 64628 4936 67180 4976
rect 67220 4936 67229 4976
rect 67854 4936 67948 4976
rect 67988 4936 67997 4976
rect 68131 4936 68140 4976
rect 68180 4936 68220 4976
rect 69667 4936 69676 4976
rect 69716 4936 70924 4976
rect 70964 4936 70973 4976
rect 71116 4936 72364 4976
rect 72404 4936 72413 4976
rect 73123 4936 73132 4976
rect 73172 4936 73181 4976
rect 74179 4936 74188 4976
rect 74228 4936 76012 4976
rect 76052 4936 76061 4976
rect 76291 4936 76300 4976
rect 76340 4936 76588 4976
rect 76628 4936 76637 4976
rect 76771 4936 76780 4976
rect 76820 4936 79276 4976
rect 79316 4936 79325 4976
rect 80899 4936 80908 4976
rect 80948 4936 86132 4976
rect 86958 4936 87052 4976
rect 87092 4936 87101 4976
rect 87630 4936 87724 4976
rect 87764 4936 87773 4976
rect 88099 4936 88108 4976
rect 88148 4936 88340 4976
rect 88398 4936 88492 4976
rect 88532 4936 88541 4976
rect 91939 4936 91948 4976
rect 91988 4936 97132 4976
rect 97172 4936 97181 4976
rect 97614 4936 97708 4976
rect 97748 4936 97757 4976
rect 97998 4936 98092 4976
rect 98132 4936 98141 4976
rect 98467 4936 98476 4976
rect 98516 4936 98525 4976
rect 63235 4892 63293 4893
rect 60067 4852 60076 4892
rect 60116 4852 61748 4892
rect 63150 4852 63244 4892
rect 63284 4852 63293 4892
rect 63427 4852 63436 4892
rect 63476 4852 66932 4892
rect 61708 4808 61748 4852
rect 63235 4851 63293 4852
rect 66892 4808 66932 4852
rect 67180 4808 67220 4936
rect 67939 4935 67997 4936
rect 68140 4892 68180 4936
rect 71116 4892 71156 4936
rect 76003 4935 76061 4936
rect 72643 4892 72701 4893
rect 73411 4892 73469 4893
rect 76588 4892 76628 4936
rect 76771 4935 76829 4936
rect 77251 4892 77309 4893
rect 67363 4852 67372 4892
rect 67412 4852 67756 4892
rect 67796 4852 68524 4892
rect 68564 4852 68573 4892
rect 69763 4852 69772 4892
rect 69812 4852 70156 4892
rect 70196 4852 70540 4892
rect 70580 4852 70828 4892
rect 70868 4852 70877 4892
rect 71107 4852 71116 4892
rect 71156 4852 71165 4892
rect 71299 4852 71308 4892
rect 71348 4852 71692 4892
rect 71732 4852 72212 4892
rect 68227 4808 68285 4809
rect 72067 4808 72125 4809
rect 59308 4768 61652 4808
rect 61708 4768 64280 4808
rect 66883 4768 66892 4808
rect 66932 4768 66941 4808
rect 67180 4768 68180 4808
rect 61612 4724 61652 4768
rect 56227 4684 56236 4724
rect 56276 4684 56524 4724
rect 56564 4684 56573 4724
rect 56803 4684 56812 4724
rect 56852 4684 57100 4724
rect 57140 4684 57149 4724
rect 57283 4684 57292 4724
rect 57332 4684 58060 4724
rect 58100 4684 58109 4724
rect 58435 4684 58444 4724
rect 58484 4684 59060 4724
rect 59107 4684 59116 4724
rect 59156 4684 60172 4724
rect 60212 4684 60221 4724
rect 61603 4684 61612 4724
rect 61652 4684 61661 4724
rect 62851 4684 62860 4724
rect 62900 4684 64108 4724
rect 64148 4684 64157 4724
rect 35020 4640 35060 4684
rect 35491 4683 35549 4684
rect 35971 4683 36029 4684
rect 56227 4683 56285 4684
rect 56803 4683 56861 4684
rect 56236 4640 56276 4683
rect 35020 4600 40108 4640
rect 40148 4600 40157 4640
rect 44323 4600 44332 4640
rect 44372 4600 44524 4640
rect 44564 4600 54028 4640
rect 54068 4600 54077 4640
rect 54499 4600 54508 4640
rect 54548 4600 56276 4640
rect 56515 4640 56573 4641
rect 64240 4640 64280 4768
rect 68140 4724 68180 4768
rect 68227 4768 68236 4808
rect 68276 4768 68332 4808
rect 68372 4768 68381 4808
rect 68803 4768 68812 4808
rect 68852 4768 69524 4808
rect 70435 4768 70444 4808
rect 70484 4768 70964 4808
rect 71982 4768 72076 4808
rect 72116 4768 72125 4808
rect 72172 4808 72212 4852
rect 72643 4852 72652 4892
rect 72692 4852 72940 4892
rect 72980 4852 73420 4892
rect 73460 4852 73469 4892
rect 73603 4852 73612 4892
rect 73652 4852 75148 4892
rect 75188 4852 75197 4892
rect 75244 4852 76396 4892
rect 76436 4852 76445 4892
rect 76588 4852 76972 4892
rect 77012 4852 77021 4892
rect 77166 4852 77260 4892
rect 77300 4852 77309 4892
rect 72643 4851 72701 4852
rect 73411 4851 73469 4852
rect 75244 4808 75284 4852
rect 77251 4851 77309 4852
rect 77539 4892 77597 4893
rect 85795 4892 85853 4893
rect 86092 4892 86132 4936
rect 87043 4935 87101 4936
rect 87715 4935 87773 4936
rect 77539 4852 77548 4892
rect 77588 4852 77836 4892
rect 77876 4852 77885 4892
rect 81763 4852 81772 4892
rect 81812 4852 82924 4892
rect 82964 4852 83500 4892
rect 83540 4852 84268 4892
rect 84308 4852 84317 4892
rect 84643 4852 84652 4892
rect 84692 4852 85612 4892
rect 85652 4852 85661 4892
rect 85795 4852 85804 4892
rect 85844 4852 85996 4892
rect 86036 4852 86045 4892
rect 86092 4852 88204 4892
rect 88244 4852 88253 4892
rect 77539 4851 77597 4852
rect 85795 4851 85853 4852
rect 85603 4808 85661 4809
rect 88300 4808 88340 4936
rect 88483 4935 88541 4936
rect 97699 4935 97757 4936
rect 98083 4935 98141 4936
rect 98476 4892 98516 4936
rect 88675 4852 88684 4892
rect 88724 4852 98516 4892
rect 72172 4768 73324 4808
rect 73364 4768 74860 4808
rect 74900 4768 75284 4808
rect 76195 4768 76204 4808
rect 76244 4768 76253 4808
rect 76300 4768 85036 4808
rect 85076 4768 85085 4808
rect 85603 4768 85612 4808
rect 85652 4768 88340 4808
rect 89635 4768 89644 4808
rect 89684 4768 93292 4808
rect 93332 4768 93341 4808
rect 68227 4767 68285 4768
rect 64387 4684 64396 4724
rect 64436 4684 67892 4724
rect 68140 4684 69292 4724
rect 69332 4684 69341 4724
rect 67555 4640 67613 4641
rect 56515 4600 56524 4640
rect 56564 4600 62764 4640
rect 62804 4600 62813 4640
rect 64240 4600 67564 4640
rect 67604 4600 67613 4640
rect 67852 4640 67892 4684
rect 68611 4640 68669 4641
rect 67852 4600 68620 4640
rect 68660 4600 68669 4640
rect 56515 4599 56573 4600
rect 67555 4599 67613 4600
rect 68611 4599 68669 4600
rect 61699 4556 61757 4557
rect 68707 4556 68765 4557
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 35587 4516 35596 4556
rect 35636 4516 36692 4556
rect 36739 4516 36748 4556
rect 36788 4516 37996 4556
rect 38036 4516 38045 4556
rect 38947 4516 38956 4556
rect 38996 4516 47980 4556
rect 48020 4516 48029 4556
rect 50179 4516 50188 4556
rect 50228 4516 50237 4556
rect 50279 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50665 4556
rect 53251 4516 53260 4556
rect 53300 4516 54316 4556
rect 54356 4516 54365 4556
rect 55747 4516 55756 4556
rect 55796 4516 58444 4556
rect 58484 4516 58493 4556
rect 61219 4516 61228 4556
rect 61268 4516 61708 4556
rect 61748 4516 61900 4556
rect 61940 4516 61949 4556
rect 62467 4516 62476 4556
rect 62516 4516 63052 4556
rect 63092 4516 63101 4556
rect 65399 4516 65408 4556
rect 65448 4516 65490 4556
rect 65530 4516 65572 4556
rect 65612 4516 65654 4556
rect 65694 4516 65736 4556
rect 65776 4516 65785 4556
rect 66796 4516 68524 4556
rect 68564 4516 68716 4556
rect 68756 4516 68765 4556
rect 69484 4556 69524 4768
rect 70723 4724 70781 4725
rect 70924 4724 70964 4768
rect 72067 4767 72125 4768
rect 71203 4724 71261 4725
rect 72643 4724 72701 4725
rect 72835 4724 72893 4725
rect 76204 4724 76244 4768
rect 76300 4724 76340 4768
rect 85603 4767 85661 4768
rect 76771 4724 76829 4725
rect 81283 4724 81341 4725
rect 88963 4724 89021 4725
rect 70638 4684 70732 4724
rect 70772 4684 70781 4724
rect 70915 4684 70924 4724
rect 70964 4684 70973 4724
rect 71118 4684 71212 4724
rect 71252 4684 71261 4724
rect 72163 4684 72172 4724
rect 72212 4684 72652 4724
rect 72692 4684 72701 4724
rect 72750 4684 72844 4724
rect 72884 4684 72893 4724
rect 73891 4684 73900 4724
rect 73940 4684 75724 4724
rect 75764 4684 76244 4724
rect 76291 4684 76300 4724
rect 76340 4684 76349 4724
rect 76686 4684 76780 4724
rect 76820 4684 76829 4724
rect 81198 4684 81292 4724
rect 81332 4684 81341 4724
rect 82147 4684 82156 4724
rect 82196 4684 82444 4724
rect 82484 4684 82493 4724
rect 83395 4684 83404 4724
rect 83444 4684 83884 4724
rect 83924 4684 83933 4724
rect 84259 4684 84268 4724
rect 84308 4684 84940 4724
rect 84980 4684 84989 4724
rect 85795 4684 85804 4724
rect 85844 4684 86764 4724
rect 86804 4684 86813 4724
rect 88878 4684 88972 4724
rect 89012 4684 89021 4724
rect 98275 4684 98284 4724
rect 98324 4684 98476 4724
rect 98516 4684 98525 4724
rect 70723 4683 70781 4684
rect 71203 4683 71261 4684
rect 72643 4683 72701 4684
rect 72835 4683 72893 4684
rect 76771 4683 76829 4684
rect 81283 4683 81341 4684
rect 88963 4683 89021 4684
rect 69955 4640 70013 4641
rect 74083 4640 74141 4641
rect 75139 4640 75197 4641
rect 69870 4600 69964 4640
rect 70004 4600 70013 4640
rect 69955 4599 70013 4600
rect 70060 4600 71596 4640
rect 71636 4600 72748 4640
rect 72788 4600 72797 4640
rect 73998 4600 74092 4640
rect 74132 4600 74141 4640
rect 75054 4600 75148 4640
rect 75188 4600 75197 4640
rect 75523 4600 75532 4640
rect 75572 4600 86572 4640
rect 86612 4600 86621 4640
rect 70060 4556 70100 4600
rect 74083 4599 74141 4600
rect 75139 4599 75197 4600
rect 71875 4556 71933 4557
rect 80419 4556 80477 4557
rect 69484 4516 69868 4556
rect 69908 4516 69917 4556
rect 70051 4516 70060 4556
rect 70100 4516 70109 4556
rect 71875 4516 71884 4556
rect 71924 4516 72076 4556
rect 72116 4516 72125 4556
rect 72547 4516 72556 4556
rect 72596 4516 72940 4556
rect 72980 4516 73708 4556
rect 73748 4516 76012 4556
rect 76052 4516 76684 4556
rect 76724 4516 76733 4556
rect 80334 4516 80428 4556
rect 80468 4516 80477 4556
rect 80519 4516 80528 4556
rect 80568 4516 80610 4556
rect 80650 4516 80692 4556
rect 80732 4516 80774 4556
rect 80814 4516 80856 4556
rect 80896 4516 80905 4556
rect 81004 4516 82732 4556
rect 82772 4516 82781 4556
rect 83779 4516 83788 4556
rect 83828 4516 84076 4556
rect 84116 4516 84125 4556
rect 84259 4516 84268 4556
rect 84308 4516 84556 4556
rect 84596 4516 84605 4556
rect 85411 4516 85420 4556
rect 85460 4516 86668 4556
rect 86708 4516 86717 4556
rect 86851 4516 86860 4556
rect 86900 4516 93580 4556
rect 93620 4516 93629 4556
rect 95639 4516 95648 4556
rect 95688 4516 95730 4556
rect 95770 4516 95812 4556
rect 95852 4516 95894 4556
rect 95934 4516 95976 4556
rect 96016 4516 96025 4556
rect 36547 4472 36605 4473
rect 13027 4432 13036 4472
rect 13076 4432 17356 4472
rect 17396 4432 17405 4472
rect 17539 4432 17548 4472
rect 17588 4432 19180 4472
rect 19220 4432 19229 4472
rect 19363 4432 19372 4472
rect 19412 4432 20812 4472
rect 20852 4432 20861 4472
rect 21187 4432 21196 4472
rect 21236 4432 21484 4472
rect 21524 4432 21533 4472
rect 21667 4432 21676 4472
rect 21716 4432 22828 4472
rect 22868 4432 24788 4472
rect 26764 4432 27244 4472
rect 27284 4432 27293 4472
rect 27907 4432 27916 4472
rect 27956 4432 30796 4472
rect 30836 4432 30845 4472
rect 31075 4432 31084 4472
rect 31124 4432 34580 4472
rect 34627 4432 34636 4472
rect 34676 4432 36556 4472
rect 36596 4432 36605 4472
rect 36652 4472 36692 4516
rect 39043 4472 39101 4473
rect 50188 4472 50228 4516
rect 61699 4515 61757 4516
rect 55555 4472 55613 4473
rect 56707 4472 56765 4473
rect 66796 4472 66836 4516
rect 68707 4515 68765 4516
rect 71875 4515 71933 4516
rect 80419 4515 80477 4516
rect 73027 4472 73085 4473
rect 77251 4472 77309 4473
rect 81004 4472 81044 4516
rect 36652 4432 39052 4472
rect 39092 4432 39101 4472
rect 39811 4432 39820 4472
rect 39860 4432 41600 4472
rect 46627 4432 46636 4472
rect 46676 4432 55564 4472
rect 55604 4432 56236 4472
rect 56276 4432 56285 4472
rect 56622 4432 56716 4472
rect 56756 4432 56765 4472
rect 56995 4432 57004 4472
rect 57044 4432 57388 4472
rect 57428 4432 57437 4472
rect 57571 4432 57580 4472
rect 57620 4432 62380 4472
rect 62420 4432 62429 4472
rect 63523 4432 63532 4472
rect 63572 4432 63724 4472
rect 63764 4432 63773 4472
rect 64195 4432 64204 4472
rect 64244 4432 66836 4472
rect 66883 4432 66892 4472
rect 66932 4432 67756 4472
rect 67796 4432 69580 4472
rect 69620 4432 71596 4472
rect 71636 4432 71980 4472
rect 72020 4432 72029 4472
rect 73027 4432 73036 4472
rect 73076 4432 73228 4472
rect 73268 4432 73277 4472
rect 77251 4432 77260 4472
rect 77300 4432 78988 4472
rect 79028 4432 79037 4472
rect 79267 4432 79276 4472
rect 79316 4432 81044 4472
rect 81475 4432 81484 4472
rect 81524 4432 87436 4472
rect 87476 4432 87485 4472
rect 17347 4431 17405 4432
rect 19363 4431 19421 4432
rect 21187 4431 21245 4432
rect 24643 4388 24701 4389
rect 26764 4388 26804 4432
rect 36547 4431 36605 4432
rect 39043 4431 39101 4432
rect 35011 4388 35069 4389
rect 35779 4388 35837 4389
rect 5059 4348 5068 4388
rect 5108 4348 5452 4388
rect 5492 4348 5501 4388
rect 13795 4348 13804 4388
rect 13844 4348 21196 4388
rect 21236 4348 21245 4388
rect 21292 4348 24268 4388
rect 24308 4348 24317 4388
rect 24558 4348 24652 4388
rect 24692 4348 26804 4388
rect 26851 4348 26860 4388
rect 26900 4348 28876 4388
rect 28916 4348 28925 4388
rect 30691 4348 30700 4388
rect 30740 4348 34252 4388
rect 34292 4348 34301 4388
rect 34926 4348 35020 4388
rect 35060 4348 35069 4388
rect 35694 4348 35788 4388
rect 35828 4348 35837 4388
rect 21292 4304 21332 4348
rect 24643 4347 24701 4348
rect 35011 4347 35069 4348
rect 35779 4347 35837 4348
rect 37795 4388 37853 4389
rect 41560 4388 41600 4432
rect 55555 4431 55613 4432
rect 56707 4431 56765 4432
rect 50371 4388 50429 4389
rect 55267 4388 55325 4389
rect 37795 4348 37804 4388
rect 37844 4348 37938 4388
rect 38755 4348 38764 4388
rect 38804 4348 41356 4388
rect 41396 4348 41405 4388
rect 41560 4348 45484 4388
rect 45524 4348 45533 4388
rect 45955 4348 45964 4388
rect 46004 4348 50380 4388
rect 50420 4348 50429 4388
rect 52195 4348 52204 4388
rect 52244 4348 54508 4388
rect 54548 4348 54557 4388
rect 55182 4348 55276 4388
rect 55316 4348 55325 4388
rect 37795 4347 37853 4348
rect 50371 4347 50429 4348
rect 55267 4347 55325 4348
rect 55843 4388 55901 4389
rect 61795 4388 61853 4389
rect 70435 4388 70493 4389
rect 55843 4348 55852 4388
rect 55892 4348 58772 4388
rect 58819 4348 58828 4388
rect 58868 4348 61228 4388
rect 61268 4348 61277 4388
rect 61795 4348 61804 4388
rect 61844 4348 63436 4388
rect 63476 4348 63485 4388
rect 64291 4348 64300 4388
rect 64340 4348 65972 4388
rect 66019 4348 66028 4388
rect 66068 4348 69004 4388
rect 69044 4348 69053 4388
rect 69100 4348 70444 4388
rect 70484 4348 71020 4388
rect 71060 4348 71069 4388
rect 55843 4347 55901 4348
rect 22723 4304 22781 4305
rect 23395 4304 23453 4305
rect 31459 4304 31517 4305
rect 7651 4264 7660 4304
rect 7700 4264 10732 4304
rect 10772 4264 10781 4304
rect 15715 4264 15724 4304
rect 15764 4264 19468 4304
rect 19508 4264 19517 4304
rect 20323 4264 20332 4304
rect 20372 4264 21332 4304
rect 22638 4264 22732 4304
rect 22772 4264 22781 4304
rect 23310 4264 23404 4304
rect 23444 4264 23453 4304
rect 25507 4264 25516 4304
rect 25556 4264 28204 4304
rect 28244 4264 31084 4304
rect 31124 4264 31133 4304
rect 31374 4264 31468 4304
rect 31508 4264 31517 4304
rect 22723 4263 22781 4264
rect 23395 4263 23453 4264
rect 31459 4263 31517 4264
rect 31651 4304 31709 4305
rect 58732 4304 58772 4348
rect 61795 4347 61853 4348
rect 65443 4304 65501 4305
rect 31651 4264 31660 4304
rect 31700 4264 32236 4304
rect 32276 4264 32285 4304
rect 32707 4264 32716 4304
rect 32756 4264 36076 4304
rect 36116 4264 36125 4304
rect 37603 4264 37612 4304
rect 37652 4264 47596 4304
rect 47636 4264 47645 4304
rect 49027 4264 49036 4304
rect 49076 4264 52972 4304
rect 53012 4264 53548 4304
rect 53588 4264 54932 4304
rect 54979 4264 54988 4304
rect 55028 4264 55604 4304
rect 56035 4264 56044 4304
rect 56084 4264 58348 4304
rect 58388 4264 58397 4304
rect 58732 4264 59500 4304
rect 59540 4264 59549 4304
rect 60163 4264 60172 4304
rect 60212 4264 65452 4304
rect 65492 4264 65501 4304
rect 65932 4304 65972 4348
rect 66883 4304 66941 4305
rect 67075 4304 67133 4305
rect 65932 4264 66892 4304
rect 66932 4264 66941 4304
rect 66990 4264 67084 4304
rect 67124 4264 67133 4304
rect 67267 4264 67276 4304
rect 67316 4264 67468 4304
rect 67508 4264 67517 4304
rect 67939 4264 67948 4304
rect 67988 4264 68332 4304
rect 68372 4264 68716 4304
rect 68756 4264 68908 4304
rect 68948 4264 68957 4304
rect 31651 4263 31709 4264
rect 19555 4220 19613 4221
rect 20227 4220 20285 4221
rect 23779 4220 23837 4221
rect 24931 4220 24989 4221
rect 28387 4220 28445 4221
rect 29923 4220 29981 4221
rect 49123 4220 49181 4221
rect 49516 4220 49556 4264
rect 49603 4220 49661 4221
rect 54892 4220 54932 4264
rect 2659 4180 2668 4220
rect 2708 4180 11020 4220
rect 11060 4180 11069 4220
rect 14563 4180 14572 4220
rect 14612 4180 17644 4220
rect 17684 4180 17693 4220
rect 19470 4180 19564 4220
rect 19604 4180 19613 4220
rect 20136 4180 20145 4220
rect 20185 4180 20236 4220
rect 20276 4180 20285 4220
rect 20515 4180 20524 4220
rect 20564 4180 21196 4220
rect 21236 4180 21245 4220
rect 21475 4180 21484 4220
rect 21524 4180 21868 4220
rect 21908 4180 21917 4220
rect 22243 4180 22252 4220
rect 22292 4180 22636 4220
rect 22676 4180 22685 4220
rect 22915 4180 22924 4220
rect 22964 4180 23596 4220
rect 23636 4180 23645 4220
rect 23694 4180 23788 4220
rect 23828 4180 23837 4220
rect 23971 4180 23980 4220
rect 24020 4180 24172 4220
rect 24212 4180 24221 4220
rect 24931 4180 24940 4220
rect 24980 4180 26860 4220
rect 26900 4180 26909 4220
rect 27427 4180 27436 4220
rect 27476 4180 27628 4220
rect 27668 4180 28012 4220
rect 28052 4180 28061 4220
rect 28387 4180 28396 4220
rect 28436 4180 28780 4220
rect 28820 4180 28829 4220
rect 29838 4180 29932 4220
rect 29972 4180 29981 4220
rect 30115 4180 30124 4220
rect 30164 4180 30316 4220
rect 30356 4180 30892 4220
rect 30932 4180 31276 4220
rect 31316 4180 31660 4220
rect 31700 4180 31709 4220
rect 33859 4180 33868 4220
rect 33908 4180 34444 4220
rect 34484 4180 34732 4220
rect 34772 4180 35020 4220
rect 35060 4180 35500 4220
rect 35540 4180 35549 4220
rect 37795 4180 37804 4220
rect 37844 4180 38188 4220
rect 38228 4180 38572 4220
rect 38612 4180 38956 4220
rect 38996 4180 39340 4220
rect 39380 4180 39389 4220
rect 41560 4180 43508 4220
rect 44611 4180 44620 4220
rect 44660 4180 45580 4220
rect 45620 4180 45629 4220
rect 47107 4180 47116 4220
rect 47156 4180 47308 4220
rect 47348 4180 49132 4220
rect 49172 4180 49181 4220
rect 49507 4180 49516 4220
rect 49556 4180 49612 4220
rect 49652 4180 49680 4220
rect 49987 4180 49996 4220
rect 50036 4180 50324 4220
rect 52099 4180 52108 4220
rect 52148 4180 52396 4220
rect 52436 4180 52684 4220
rect 52724 4180 52876 4220
rect 52916 4180 53356 4220
rect 53396 4180 53405 4220
rect 53452 4180 54796 4220
rect 54836 4180 54845 4220
rect 54892 4180 55084 4220
rect 55124 4180 55133 4220
rect 19555 4179 19613 4180
rect 20227 4179 20285 4180
rect 23779 4179 23837 4180
rect 24931 4179 24989 4180
rect 28387 4179 28445 4180
rect 29923 4179 29981 4180
rect 7075 4136 7133 4137
rect 12067 4136 12125 4137
rect 25699 4136 25757 4137
rect 30595 4136 30653 4137
rect 32899 4136 32957 4137
rect 34051 4136 34109 4137
rect 39043 4136 39101 4137
rect 41443 4136 41501 4137
rect 4579 4096 4588 4136
rect 4628 4096 7084 4136
rect 7124 4096 7133 4136
rect 7267 4096 7276 4136
rect 7316 4096 10540 4136
rect 10580 4096 10589 4136
rect 11107 4096 11116 4136
rect 11156 4096 12076 4136
rect 12116 4096 12125 4136
rect 7075 4095 7133 4096
rect 12067 4095 12125 4096
rect 14188 4096 14764 4136
rect 14804 4096 14813 4136
rect 18115 4096 18124 4136
rect 18164 4096 21812 4136
rect 14188 3968 14228 4096
rect 17155 4052 17213 4053
rect 21772 4052 21812 4096
rect 21964 4096 24268 4136
rect 24308 4096 24317 4136
rect 25614 4096 25708 4136
rect 25748 4096 25757 4136
rect 27715 4096 27724 4136
rect 27764 4096 28396 4136
rect 28436 4096 28445 4136
rect 28579 4096 28588 4136
rect 28628 4096 30548 4136
rect 21964 4052 22004 4096
rect 25699 4095 25757 4096
rect 23971 4052 24029 4053
rect 17155 4012 17164 4052
rect 17204 4012 17644 4052
rect 17684 4012 17693 4052
rect 17740 4012 21100 4052
rect 21140 4012 21149 4052
rect 21772 4012 22004 4052
rect 23886 4012 23980 4052
rect 24020 4012 24029 4052
rect 26083 4012 26092 4052
rect 26132 4012 28012 4052
rect 28052 4012 28061 4052
rect 28960 4012 29452 4052
rect 29492 4012 29501 4052
rect 17155 4011 17213 4012
rect 17740 3968 17780 4012
rect 23971 4011 24029 4012
rect 19747 3968 19805 3969
rect 4003 3928 4012 3968
rect 4052 3928 4204 3968
rect 4244 3928 4253 3968
rect 14179 3928 14188 3968
rect 14228 3928 14237 3968
rect 14755 3928 14764 3968
rect 14804 3928 16108 3968
rect 16148 3928 16157 3968
rect 16579 3928 16588 3968
rect 16628 3928 16876 3968
rect 16916 3928 16925 3968
rect 17644 3928 17780 3968
rect 19662 3928 19756 3968
rect 19796 3928 19805 3968
rect 17644 3884 17684 3928
rect 19747 3927 19805 3928
rect 19939 3968 19997 3969
rect 28960 3968 29000 4012
rect 19939 3928 19948 3968
rect 19988 3928 20082 3968
rect 20140 3928 24556 3968
rect 24596 3928 24605 3968
rect 27235 3928 27244 3968
rect 27284 3928 29000 3968
rect 29059 3968 29117 3969
rect 30508 3968 30548 4096
rect 30595 4096 30604 4136
rect 30644 4096 31988 4136
rect 32035 4096 32044 4136
rect 32084 4096 32716 4136
rect 32756 4096 32765 4136
rect 32899 4096 32908 4136
rect 32948 4096 33004 4136
rect 33044 4096 33053 4136
rect 33966 4096 34060 4136
rect 34100 4096 34109 4136
rect 34243 4096 34252 4136
rect 34292 4096 35116 4136
rect 35156 4096 35165 4136
rect 38755 4096 38764 4136
rect 38804 4096 39052 4136
rect 39092 4096 39101 4136
rect 40291 4096 40300 4136
rect 40340 4096 40588 4136
rect 40628 4096 40637 4136
rect 40867 4096 40876 4136
rect 40916 4096 41068 4136
rect 41108 4096 41117 4136
rect 41358 4096 41452 4136
rect 41492 4096 41501 4136
rect 30595 4095 30653 4096
rect 31948 4052 31988 4096
rect 32899 4095 32957 4096
rect 34051 4095 34109 4096
rect 39043 4095 39101 4096
rect 41443 4095 41501 4096
rect 41560 4052 41600 4180
rect 42595 4136 42653 4137
rect 42979 4136 43037 4137
rect 43363 4136 43421 4137
rect 42510 4096 42604 4136
rect 42644 4096 42653 4136
rect 42894 4096 42988 4136
rect 43028 4096 43037 4136
rect 43278 4096 43372 4136
rect 43412 4096 43421 4136
rect 43468 4136 43508 4180
rect 49123 4179 49181 4180
rect 49603 4179 49661 4180
rect 50284 4136 50324 4180
rect 53452 4136 53492 4180
rect 54115 4136 54173 4137
rect 43468 4096 46444 4136
rect 46484 4096 46493 4136
rect 50275 4096 50284 4136
rect 50324 4096 50956 4136
rect 50996 4096 52588 4136
rect 52628 4096 53492 4136
rect 54030 4096 54124 4136
rect 54164 4096 54173 4136
rect 54796 4136 54836 4180
rect 54796 4096 54988 4136
rect 55028 4096 55037 4136
rect 42595 4095 42653 4096
rect 42979 4095 43037 4096
rect 43363 4095 43421 4096
rect 54115 4095 54173 4096
rect 47299 4052 47357 4053
rect 55564 4052 55604 4264
rect 65443 4263 65501 4264
rect 66883 4263 66941 4264
rect 67075 4263 67133 4264
rect 57955 4220 58013 4221
rect 64771 4220 64829 4221
rect 69100 4220 69140 4348
rect 70435 4347 70493 4348
rect 71980 4304 72020 4432
rect 73027 4431 73085 4432
rect 77251 4431 77309 4432
rect 81763 4388 81821 4389
rect 85891 4388 85949 4389
rect 72259 4348 72268 4388
rect 72308 4348 73516 4388
rect 73556 4348 73565 4388
rect 75811 4348 75820 4388
rect 75860 4348 76588 4388
rect 76628 4348 76637 4388
rect 76771 4348 76780 4388
rect 76820 4348 77164 4388
rect 77204 4348 80908 4388
rect 80948 4348 80957 4388
rect 81678 4348 81772 4388
rect 81812 4348 83404 4388
rect 83444 4348 83692 4388
rect 83732 4348 83741 4388
rect 85891 4348 85900 4388
rect 85940 4348 86380 4388
rect 86420 4348 86429 4388
rect 81763 4347 81821 4348
rect 85891 4347 85949 4348
rect 69283 4264 69292 4304
rect 69332 4264 70060 4304
rect 70100 4264 70109 4304
rect 71980 4264 72788 4304
rect 74467 4264 74476 4304
rect 74516 4264 74668 4304
rect 74708 4264 75860 4304
rect 76387 4264 76396 4304
rect 76436 4264 77644 4304
rect 77684 4264 77693 4304
rect 79075 4264 79084 4304
rect 79124 4264 80620 4304
rect 80660 4264 80669 4304
rect 80995 4264 81004 4304
rect 81044 4264 81580 4304
rect 81620 4264 81629 4304
rect 83971 4264 83980 4304
rect 84020 4264 85324 4304
rect 85364 4264 85373 4304
rect 85699 4264 85708 4304
rect 85748 4264 86764 4304
rect 86804 4264 86813 4304
rect 89731 4264 89740 4304
rect 89780 4264 89932 4304
rect 89972 4264 89981 4304
rect 97795 4264 97804 4304
rect 97844 4264 98956 4304
rect 98996 4264 99005 4304
rect 72748 4220 72788 4264
rect 73411 4220 73469 4221
rect 75820 4220 75860 4264
rect 77539 4220 77597 4221
rect 56515 4180 56524 4220
rect 56564 4180 57100 4220
rect 57140 4180 57149 4220
rect 57870 4180 57964 4220
rect 58004 4180 58013 4220
rect 58819 4180 58828 4220
rect 58868 4180 59404 4220
rect 59444 4180 59453 4220
rect 59875 4180 59884 4220
rect 59924 4209 60596 4220
rect 59924 4180 60460 4209
rect 57955 4179 58013 4180
rect 60451 4169 60460 4180
rect 60500 4180 60596 4209
rect 62275 4180 62284 4220
rect 62324 4180 64588 4220
rect 64628 4180 64637 4220
rect 64686 4180 64780 4220
rect 64820 4180 64829 4220
rect 65635 4180 65644 4220
rect 65684 4180 68044 4220
rect 68084 4180 68093 4220
rect 68136 4180 68145 4220
rect 68185 4180 69140 4220
rect 70243 4180 70252 4220
rect 70292 4180 70444 4220
rect 70484 4180 70828 4220
rect 70868 4180 71212 4220
rect 71252 4180 71261 4220
rect 71779 4180 71788 4220
rect 71828 4180 72172 4220
rect 72212 4180 72221 4220
rect 72355 4180 72364 4220
rect 72404 4180 72692 4220
rect 72739 4180 72748 4220
rect 72788 4180 72797 4220
rect 73315 4180 73324 4220
rect 73364 4180 73420 4220
rect 73460 4180 75764 4220
rect 75811 4180 75820 4220
rect 75860 4180 75869 4220
rect 76003 4180 76012 4220
rect 76052 4180 76780 4220
rect 76820 4180 76829 4220
rect 77347 4180 77356 4220
rect 77396 4180 77548 4220
rect 77588 4180 77597 4220
rect 78403 4180 78412 4220
rect 78452 4180 81292 4220
rect 81332 4180 81341 4220
rect 81388 4180 84460 4220
rect 84500 4180 84509 4220
rect 86092 4180 95156 4220
rect 60500 4169 60509 4180
rect 56803 4136 56861 4137
rect 55651 4096 55660 4136
rect 55700 4096 56812 4136
rect 56852 4096 56861 4136
rect 58051 4096 58060 4136
rect 58100 4096 58540 4136
rect 58580 4096 58589 4136
rect 56803 4095 56861 4096
rect 60451 4052 60509 4053
rect 30883 4012 30892 4052
rect 30932 4012 31852 4052
rect 31892 4012 31901 4052
rect 31948 4012 34636 4052
rect 34676 4012 36172 4052
rect 36212 4012 36221 4052
rect 38563 4012 38572 4052
rect 38612 4012 41600 4052
rect 42787 4012 42796 4052
rect 42836 4012 45388 4052
rect 45428 4012 45437 4052
rect 46051 4012 46060 4052
rect 46100 4012 47308 4052
rect 47348 4012 47357 4052
rect 50179 4012 50188 4052
rect 50228 4012 51244 4052
rect 51284 4012 51293 4052
rect 51619 4012 51628 4052
rect 51668 4012 54796 4052
rect 54836 4012 54845 4052
rect 55564 4012 55988 4052
rect 56131 4012 56140 4052
rect 56180 4012 56524 4052
rect 56564 4012 57580 4052
rect 57620 4012 57629 4052
rect 57676 4012 60076 4052
rect 60116 4012 60125 4052
rect 60366 4012 60460 4052
rect 60500 4012 60509 4052
rect 47299 4011 47357 4012
rect 31267 3968 31325 3969
rect 49507 3968 49565 3969
rect 49699 3968 49757 3969
rect 29059 3928 29068 3968
rect 29108 3928 29261 3968
rect 29301 3928 29310 3968
rect 30508 3928 31276 3968
rect 31316 3928 31325 3968
rect 33571 3928 33580 3968
rect 33620 3928 35300 3968
rect 37795 3928 37804 3968
rect 37844 3928 37853 3968
rect 38179 3928 38188 3968
rect 38228 3928 38668 3968
rect 38708 3928 38717 3968
rect 39331 3928 39340 3968
rect 39380 3928 43028 3968
rect 43171 3928 43180 3968
rect 43220 3928 45772 3968
rect 45812 3928 45821 3968
rect 49219 3928 49228 3968
rect 49268 3928 49516 3968
rect 49556 3928 49565 3968
rect 49614 3928 49708 3968
rect 49748 3928 49757 3968
rect 52771 3928 52780 3968
rect 52820 3928 53740 3968
rect 53780 3928 53789 3968
rect 54019 3928 54028 3968
rect 54068 3928 55852 3968
rect 55892 3928 55901 3968
rect 19939 3927 19997 3928
rect 20140 3884 20180 3928
rect 29059 3927 29117 3928
rect 31267 3927 31325 3928
rect 35260 3884 35300 3928
rect 37804 3884 37844 3928
rect 42988 3884 43028 3928
rect 49507 3927 49565 3928
rect 49699 3927 49757 3928
rect 49891 3884 49949 3885
rect 55843 3884 55901 3885
rect 15043 3844 15052 3884
rect 15092 3844 17684 3884
rect 17731 3844 17740 3884
rect 17780 3844 20180 3884
rect 20419 3844 20428 3884
rect 20468 3844 21388 3884
rect 21428 3844 21437 3884
rect 22051 3844 22060 3884
rect 22100 3844 22540 3884
rect 22580 3844 25132 3884
rect 25172 3844 28492 3884
rect 28532 3844 30508 3884
rect 30548 3844 30557 3884
rect 35260 3844 35596 3884
rect 35636 3844 35645 3884
rect 37804 3844 42220 3884
rect 42260 3844 42269 3884
rect 42979 3844 42988 3884
rect 43028 3844 43037 3884
rect 49806 3844 49900 3884
rect 49940 3844 49949 3884
rect 53635 3844 53644 3884
rect 53684 3844 55852 3884
rect 55892 3844 55901 3884
rect 55948 3884 55988 4012
rect 56419 3928 56428 3968
rect 56468 3928 57388 3968
rect 57428 3928 57437 3968
rect 57676 3884 57716 4012
rect 60451 4011 60509 4012
rect 60556 3969 60596 4180
rect 64771 4179 64829 4180
rect 61987 4136 62045 4137
rect 66211 4136 66269 4137
rect 68611 4136 68669 4137
rect 68995 4136 69053 4137
rect 69475 4136 69533 4137
rect 61902 4096 61996 4136
rect 62036 4096 62045 4136
rect 66019 4096 66028 4136
rect 66068 4096 66220 4136
rect 66260 4096 66269 4136
rect 66403 4096 66412 4136
rect 66452 4096 68428 4136
rect 68468 4096 68477 4136
rect 68611 4096 68620 4136
rect 68660 4096 68669 4136
rect 68910 4096 69004 4136
rect 69044 4096 69053 4136
rect 69390 4096 69484 4136
rect 69524 4096 69533 4136
rect 61987 4095 62045 4096
rect 66211 4095 66269 4096
rect 68611 4095 68669 4096
rect 68995 4095 69053 4096
rect 69475 4095 69533 4096
rect 70435 4136 70493 4137
rect 72652 4136 72692 4180
rect 73411 4179 73469 4180
rect 75235 4136 75293 4137
rect 75619 4136 75677 4137
rect 70435 4096 70444 4136
rect 70484 4096 70580 4136
rect 71299 4096 71308 4136
rect 71348 4096 72556 4136
rect 72596 4096 72605 4136
rect 72652 4096 73132 4136
rect 73172 4096 73181 4136
rect 73324 4096 73900 4136
rect 73940 4096 73949 4136
rect 74371 4096 74380 4136
rect 74420 4096 75052 4136
rect 75092 4096 75101 4136
rect 75150 4096 75244 4136
rect 75284 4096 75293 4136
rect 75534 4096 75628 4136
rect 75668 4096 75677 4136
rect 75724 4136 75764 4180
rect 76012 4136 76052 4180
rect 77539 4179 77597 4180
rect 79747 4136 79805 4137
rect 81388 4136 81428 4180
rect 86092 4136 86132 4180
rect 75724 4096 76052 4136
rect 76099 4096 76108 4136
rect 76148 4096 76396 4136
rect 76436 4096 76445 4136
rect 76675 4096 76684 4136
rect 76724 4096 77164 4136
rect 77204 4096 78795 4136
rect 78835 4096 78844 4136
rect 78979 4096 78988 4136
rect 79028 4096 79756 4136
rect 79796 4096 79805 4136
rect 80035 4096 80044 4136
rect 80084 4096 80428 4136
rect 80468 4096 80477 4136
rect 80899 4096 80908 4136
rect 80948 4096 81428 4136
rect 81880 4096 82540 4136
rect 82580 4096 82589 4136
rect 82723 4096 82732 4136
rect 82772 4096 83212 4136
rect 83252 4096 83261 4136
rect 84355 4096 84364 4136
rect 84404 4096 86132 4136
rect 86275 4136 86333 4137
rect 95116 4136 95156 4180
rect 86275 4096 86284 4136
rect 86324 4096 86418 4136
rect 88387 4096 88396 4136
rect 88436 4096 88445 4136
rect 89827 4096 89836 4136
rect 89876 4096 91660 4136
rect 91700 4096 91709 4136
rect 93283 4096 93292 4136
rect 93332 4096 93868 4136
rect 93908 4096 93917 4136
rect 95107 4096 95116 4136
rect 95156 4096 95165 4136
rect 97219 4096 97228 4136
rect 97268 4096 98572 4136
rect 98612 4096 98621 4136
rect 70435 4095 70493 4096
rect 64771 4052 64829 4053
rect 60643 4012 60652 4052
rect 60692 4012 63628 4052
rect 63668 4012 63677 4052
rect 64686 4012 64780 4052
rect 64820 4012 64829 4052
rect 64771 4011 64829 4012
rect 66403 4052 66461 4053
rect 68620 4052 68660 4095
rect 70540 4052 70580 4096
rect 73324 4052 73364 4096
rect 75235 4095 75293 4096
rect 75619 4095 75677 4096
rect 79747 4095 79805 4096
rect 73507 4052 73565 4053
rect 75715 4052 75773 4053
rect 77251 4052 77309 4053
rect 81880 4052 81920 4096
rect 86275 4095 86333 4096
rect 66403 4012 66412 4052
rect 66452 4012 68524 4052
rect 68564 4012 68573 4052
rect 68620 4012 69100 4052
rect 69140 4012 69149 4052
rect 69571 4012 69580 4052
rect 69620 4012 70444 4052
rect 70484 4012 70493 4052
rect 70540 4012 70636 4052
rect 70676 4012 70685 4052
rect 71395 4012 71404 4052
rect 71444 4012 73364 4052
rect 73422 4012 73516 4052
rect 73556 4012 73565 4052
rect 74851 4012 74860 4052
rect 74900 4012 75532 4052
rect 75572 4012 75581 4052
rect 75715 4012 75724 4052
rect 75764 4012 77260 4052
rect 77300 4012 77309 4052
rect 66403 4011 66461 4012
rect 73507 4011 73565 4012
rect 75715 4011 75773 4012
rect 77251 4011 77309 4012
rect 77452 4012 81920 4052
rect 85123 4012 85132 4052
rect 85172 4012 85516 4052
rect 85556 4012 85565 4052
rect 60547 3968 60605 3969
rect 66883 3968 66941 3969
rect 70531 3968 70589 3969
rect 71779 3968 71837 3969
rect 77452 3968 77492 4012
rect 84259 3968 84317 3969
rect 88396 3968 88436 4096
rect 94243 4012 94252 4052
rect 94292 4012 94924 4052
rect 94964 4012 94973 4052
rect 60462 3928 60556 3968
rect 60596 3928 64280 3968
rect 64579 3928 64588 3968
rect 64628 3928 65836 3968
rect 65876 3928 65885 3968
rect 66211 3928 66220 3968
rect 66260 3928 66269 3968
rect 66883 3928 66892 3968
rect 66932 3928 68140 3968
rect 68180 3928 68189 3968
rect 70531 3928 70540 3968
rect 70580 3928 71020 3968
rect 71060 3928 71069 3968
rect 71694 3928 71788 3968
rect 71828 3928 71837 3968
rect 72163 3928 72172 3968
rect 72212 3928 77492 3968
rect 79555 3928 79564 3968
rect 79604 3928 79852 3968
rect 79892 3928 79901 3968
rect 80323 3928 80332 3968
rect 80372 3928 80381 3968
rect 82147 3928 82156 3968
rect 82196 3928 82444 3968
rect 82484 3928 82493 3968
rect 84259 3928 84268 3968
rect 84308 3928 84364 3968
rect 84404 3928 84413 3968
rect 85027 3928 85036 3968
rect 85076 3928 87244 3968
rect 87284 3928 87293 3968
rect 88195 3928 88204 3968
rect 88244 3928 88436 3968
rect 90787 3928 90796 3968
rect 90836 3928 91468 3968
rect 91508 3928 91517 3968
rect 91747 3928 91756 3968
rect 91796 3928 92236 3968
rect 92276 3928 92285 3968
rect 94051 3928 94060 3968
rect 94100 3928 94540 3968
rect 94580 3928 94589 3968
rect 94723 3928 94732 3968
rect 94772 3928 94781 3968
rect 96163 3928 96172 3968
rect 96212 3928 96844 3968
rect 96884 3928 96893 3968
rect 98371 3928 98380 3968
rect 98420 3928 98764 3968
rect 98804 3928 98813 3968
rect 60547 3927 60605 3928
rect 58531 3884 58589 3885
rect 62083 3884 62141 3885
rect 64240 3884 64280 3928
rect 66220 3884 66260 3928
rect 66883 3927 66941 3928
rect 70531 3927 70589 3928
rect 55948 3844 57716 3884
rect 58446 3844 58540 3884
rect 58580 3844 58589 3884
rect 61998 3844 62092 3884
rect 62132 3844 62141 3884
rect 63043 3844 63052 3884
rect 63092 3844 63340 3884
rect 63380 3844 63389 3884
rect 64240 3844 64684 3884
rect 64724 3844 64733 3884
rect 64867 3844 64876 3884
rect 64916 3844 66260 3884
rect 66787 3884 66845 3885
rect 68227 3884 68285 3885
rect 70723 3884 70781 3885
rect 66787 3844 66796 3884
rect 66836 3844 67756 3884
rect 67796 3844 67805 3884
rect 68227 3844 68236 3884
rect 68276 3844 70580 3884
rect 70627 3844 70636 3884
rect 70676 3844 70732 3884
rect 70772 3844 70781 3884
rect 71020 3884 71060 3928
rect 71779 3927 71837 3928
rect 75139 3884 75197 3885
rect 80332 3884 80372 3928
rect 84259 3927 84317 3928
rect 86851 3884 86909 3885
rect 94732 3884 94772 3928
rect 71020 3844 75092 3884
rect 49891 3843 49949 3844
rect 55843 3843 55901 3844
rect 58531 3843 58589 3844
rect 62083 3843 62141 3844
rect 66787 3843 66845 3844
rect 68227 3843 68285 3844
rect 23875 3800 23933 3801
rect 35587 3800 35645 3801
rect 38083 3800 38141 3801
rect 40291 3800 40349 3801
rect 41059 3800 41117 3801
rect 57091 3800 57149 3801
rect 67075 3800 67133 3801
rect 67843 3800 67901 3801
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4675 3760 4684 3800
rect 4724 3760 7372 3800
rect 7412 3760 7421 3800
rect 15139 3760 15148 3800
rect 15188 3760 15628 3800
rect 15668 3760 15677 3800
rect 15907 3760 15916 3800
rect 15956 3760 17548 3800
rect 17588 3760 17597 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 22435 3760 22444 3800
rect 22484 3760 23884 3800
rect 23924 3760 23933 3800
rect 24643 3760 24652 3800
rect 24692 3760 27628 3800
rect 27668 3760 27677 3800
rect 28675 3760 28684 3800
rect 28724 3760 29260 3800
rect 29300 3760 29309 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 35299 3760 35308 3800
rect 35348 3760 35596 3800
rect 35636 3760 35645 3800
rect 35875 3760 35884 3800
rect 35924 3760 36844 3800
rect 36884 3760 36893 3800
rect 38083 3760 38092 3800
rect 38132 3760 38764 3800
rect 38804 3760 38813 3800
rect 40206 3760 40300 3800
rect 40340 3760 40349 3800
rect 40974 3760 41068 3800
rect 41108 3760 41117 3800
rect 41251 3760 41260 3800
rect 41300 3760 43276 3800
rect 43316 3760 43325 3800
rect 43555 3760 43564 3800
rect 43604 3760 46156 3800
rect 46196 3760 46205 3800
rect 46819 3760 46828 3800
rect 46868 3760 47500 3800
rect 47540 3760 47549 3800
rect 49039 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49425 3800
rect 49507 3760 49516 3800
rect 49556 3760 50092 3800
rect 50132 3760 50141 3800
rect 50188 3760 52628 3800
rect 52867 3760 52876 3800
rect 52916 3760 54124 3800
rect 54164 3760 54173 3800
rect 55267 3760 55276 3800
rect 55316 3760 57100 3800
rect 57140 3760 57149 3800
rect 58243 3760 58252 3800
rect 58292 3760 58732 3800
rect 58772 3760 58781 3800
rect 60643 3760 60652 3800
rect 60692 3760 62572 3800
rect 62612 3760 62621 3800
rect 64159 3760 64168 3800
rect 64208 3760 64250 3800
rect 64290 3760 64332 3800
rect 64372 3760 64414 3800
rect 64454 3760 64496 3800
rect 64536 3760 64545 3800
rect 64771 3760 64780 3800
rect 64820 3760 65260 3800
rect 65300 3760 65309 3800
rect 65443 3760 65452 3800
rect 65492 3760 65932 3800
rect 65972 3760 65981 3800
rect 66990 3760 67084 3800
rect 67124 3760 67133 3800
rect 67758 3760 67852 3800
rect 67892 3760 67901 3800
rect 23875 3759 23933 3760
rect 35587 3759 35645 3760
rect 38083 3759 38141 3760
rect 40291 3759 40349 3760
rect 41059 3759 41117 3760
rect 14467 3716 14525 3717
rect 16387 3716 16445 3717
rect 20131 3716 20189 3717
rect 14467 3676 14476 3716
rect 14516 3676 15052 3716
rect 15092 3676 15101 3716
rect 15427 3676 15436 3716
rect 15476 3676 15724 3716
rect 15764 3676 15773 3716
rect 16387 3676 16396 3716
rect 16436 3676 20140 3716
rect 20180 3676 20189 3716
rect 14467 3675 14525 3676
rect 16387 3675 16445 3676
rect 20131 3675 20189 3676
rect 20323 3716 20381 3717
rect 20611 3716 20669 3717
rect 24451 3716 24509 3717
rect 50188 3716 50228 3760
rect 20323 3676 20332 3716
rect 20372 3676 20620 3716
rect 20660 3676 20669 3716
rect 20899 3676 20908 3716
rect 20948 3676 23116 3716
rect 23156 3676 23165 3716
rect 24451 3676 24460 3716
rect 24500 3676 28492 3716
rect 28532 3676 28541 3716
rect 30499 3676 30508 3716
rect 30548 3676 35020 3716
rect 35060 3676 37996 3716
rect 38036 3676 43468 3716
rect 43508 3676 43517 3716
rect 48547 3676 48556 3716
rect 48596 3676 50228 3716
rect 52195 3676 52204 3716
rect 52244 3676 52492 3716
rect 52532 3676 52541 3716
rect 20323 3675 20381 3676
rect 20611 3675 20669 3676
rect 24451 3675 24509 3676
rect 25411 3632 25469 3633
rect 11971 3592 11980 3632
rect 12020 3592 22348 3632
rect 22388 3592 22397 3632
rect 22723 3592 22732 3632
rect 22772 3592 23884 3632
rect 23924 3592 23933 3632
rect 25326 3592 25420 3632
rect 25460 3592 25469 3632
rect 25411 3591 25469 3592
rect 26371 3632 26429 3633
rect 26371 3592 26380 3632
rect 26420 3592 26572 3632
rect 26612 3592 26621 3632
rect 31939 3592 31948 3632
rect 31988 3592 31997 3632
rect 33091 3592 33100 3632
rect 33140 3592 34252 3632
rect 34292 3592 34301 3632
rect 35107 3592 35116 3632
rect 35156 3592 39052 3632
rect 39092 3592 39101 3632
rect 39523 3592 39532 3632
rect 39572 3592 42604 3632
rect 42644 3592 42653 3632
rect 42883 3592 42892 3632
rect 42932 3592 46732 3632
rect 46772 3592 46781 3632
rect 48931 3592 48940 3632
rect 48980 3592 49420 3632
rect 49460 3592 49469 3632
rect 26371 3591 26429 3592
rect 19843 3548 19901 3549
rect 20899 3548 20957 3549
rect 21571 3548 21629 3549
rect 31948 3548 31988 3592
rect 52588 3548 52628 3760
rect 57091 3759 57149 3760
rect 67075 3759 67133 3760
rect 67843 3759 67901 3760
rect 68323 3800 68381 3801
rect 70540 3800 70580 3844
rect 70723 3843 70781 3844
rect 75052 3800 75092 3844
rect 75139 3844 75148 3884
rect 75188 3844 75628 3884
rect 75668 3844 75677 3884
rect 77059 3844 77068 3884
rect 77108 3844 77204 3884
rect 78019 3844 78028 3884
rect 78068 3844 80372 3884
rect 80611 3844 80620 3884
rect 80660 3844 85900 3884
rect 85940 3844 85949 3884
rect 86851 3844 86860 3884
rect 86900 3844 94772 3884
rect 75139 3843 75197 3844
rect 75331 3800 75389 3801
rect 77059 3800 77117 3801
rect 68323 3760 68332 3800
rect 68372 3760 70060 3800
rect 70100 3760 70109 3800
rect 70540 3760 71404 3800
rect 71444 3760 71453 3800
rect 71971 3760 71980 3800
rect 72020 3760 73900 3800
rect 73940 3760 73949 3800
rect 75052 3760 75340 3800
rect 75380 3760 75389 3800
rect 75523 3760 75532 3800
rect 75572 3760 77068 3800
rect 77108 3760 77117 3800
rect 77164 3800 77204 3844
rect 86851 3843 86909 3844
rect 79747 3800 79805 3801
rect 81475 3800 81533 3801
rect 77164 3760 77740 3800
rect 77780 3760 77789 3800
rect 78211 3760 78220 3800
rect 78260 3760 78988 3800
rect 79028 3760 79037 3800
rect 79279 3760 79288 3800
rect 79328 3760 79370 3800
rect 79410 3760 79452 3800
rect 79492 3760 79534 3800
rect 79574 3760 79616 3800
rect 79656 3760 79665 3800
rect 79747 3760 79756 3800
rect 79796 3760 80716 3800
rect 80756 3760 81196 3800
rect 81236 3760 81245 3800
rect 81475 3760 81484 3800
rect 81524 3760 83596 3800
rect 83636 3760 83645 3800
rect 84451 3760 84460 3800
rect 84500 3760 86860 3800
rect 86900 3760 86909 3800
rect 91939 3760 91948 3800
rect 91988 3760 92620 3800
rect 92660 3760 92669 3800
rect 92899 3760 92908 3800
rect 92948 3760 93388 3800
rect 93428 3760 93437 3800
rect 94399 3760 94408 3800
rect 94448 3760 94490 3800
rect 94530 3760 94572 3800
rect 94612 3760 94654 3800
rect 94694 3760 94736 3800
rect 94776 3760 94785 3800
rect 95587 3760 95596 3800
rect 95636 3760 96076 3800
rect 96116 3760 96125 3800
rect 68323 3759 68381 3760
rect 75331 3759 75389 3760
rect 77059 3759 77117 3760
rect 79747 3759 79805 3760
rect 81475 3759 81533 3760
rect 63811 3716 63869 3717
rect 80611 3716 80669 3717
rect 53347 3676 53356 3716
rect 53396 3676 61132 3716
rect 61172 3676 61181 3716
rect 61507 3676 61516 3716
rect 61556 3676 63572 3716
rect 63427 3632 63485 3633
rect 54787 3592 54796 3632
rect 54836 3592 55372 3632
rect 55412 3592 55421 3632
rect 56035 3592 56044 3632
rect 56084 3592 58156 3632
rect 58196 3592 58205 3632
rect 59683 3592 59692 3632
rect 59732 3592 63436 3632
rect 63476 3592 63485 3632
rect 63427 3591 63485 3592
rect 60259 3548 60317 3549
rect 8140 3508 18604 3548
rect 18644 3508 18653 3548
rect 18883 3508 18892 3548
rect 18932 3508 19372 3548
rect 19412 3508 19421 3548
rect 19843 3508 19852 3548
rect 19892 3508 20180 3548
rect 20515 3508 20524 3548
rect 20564 3508 20908 3548
rect 20948 3508 20957 3548
rect 21486 3508 21580 3548
rect 21620 3508 21629 3548
rect 21763 3508 21772 3548
rect 21812 3508 22636 3548
rect 22676 3508 22685 3548
rect 26659 3508 26668 3548
rect 26708 3508 27668 3548
rect 31948 3508 33716 3548
rect 34915 3508 34924 3548
rect 34964 3508 40588 3548
rect 40628 3508 40637 3548
rect 40867 3508 40876 3548
rect 40916 3508 41356 3548
rect 41396 3508 41405 3548
rect 42019 3508 42028 3548
rect 42068 3508 44332 3548
rect 44372 3508 44381 3548
rect 48163 3508 48172 3548
rect 48212 3508 49036 3548
rect 49076 3508 49085 3548
rect 51427 3508 51436 3548
rect 51476 3508 52492 3548
rect 52532 3508 52541 3548
rect 52588 3508 59212 3548
rect 59252 3508 59261 3548
rect 60174 3508 60268 3548
rect 60308 3508 60317 3548
rect 61219 3508 61228 3548
rect 61268 3508 62284 3548
rect 62324 3508 62333 3548
rect 1219 3464 1277 3465
rect 1603 3464 1661 3465
rect 1987 3464 2045 3465
rect 2371 3464 2429 3465
rect 6211 3464 6269 3465
rect 6979 3464 7037 3465
rect 8140 3464 8180 3508
rect 19843 3507 19901 3508
rect 16195 3464 16253 3465
rect 17155 3464 17213 3465
rect 17443 3464 17501 3465
rect 18499 3464 18557 3465
rect 19267 3464 19325 3465
rect 20140 3464 20180 3508
rect 20899 3507 20957 3508
rect 21571 3507 21629 3508
rect 21955 3464 22013 3465
rect 22147 3464 22205 3465
rect 23491 3464 23549 3465
rect 27628 3464 27668 3508
rect 28099 3464 28157 3465
rect 31939 3464 31997 3465
rect 1134 3424 1228 3464
rect 1268 3424 1277 3464
rect 1518 3424 1612 3464
rect 1652 3424 1661 3464
rect 1902 3424 1996 3464
rect 2036 3424 2045 3464
rect 2286 3424 2380 3464
rect 2420 3424 2429 3464
rect 3331 3424 3340 3464
rect 3380 3424 3532 3464
rect 3572 3424 3581 3464
rect 4291 3424 4300 3464
rect 4340 3424 6220 3464
rect 6260 3424 6269 3464
rect 6894 3424 6988 3464
rect 7028 3424 7037 3464
rect 8131 3424 8140 3464
rect 8180 3424 8189 3464
rect 10051 3424 10060 3464
rect 10100 3424 15764 3464
rect 15811 3424 15820 3464
rect 15860 3424 16204 3464
rect 16244 3424 16253 3464
rect 16771 3424 16780 3464
rect 16820 3424 16972 3464
rect 17012 3424 17021 3464
rect 17155 3424 17164 3464
rect 17204 3424 17298 3464
rect 17347 3424 17356 3464
rect 17396 3424 17452 3464
rect 17492 3424 17501 3464
rect 18414 3424 18508 3464
rect 18548 3424 18557 3464
rect 19182 3424 19276 3464
rect 19316 3424 19325 3464
rect 20035 3424 20044 3464
rect 20084 3424 20093 3464
rect 20140 3424 21196 3464
rect 21236 3424 21245 3464
rect 21955 3424 21964 3464
rect 22004 3424 22098 3464
rect 22147 3424 22156 3464
rect 22196 3424 23116 3464
rect 23156 3424 23165 3464
rect 23406 3424 23500 3464
rect 23540 3424 23549 3464
rect 25411 3424 25420 3464
rect 25460 3424 27436 3464
rect 27476 3424 27485 3464
rect 27619 3424 27628 3464
rect 27668 3424 27677 3464
rect 28014 3424 28108 3464
rect 28148 3424 28157 3464
rect 29635 3424 29644 3464
rect 29684 3424 30316 3464
rect 30356 3424 30365 3464
rect 31854 3424 31948 3464
rect 31988 3424 31997 3464
rect 1219 3423 1277 3424
rect 1603 3423 1661 3424
rect 1987 3423 2045 3424
rect 2371 3423 2429 3424
rect 6211 3423 6269 3424
rect 6979 3423 7037 3424
rect 1027 3340 1036 3380
rect 1076 3340 2572 3380
rect 2612 3340 2621 3380
rect 14371 3340 14380 3380
rect 14420 3340 14764 3380
rect 14804 3340 14813 3380
rect 15724 3296 15764 3424
rect 16195 3423 16253 3424
rect 17155 3423 17213 3424
rect 17443 3423 17501 3424
rect 18499 3423 18557 3424
rect 19267 3423 19325 3424
rect 18691 3380 18749 3381
rect 15907 3340 15916 3380
rect 15956 3340 18700 3380
rect 18740 3340 18749 3380
rect 20044 3380 20084 3424
rect 21955 3423 22013 3424
rect 22147 3423 22205 3424
rect 23491 3423 23549 3424
rect 28099 3423 28157 3424
rect 31939 3423 31997 3424
rect 32131 3464 32189 3465
rect 33676 3464 33716 3508
rect 60259 3507 60317 3508
rect 36067 3464 36125 3465
rect 32131 3424 32140 3464
rect 32180 3424 33580 3464
rect 33620 3424 33629 3464
rect 33676 3424 35692 3464
rect 35732 3424 35741 3464
rect 35982 3424 36076 3464
rect 36116 3424 36125 3464
rect 32131 3423 32189 3424
rect 36067 3423 36125 3424
rect 36547 3464 36605 3465
rect 43363 3464 43421 3465
rect 47971 3464 48029 3465
rect 56899 3464 56957 3465
rect 36547 3424 36556 3464
rect 36596 3424 38380 3464
rect 38420 3424 38429 3464
rect 38947 3424 38956 3464
rect 38996 3424 41836 3464
rect 41876 3424 41885 3464
rect 43278 3424 43372 3464
rect 43412 3424 43421 3464
rect 44707 3424 44716 3464
rect 44756 3424 44765 3464
rect 47886 3424 47980 3464
rect 48020 3424 48029 3464
rect 49123 3424 49132 3464
rect 49172 3424 49652 3464
rect 51811 3424 51820 3464
rect 51860 3424 52396 3464
rect 52436 3424 52445 3464
rect 56814 3424 56908 3464
rect 56948 3424 56957 3464
rect 36547 3423 36605 3424
rect 43363 3423 43421 3424
rect 30019 3380 30077 3381
rect 34339 3380 34397 3381
rect 20044 3340 23308 3380
rect 23348 3340 23357 3380
rect 25987 3340 25996 3380
rect 26036 3340 26045 3380
rect 26179 3340 26188 3380
rect 26228 3340 26380 3380
rect 26420 3340 26429 3380
rect 29934 3340 30028 3380
rect 30068 3340 30077 3380
rect 31747 3340 31756 3380
rect 31796 3340 33100 3380
rect 33140 3340 33149 3380
rect 34339 3340 34348 3380
rect 34388 3340 37364 3380
rect 37411 3340 37420 3380
rect 37460 3340 38860 3380
rect 38900 3340 38909 3380
rect 40483 3340 40492 3380
rect 40532 3340 42124 3380
rect 42164 3340 42173 3380
rect 43939 3340 43948 3380
rect 43988 3340 44620 3380
rect 44660 3340 44669 3380
rect 18691 3339 18749 3340
rect 20323 3296 20381 3297
rect 7747 3256 7756 3296
rect 7796 3256 9620 3296
rect 10819 3256 10828 3296
rect 10868 3256 15148 3296
rect 15188 3256 15197 3296
rect 15724 3256 20332 3296
rect 20372 3256 20381 3296
rect 9580 3212 9620 3256
rect 20323 3255 20381 3256
rect 20803 3296 20861 3297
rect 25996 3296 26036 3340
rect 30019 3339 30077 3340
rect 34339 3339 34397 3340
rect 20803 3256 20812 3296
rect 20852 3256 20946 3296
rect 25996 3256 27724 3296
rect 27764 3256 27773 3296
rect 34636 3256 35788 3296
rect 35828 3256 35837 3296
rect 36931 3256 36940 3296
rect 36980 3256 37228 3296
rect 37268 3256 37277 3296
rect 20803 3255 20861 3256
rect 20707 3212 20765 3213
rect 1411 3172 1420 3212
rect 1460 3172 1612 3212
rect 1652 3172 1661 3212
rect 2179 3172 2188 3212
rect 2228 3172 2380 3212
rect 2420 3172 2429 3212
rect 2563 3172 2572 3212
rect 2612 3172 3628 3212
rect 3668 3172 3677 3212
rect 4675 3172 4684 3212
rect 4724 3172 4876 3212
rect 4916 3172 4925 3212
rect 5251 3172 5260 3212
rect 5300 3172 5740 3212
rect 5780 3172 5789 3212
rect 7555 3172 7564 3212
rect 7604 3172 8524 3212
rect 8564 3172 8573 3212
rect 9580 3172 14036 3212
rect 14083 3172 14092 3212
rect 14132 3172 14380 3212
rect 14420 3172 14429 3212
rect 15427 3172 15436 3212
rect 15476 3172 15916 3212
rect 15956 3172 15965 3212
rect 17155 3172 17164 3212
rect 17204 3172 19660 3212
rect 19700 3172 19709 3212
rect 20227 3172 20236 3212
rect 20276 3172 20716 3212
rect 20756 3172 20765 3212
rect 20995 3172 21004 3212
rect 21044 3172 23116 3212
rect 23156 3172 23165 3212
rect 25219 3172 25228 3212
rect 25268 3172 26956 3212
rect 26996 3172 27005 3212
rect 27907 3172 27916 3212
rect 27956 3172 29000 3212
rect 30211 3172 30220 3212
rect 30260 3172 31564 3212
rect 31604 3172 31613 3212
rect 13996 3128 14036 3172
rect 20707 3171 20765 3172
rect 20899 3128 20957 3129
rect 3235 3088 3244 3128
rect 3284 3088 3532 3128
rect 3572 3088 3581 3128
rect 7363 3088 7372 3128
rect 7412 3088 8372 3128
rect 10435 3088 10444 3128
rect 10484 3088 13900 3128
rect 13940 3088 13949 3128
rect 13996 3088 17260 3128
rect 17300 3088 17309 3128
rect 20814 3088 20908 3128
rect 20948 3088 20957 3128
rect 28960 3128 29000 3172
rect 34636 3128 34676 3256
rect 35491 3172 35500 3212
rect 35540 3172 36980 3212
rect 28960 3088 30316 3128
rect 30356 3088 30365 3128
rect 31267 3088 31276 3128
rect 31316 3088 34676 3128
rect 34723 3128 34781 3129
rect 36940 3128 36980 3172
rect 37324 3128 37364 3340
rect 37795 3296 37853 3297
rect 39715 3296 39773 3297
rect 44716 3296 44756 3424
rect 47971 3423 48029 3424
rect 45091 3340 45100 3380
rect 45140 3340 46252 3380
rect 46292 3340 46301 3380
rect 49315 3340 49324 3380
rect 49364 3340 49516 3380
rect 49556 3340 49565 3380
rect 49612 3297 49652 3424
rect 56899 3423 56957 3424
rect 57379 3464 57437 3465
rect 58147 3464 58205 3465
rect 60739 3464 60797 3465
rect 63532 3464 63572 3676
rect 63811 3676 63820 3716
rect 63860 3676 64972 3716
rect 65012 3676 65021 3716
rect 66211 3676 66220 3716
rect 66260 3676 66700 3716
rect 66740 3676 66749 3716
rect 68131 3676 68140 3716
rect 68180 3676 68524 3716
rect 68564 3676 68573 3716
rect 68620 3676 80620 3716
rect 80660 3676 80669 3716
rect 82243 3676 82252 3716
rect 82292 3676 82444 3716
rect 82484 3676 82493 3716
rect 83395 3676 83404 3716
rect 83444 3676 98188 3716
rect 98228 3676 98237 3716
rect 63811 3675 63869 3676
rect 63715 3632 63773 3633
rect 68620 3632 68660 3676
rect 80611 3675 80669 3676
rect 76579 3632 76637 3633
rect 81859 3632 81917 3633
rect 63715 3592 63724 3632
rect 63764 3592 68660 3632
rect 70147 3592 70156 3632
rect 70196 3592 70924 3632
rect 70964 3592 70973 3632
rect 71779 3592 71788 3632
rect 71828 3592 73132 3632
rect 73172 3592 73181 3632
rect 73507 3592 73516 3632
rect 73556 3592 75436 3632
rect 75476 3592 75485 3632
rect 76579 3592 76588 3632
rect 76628 3592 76684 3632
rect 76724 3592 76733 3632
rect 77347 3592 77356 3632
rect 77396 3592 78700 3632
rect 78740 3592 78749 3632
rect 79180 3592 81868 3632
rect 81908 3592 81917 3632
rect 83203 3592 83212 3632
rect 83252 3592 84940 3632
rect 84980 3592 84989 3632
rect 85123 3592 85132 3632
rect 85172 3592 87052 3632
rect 87092 3592 87101 3632
rect 93091 3592 93100 3632
rect 93140 3592 93772 3632
rect 93812 3592 93821 3632
rect 97411 3592 97420 3632
rect 97460 3592 98860 3632
rect 98900 3592 98909 3632
rect 63715 3591 63773 3592
rect 76579 3591 76637 3592
rect 79180 3548 79220 3592
rect 81859 3591 81917 3592
rect 63907 3508 63916 3548
rect 63956 3508 64972 3548
rect 65012 3508 65021 3548
rect 66307 3508 66316 3548
rect 66356 3508 70100 3548
rect 70243 3508 70252 3548
rect 70292 3508 72076 3548
rect 72116 3508 72125 3548
rect 73699 3508 73708 3548
rect 73748 3508 78220 3548
rect 78260 3508 78269 3548
rect 78508 3508 79220 3548
rect 79267 3508 79276 3548
rect 79316 3508 82636 3548
rect 82676 3508 82685 3548
rect 82915 3508 82924 3548
rect 82964 3508 86860 3548
rect 86900 3508 86909 3548
rect 87139 3508 87148 3548
rect 87188 3508 87820 3548
rect 87860 3508 87869 3548
rect 87916 3508 90740 3548
rect 91171 3508 91180 3548
rect 91220 3508 91852 3548
rect 91892 3508 91901 3548
rect 67459 3464 67517 3465
rect 69379 3464 69437 3465
rect 57379 3424 57388 3464
rect 57428 3424 57772 3464
rect 57812 3424 57821 3464
rect 58062 3424 58156 3464
rect 58196 3424 58205 3464
rect 60654 3424 60748 3464
rect 60788 3424 60797 3464
rect 57379 3423 57437 3424
rect 58147 3423 58205 3424
rect 60739 3423 60797 3424
rect 61720 3424 63244 3464
rect 63284 3424 63293 3464
rect 63532 3424 65164 3464
rect 65204 3424 65213 3464
rect 65923 3424 65932 3464
rect 65972 3424 66988 3464
rect 67028 3424 67037 3464
rect 67374 3424 67468 3464
rect 67508 3424 67517 3464
rect 69294 3424 69388 3464
rect 69428 3424 69437 3464
rect 70060 3464 70100 3508
rect 70339 3464 70397 3465
rect 76291 3464 76349 3465
rect 70060 3424 70348 3464
rect 70388 3424 70397 3464
rect 74179 3424 74188 3464
rect 74228 3424 75148 3464
rect 75188 3424 75197 3464
rect 76206 3424 76300 3464
rect 76340 3424 76349 3464
rect 61720 3380 61760 3424
rect 67459 3423 67517 3424
rect 69379 3423 69437 3424
rect 70339 3423 70397 3424
rect 76291 3423 76349 3424
rect 76771 3464 76829 3465
rect 78508 3464 78548 3508
rect 80131 3464 80189 3465
rect 87916 3464 87956 3508
rect 89251 3464 89309 3465
rect 76771 3424 76780 3464
rect 76820 3424 78548 3464
rect 78595 3424 78604 3464
rect 78644 3424 78653 3464
rect 78787 3424 78796 3464
rect 78836 3424 79372 3464
rect 79412 3424 79421 3464
rect 80046 3424 80140 3464
rect 80180 3424 80189 3464
rect 80515 3424 80524 3464
rect 80564 3424 81100 3464
rect 81140 3424 81149 3464
rect 82051 3424 82060 3464
rect 82100 3424 82828 3464
rect 82868 3424 82877 3464
rect 83875 3424 83884 3464
rect 83924 3424 87956 3464
rect 88579 3424 88588 3464
rect 88628 3424 89260 3464
rect 89300 3424 89309 3464
rect 90700 3464 90740 3508
rect 94723 3464 94781 3465
rect 95107 3464 95165 3465
rect 95491 3464 95549 3465
rect 95875 3464 95933 3465
rect 96643 3464 96701 3465
rect 97411 3464 97469 3465
rect 97795 3464 97853 3465
rect 90700 3424 91660 3464
rect 91700 3424 91709 3464
rect 92035 3424 92044 3464
rect 92084 3424 92093 3464
rect 94638 3424 94732 3464
rect 94772 3424 94781 3464
rect 95022 3424 95116 3464
rect 95156 3424 95165 3464
rect 95406 3424 95500 3464
rect 95540 3424 95549 3464
rect 95790 3424 95884 3464
rect 95924 3424 95933 3464
rect 96558 3424 96652 3464
rect 96692 3424 96701 3464
rect 97326 3424 97420 3464
rect 97460 3424 97469 3464
rect 97710 3424 97804 3464
rect 97844 3424 97853 3464
rect 76771 3423 76829 3424
rect 70819 3380 70877 3381
rect 78604 3380 78644 3424
rect 80131 3423 80189 3424
rect 89251 3423 89309 3424
rect 85699 3380 85757 3381
rect 86083 3380 86141 3381
rect 92044 3380 92084 3424
rect 94723 3423 94781 3424
rect 95107 3423 95165 3424
rect 95491 3423 95549 3424
rect 95875 3423 95933 3424
rect 96643 3423 96701 3424
rect 97411 3423 97469 3424
rect 97795 3423 97853 3424
rect 97987 3464 98045 3465
rect 97987 3424 97996 3464
rect 98036 3424 98572 3464
rect 98612 3424 98621 3464
rect 97987 3423 98045 3424
rect 53635 3340 53644 3380
rect 53684 3340 55468 3380
rect 55508 3340 55517 3380
rect 57187 3340 57196 3380
rect 57236 3340 61760 3380
rect 62563 3340 62572 3380
rect 62612 3340 62621 3380
rect 62755 3340 62764 3380
rect 62804 3340 66452 3380
rect 66499 3340 66508 3380
rect 66548 3340 66700 3380
rect 66740 3340 66749 3380
rect 67075 3340 67084 3380
rect 67124 3340 70828 3380
rect 70868 3340 70877 3380
rect 71875 3340 71884 3380
rect 71924 3340 72500 3380
rect 72547 3340 72556 3380
rect 72596 3340 78644 3380
rect 79171 3340 79180 3380
rect 79220 3340 79229 3380
rect 79660 3340 79756 3380
rect 79796 3340 79805 3380
rect 85123 3340 85132 3380
rect 85172 3340 85420 3380
rect 85460 3340 85469 3380
rect 85614 3340 85708 3380
rect 85748 3340 85757 3380
rect 85998 3340 86092 3380
rect 86132 3340 86141 3380
rect 86851 3340 86860 3380
rect 86900 3340 92084 3380
rect 93667 3340 93676 3380
rect 93716 3340 94156 3380
rect 94196 3340 94205 3380
rect 97315 3340 97324 3380
rect 97364 3340 97996 3380
rect 98036 3340 98045 3380
rect 49219 3296 49277 3297
rect 49603 3296 49661 3297
rect 62572 3296 62612 3340
rect 63139 3296 63197 3297
rect 63811 3296 63869 3297
rect 66412 3296 66452 3340
rect 70819 3339 70877 3340
rect 68227 3296 68285 3297
rect 70627 3296 70685 3297
rect 72460 3296 72500 3340
rect 72739 3296 72797 3297
rect 75811 3296 75869 3297
rect 79180 3296 79220 3340
rect 37795 3256 37804 3296
rect 37844 3256 39532 3296
rect 39572 3256 39581 3296
rect 39715 3256 39724 3296
rect 39764 3256 40684 3296
rect 40724 3256 40733 3296
rect 40780 3256 44756 3296
rect 46600 3256 46636 3296
rect 46676 3256 46685 3296
rect 49134 3256 49228 3296
rect 49268 3256 49277 3296
rect 49518 3256 49612 3296
rect 49652 3256 49661 3296
rect 54787 3256 54796 3296
rect 54836 3256 54988 3296
rect 55028 3256 55037 3296
rect 55267 3256 55276 3296
rect 55316 3256 62612 3296
rect 63054 3256 63148 3296
rect 63188 3256 63197 3296
rect 63523 3256 63532 3296
rect 63572 3256 63820 3296
rect 63860 3256 63869 3296
rect 37795 3255 37853 3256
rect 39715 3255 39773 3256
rect 37507 3172 37516 3212
rect 37556 3172 39916 3212
rect 39956 3172 39965 3212
rect 34723 3088 34732 3128
rect 34772 3088 36884 3128
rect 36931 3088 36940 3128
rect 36980 3088 36989 3128
rect 37324 3088 39148 3128
rect 39188 3088 39197 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 6211 2920 6220 2960
rect 6260 2920 7372 2960
rect 7412 2920 7421 2960
rect 8332 2792 8372 3088
rect 20899 3087 20957 3088
rect 34723 3087 34781 3088
rect 19651 3044 19709 3045
rect 36844 3044 36884 3088
rect 40780 3044 40820 3256
rect 41539 3212 41597 3213
rect 46600 3212 46640 3256
rect 49219 3255 49277 3256
rect 49603 3255 49661 3256
rect 63139 3255 63197 3256
rect 63811 3255 63869 3256
rect 64240 3256 64780 3296
rect 64820 3256 64829 3296
rect 66412 3256 68236 3296
rect 68276 3256 68285 3296
rect 70541 3256 70550 3296
rect 70590 3256 70636 3296
rect 70676 3256 70685 3296
rect 71299 3256 71308 3296
rect 71348 3256 71788 3296
rect 71828 3256 71837 3296
rect 72451 3256 72460 3296
rect 72500 3256 72509 3296
rect 72739 3256 72748 3296
rect 72788 3256 72844 3296
rect 72884 3256 72893 3296
rect 73123 3256 73132 3296
rect 73172 3256 75820 3296
rect 75860 3256 75869 3296
rect 76963 3256 76972 3296
rect 77012 3256 79220 3296
rect 59491 3212 59549 3213
rect 60547 3212 60605 3213
rect 41539 3172 41548 3212
rect 41588 3172 46640 3212
rect 48931 3172 48940 3212
rect 48980 3172 50188 3212
rect 50228 3172 50237 3212
rect 53443 3172 53452 3212
rect 53492 3172 55852 3212
rect 55892 3172 55901 3212
rect 56803 3172 56812 3212
rect 56852 3172 57100 3212
rect 57140 3172 57149 3212
rect 59406 3172 59500 3212
rect 59540 3172 59549 3212
rect 59683 3172 59692 3212
rect 59732 3172 60268 3212
rect 60308 3172 60556 3212
rect 60596 3172 60605 3212
rect 60739 3172 60748 3212
rect 60788 3172 63436 3212
rect 63476 3172 63485 3212
rect 41539 3171 41597 3172
rect 59491 3171 59549 3172
rect 60547 3171 60605 3172
rect 55267 3128 55325 3129
rect 41539 3088 41548 3128
rect 41588 3088 44236 3128
rect 44276 3088 44285 3128
rect 48739 3088 48748 3128
rect 48788 3088 55276 3128
rect 55316 3088 55325 3128
rect 58915 3088 58924 3128
rect 58964 3088 61652 3128
rect 61795 3088 61804 3128
rect 61844 3088 61996 3128
rect 62036 3088 62045 3128
rect 62179 3088 62188 3128
rect 62228 3088 63916 3128
rect 63956 3088 63965 3128
rect 55267 3087 55325 3088
rect 54115 3044 54173 3045
rect 61612 3044 61652 3088
rect 63139 3044 63197 3045
rect 64240 3044 64280 3256
rect 68227 3255 68285 3256
rect 70627 3255 70685 3256
rect 72739 3255 72797 3256
rect 75811 3255 75869 3256
rect 78787 3212 78845 3213
rect 79660 3212 79700 3340
rect 85699 3339 85757 3340
rect 86083 3339 86141 3340
rect 81667 3256 81676 3296
rect 81716 3256 89300 3296
rect 87043 3212 87101 3213
rect 89260 3212 89300 3256
rect 90700 3256 94348 3296
rect 94388 3256 94397 3296
rect 90700 3212 90740 3256
rect 64387 3172 64396 3212
rect 64436 3172 64588 3212
rect 64628 3172 64637 3212
rect 65731 3172 65740 3212
rect 65780 3172 66028 3212
rect 66068 3172 66077 3212
rect 66307 3172 66316 3212
rect 66356 3172 68428 3212
rect 68468 3172 68477 3212
rect 71203 3172 71212 3212
rect 71252 3172 73420 3212
rect 73460 3172 73469 3212
rect 75331 3172 75340 3212
rect 75380 3172 75389 3212
rect 78787 3172 78796 3212
rect 78836 3172 79700 3212
rect 81091 3172 81100 3212
rect 81140 3172 84172 3212
rect 84212 3172 84221 3212
rect 86958 3172 87052 3212
rect 87092 3172 87101 3212
rect 87427 3172 87436 3212
rect 87476 3172 89164 3212
rect 89204 3172 89213 3212
rect 89260 3172 90740 3212
rect 93187 3172 93196 3212
rect 93236 3172 94540 3212
rect 94580 3172 94589 3212
rect 97027 3172 97036 3212
rect 97076 3172 98380 3212
rect 98420 3172 98429 3212
rect 75340 3128 75380 3172
rect 78787 3171 78845 3172
rect 87043 3171 87101 3172
rect 81667 3128 81725 3129
rect 72739 3088 72748 3128
rect 72788 3088 75380 3128
rect 77731 3088 77740 3128
rect 77780 3088 81044 3128
rect 8419 3004 8428 3044
rect 8468 3004 13364 3044
rect 13507 3004 13516 3044
rect 13556 3004 19660 3044
rect 19700 3004 19709 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 36844 3004 37516 3044
rect 37556 3004 37565 3044
rect 37780 3004 38284 3044
rect 38324 3004 40820 3044
rect 43171 3004 43180 3044
rect 43220 3004 46348 3044
rect 46388 3004 46397 3044
rect 46627 3004 46636 3044
rect 46676 3004 47404 3044
rect 47444 3004 47453 3044
rect 48643 3004 48652 3044
rect 48692 3004 49228 3044
rect 49268 3004 49277 3044
rect 50279 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50665 3044
rect 54115 3004 54124 3044
rect 54164 3004 61516 3044
rect 61556 3004 61565 3044
rect 61612 3004 63148 3044
rect 63188 3004 63197 3044
rect 13324 2960 13364 3004
rect 19651 3003 19709 3004
rect 17155 2960 17213 2961
rect 37780 2960 37820 3004
rect 54115 3003 54173 3004
rect 63139 3003 63197 3004
rect 63724 3004 64280 3044
rect 65399 3004 65408 3044
rect 65448 3004 65490 3044
rect 65530 3004 65572 3044
rect 65612 3004 65654 3044
rect 65694 3004 65736 3044
rect 65776 3004 65785 3044
rect 74371 3004 74380 3044
rect 74420 3004 75244 3044
rect 75284 3004 75293 3044
rect 75907 3004 75916 3044
rect 75956 3004 80468 3044
rect 80519 3004 80528 3044
rect 80568 3004 80610 3044
rect 80650 3004 80692 3044
rect 80732 3004 80774 3044
rect 80814 3004 80856 3044
rect 80896 3004 80905 3044
rect 54883 2960 54941 2961
rect 13324 2920 17164 2960
rect 17204 2920 17213 2960
rect 32131 2920 32140 2960
rect 32180 2920 34636 2960
rect 34676 2920 34685 2960
rect 35779 2920 35788 2960
rect 35828 2920 37820 2960
rect 38467 2920 38476 2960
rect 38516 2920 42892 2960
rect 42932 2920 42941 2960
rect 43075 2920 43084 2960
rect 43124 2920 43468 2960
rect 43508 2920 43517 2960
rect 43939 2920 43948 2960
rect 43988 2920 46924 2960
rect 46964 2920 46973 2960
rect 47491 2920 47500 2960
rect 47540 2920 51092 2960
rect 17155 2919 17213 2920
rect 19459 2876 19517 2877
rect 33667 2876 33725 2877
rect 34531 2876 34589 2877
rect 38476 2876 38516 2920
rect 41539 2876 41597 2877
rect 51052 2876 51092 2920
rect 54883 2920 54892 2960
rect 54932 2920 62284 2960
rect 62324 2920 62333 2960
rect 54883 2919 54941 2920
rect 57187 2876 57245 2877
rect 61891 2876 61949 2877
rect 13891 2836 13900 2876
rect 13940 2836 19468 2876
rect 19508 2836 19517 2876
rect 30595 2836 30604 2876
rect 30644 2836 32044 2876
rect 32084 2836 32093 2876
rect 33667 2836 33676 2876
rect 33716 2836 33868 2876
rect 33908 2836 33917 2876
rect 34531 2836 34540 2876
rect 34580 2836 38516 2876
rect 39043 2836 39052 2876
rect 39092 2836 41548 2876
rect 41588 2836 41597 2876
rect 43555 2836 43564 2876
rect 43604 2836 46540 2876
rect 46580 2836 46589 2876
rect 50467 2836 50476 2876
rect 50516 2836 50956 2876
rect 50996 2836 51005 2876
rect 51052 2836 55276 2876
rect 55316 2836 55325 2876
rect 57187 2836 57196 2876
rect 57236 2836 61228 2876
rect 61268 2836 61277 2876
rect 61806 2836 61900 2876
rect 61940 2836 61949 2876
rect 19459 2835 19517 2836
rect 33667 2835 33725 2836
rect 34531 2835 34589 2836
rect 41539 2835 41597 2836
rect 57187 2835 57245 2836
rect 61891 2835 61949 2836
rect 19363 2792 19421 2793
rect 46627 2792 46685 2793
rect 8332 2752 19372 2792
rect 19412 2752 19421 2792
rect 29059 2752 29068 2792
rect 29108 2752 31276 2792
rect 31316 2752 31325 2792
rect 31747 2752 31756 2792
rect 31796 2752 34060 2792
rect 34100 2752 34109 2792
rect 39235 2752 39244 2792
rect 39284 2752 43508 2792
rect 44323 2752 44332 2792
rect 44372 2752 46636 2792
rect 46676 2752 46685 2792
rect 19363 2751 19421 2752
rect 16579 2708 16637 2709
rect 38851 2708 38909 2709
rect 43468 2708 43508 2752
rect 46627 2751 46685 2752
rect 46819 2792 46877 2793
rect 60355 2792 60413 2793
rect 63724 2792 63764 3004
rect 73795 2960 73853 2961
rect 63907 2920 63916 2960
rect 63956 2920 64300 2960
rect 64340 2920 64349 2960
rect 64963 2920 64972 2960
rect 65012 2920 67276 2960
rect 67316 2920 67325 2960
rect 68227 2920 68236 2960
rect 68276 2920 73804 2960
rect 73844 2920 73853 2960
rect 74755 2920 74764 2960
rect 74804 2920 78028 2960
rect 78068 2920 78077 2960
rect 73795 2919 73853 2920
rect 80428 2876 80468 3004
rect 81004 2960 81044 3088
rect 81667 3088 81676 3128
rect 81716 3088 88724 3128
rect 81667 3087 81725 3088
rect 81283 3044 81341 3045
rect 81283 3004 81292 3044
rect 81332 3004 88588 3044
rect 88628 3004 88637 3044
rect 81283 3003 81341 3004
rect 88684 2960 88724 3088
rect 89356 3088 92812 3128
rect 92852 3088 92861 3128
rect 89356 2960 89396 3088
rect 95639 3004 95648 3044
rect 95688 3004 95730 3044
rect 95770 3004 95812 3044
rect 95852 3004 95894 3044
rect 95934 3004 95976 3044
rect 96016 3004 96025 3044
rect 98083 3004 98092 3044
rect 98132 3004 98380 3044
rect 98420 3004 98429 3044
rect 81004 2920 86668 2960
rect 86708 2920 86717 2960
rect 88684 2920 89396 2960
rect 90700 2920 96940 2960
rect 96980 2920 96989 2960
rect 81859 2876 81917 2877
rect 90700 2876 90740 2920
rect 64579 2836 64588 2876
rect 64628 2836 66796 2876
rect 66836 2836 66845 2876
rect 66979 2836 66988 2876
rect 67028 2836 69580 2876
rect 69620 2836 69629 2876
rect 76483 2836 76492 2876
rect 76532 2836 79564 2876
rect 79604 2836 79613 2876
rect 80428 2836 81812 2876
rect 81772 2792 81812 2836
rect 81859 2836 81868 2876
rect 81908 2836 90740 2876
rect 95683 2836 95692 2876
rect 95732 2836 96364 2876
rect 96404 2836 96413 2876
rect 81859 2835 81917 2836
rect 46819 2752 46828 2792
rect 46868 2752 47116 2792
rect 47156 2752 47165 2792
rect 48355 2752 48364 2792
rect 48404 2752 54604 2792
rect 54644 2752 54653 2792
rect 57091 2752 57100 2792
rect 57140 2752 57868 2792
rect 57908 2752 57917 2792
rect 60355 2752 60364 2792
rect 60404 2752 63764 2792
rect 63811 2752 63820 2792
rect 63860 2752 66124 2792
rect 66164 2752 66173 2792
rect 66499 2752 66508 2792
rect 66548 2752 68812 2792
rect 68852 2752 68861 2792
rect 75139 2752 75148 2792
rect 75188 2752 78412 2792
rect 78452 2752 78461 2792
rect 78883 2752 78892 2792
rect 78932 2752 81716 2792
rect 81772 2752 91276 2792
rect 91316 2752 91325 2792
rect 46819 2751 46877 2752
rect 60355 2751 60413 2752
rect 81676 2708 81716 2752
rect 16494 2668 16588 2708
rect 16628 2668 16637 2708
rect 27043 2668 27052 2708
rect 27092 2668 28492 2708
rect 28532 2668 28541 2708
rect 28675 2668 28684 2708
rect 28724 2668 31180 2708
rect 31220 2668 31229 2708
rect 32515 2668 32524 2708
rect 32564 2668 35212 2708
rect 35252 2668 35261 2708
rect 38851 2668 38860 2708
rect 38900 2668 41548 2708
rect 41588 2668 41597 2708
rect 41731 2668 41740 2708
rect 41780 2668 41789 2708
rect 42211 2668 42220 2708
rect 42260 2668 42508 2708
rect 42548 2668 42557 2708
rect 43468 2668 45292 2708
rect 45332 2668 45341 2708
rect 45859 2668 45868 2708
rect 45908 2668 48748 2708
rect 48788 2668 48797 2708
rect 57667 2668 57676 2708
rect 57716 2668 58828 2708
rect 58868 2668 58877 2708
rect 59971 2668 59980 2708
rect 60020 2668 63916 2708
rect 63956 2668 63965 2708
rect 65923 2668 65932 2708
rect 65972 2668 68044 2708
rect 68084 2668 68093 2708
rect 72067 2668 72076 2708
rect 72116 2668 74956 2708
rect 74996 2668 75005 2708
rect 81676 2668 82252 2708
rect 82292 2668 82301 2708
rect 87715 2668 87724 2708
rect 87764 2668 88108 2708
rect 88148 2668 88157 2708
rect 88579 2668 88588 2708
rect 88628 2668 96268 2708
rect 96308 2668 96317 2708
rect 16579 2667 16637 2668
rect 38851 2667 38909 2668
rect 16675 2624 16733 2625
rect 41740 2624 41780 2668
rect 75907 2624 75965 2625
rect 85987 2624 86045 2625
rect 8323 2584 8332 2624
rect 8372 2584 9524 2624
rect 15523 2584 15532 2624
rect 15572 2584 16532 2624
rect 16590 2584 16684 2624
rect 16724 2584 16733 2624
rect 9484 2540 9524 2584
rect 16492 2540 16532 2584
rect 16675 2583 16733 2584
rect 17452 2584 17548 2624
rect 17588 2584 17597 2624
rect 41740 2584 43852 2624
rect 43892 2584 43901 2624
rect 44707 2584 44716 2624
rect 44756 2584 46636 2624
rect 46676 2584 46685 2624
rect 46732 2584 48268 2624
rect 48308 2584 48317 2624
rect 58828 2584 59500 2624
rect 59540 2584 59549 2624
rect 65347 2584 65356 2624
rect 65396 2584 67660 2624
rect 67700 2584 67709 2624
rect 68803 2584 68812 2624
rect 68852 2584 71116 2624
rect 71156 2584 71165 2624
rect 71587 2584 71596 2624
rect 71636 2584 74188 2624
rect 74228 2584 74237 2624
rect 74956 2584 75916 2624
rect 75956 2584 75965 2624
rect 85902 2584 85996 2624
rect 86036 2584 86045 2624
rect 86659 2584 86668 2624
rect 86708 2584 90892 2624
rect 90932 2584 90941 2624
rect 96652 2584 97996 2624
rect 98036 2584 98045 2624
rect 1603 2500 1612 2540
rect 1652 2500 1661 2540
rect 1795 2500 1804 2540
rect 1844 2500 2956 2540
rect 2996 2500 3005 2540
rect 9475 2500 9484 2540
rect 9524 2500 9533 2540
rect 13572 2500 13612 2540
rect 13652 2500 13661 2540
rect 16492 2500 16724 2540
rect 1612 2372 1652 2500
rect 13612 2456 13652 2500
rect 15619 2456 15677 2457
rect 16684 2456 16724 2500
rect 17452 2456 17492 2584
rect 21379 2540 21437 2541
rect 46732 2540 46772 2584
rect 58828 2540 58868 2584
rect 74956 2540 74996 2584
rect 75907 2583 75965 2584
rect 85987 2583 86045 2584
rect 76099 2540 76157 2541
rect 87619 2540 87677 2541
rect 96652 2540 96692 2584
rect 21379 2500 21388 2540
rect 21428 2500 21484 2540
rect 21524 2500 21533 2540
rect 23652 2500 23692 2540
rect 23732 2500 23741 2540
rect 25572 2500 25612 2540
rect 25652 2500 25661 2540
rect 41155 2500 41164 2540
rect 41204 2500 41740 2540
rect 41780 2500 41789 2540
rect 41923 2500 41932 2540
rect 41972 2500 42892 2540
rect 42932 2500 42941 2540
rect 45475 2500 45484 2540
rect 45524 2500 46772 2540
rect 58819 2500 58828 2540
rect 58868 2500 58877 2540
rect 59971 2500 59980 2540
rect 60020 2500 60364 2540
rect 60404 2500 60413 2540
rect 74947 2500 74956 2540
rect 74996 2500 75005 2540
rect 76014 2500 76108 2540
rect 76148 2500 76157 2540
rect 85891 2500 85900 2540
rect 85940 2500 86036 2540
rect 86563 2500 86572 2540
rect 86612 2500 86956 2540
rect 86996 2500 87005 2540
rect 87534 2500 87628 2540
rect 87668 2500 87677 2540
rect 89316 2500 89356 2540
rect 89396 2500 89405 2540
rect 96643 2500 96652 2540
rect 96692 2500 96701 2540
rect 21379 2499 21437 2500
rect 23692 2456 23732 2500
rect 25612 2456 25652 2500
rect 76099 2499 76157 2500
rect 85891 2456 85949 2457
rect 5443 2416 5452 2456
rect 5492 2416 11360 2456
rect 13612 2416 14284 2456
rect 14324 2416 14333 2456
rect 15619 2416 15628 2456
rect 15668 2416 16396 2456
rect 16436 2416 16445 2456
rect 16684 2416 16972 2456
rect 17012 2416 17021 2456
rect 17452 2416 20044 2456
rect 20084 2416 20093 2456
rect 23692 2416 25228 2456
rect 25268 2416 25277 2456
rect 25612 2416 27532 2456
rect 27572 2416 27581 2456
rect 37219 2416 37228 2456
rect 37268 2416 44908 2456
rect 44948 2416 44957 2456
rect 45571 2416 45580 2456
rect 45620 2416 60692 2456
rect 61123 2416 61132 2456
rect 61172 2416 62668 2456
rect 62708 2416 62717 2456
rect 75523 2416 75532 2456
rect 75572 2416 76588 2456
rect 76628 2416 76637 2456
rect 76771 2416 76780 2456
rect 76820 2416 81332 2456
rect 84931 2416 84940 2456
rect 84980 2416 85900 2456
rect 85940 2416 85949 2456
rect 85996 2456 86036 2500
rect 87619 2499 87677 2500
rect 86179 2456 86237 2457
rect 89356 2456 89396 2500
rect 85996 2416 86188 2456
rect 86228 2416 86237 2456
rect 88867 2416 88876 2456
rect 88916 2416 89396 2456
rect 11320 2372 11360 2416
rect 15619 2415 15677 2416
rect 60652 2372 60692 2416
rect 62083 2372 62141 2373
rect 1612 2332 2572 2372
rect 2612 2332 2621 2372
rect 5827 2332 5836 2372
rect 5876 2332 6320 2372
rect 7939 2332 7948 2372
rect 7988 2332 9100 2372
rect 9140 2332 9149 2372
rect 11320 2332 29000 2372
rect 33955 2332 33964 2372
rect 34004 2332 34444 2372
rect 34484 2332 34493 2372
rect 38083 2332 38092 2372
rect 38132 2332 38476 2372
rect 38516 2332 38525 2372
rect 40771 2332 40780 2372
rect 40820 2332 41164 2372
rect 41204 2332 41213 2372
rect 54595 2332 54604 2372
rect 54644 2332 55756 2372
rect 55796 2332 55805 2372
rect 59011 2332 59020 2372
rect 59060 2332 60460 2372
rect 60500 2332 60509 2372
rect 60652 2332 62092 2372
rect 62132 2332 62141 2372
rect 62275 2332 62284 2372
rect 62324 2332 63340 2372
rect 63380 2332 63389 2372
rect 69763 2332 69772 2372
rect 69812 2332 70444 2372
rect 70484 2332 70493 2372
rect 76675 2332 76684 2372
rect 76724 2332 78028 2372
rect 78068 2332 78077 2372
rect 78211 2332 78220 2372
rect 78260 2332 79660 2372
rect 79700 2332 79709 2372
rect 6280 2288 6320 2332
rect 16579 2288 16637 2289
rect 28960 2288 29000 2332
rect 62083 2331 62141 2332
rect 56611 2288 56669 2289
rect 81292 2288 81332 2416
rect 85891 2415 85949 2416
rect 86179 2415 86237 2416
rect 87619 2372 87677 2373
rect 82051 2332 82060 2372
rect 82100 2332 85324 2372
rect 85364 2332 85373 2372
rect 85891 2332 85900 2372
rect 85940 2332 87628 2372
rect 87668 2332 87677 2372
rect 89347 2332 89356 2372
rect 89396 2332 90700 2372
rect 90740 2332 90749 2372
rect 97987 2332 97996 2372
rect 98036 2332 98476 2372
rect 98516 2332 98525 2372
rect 87619 2331 87677 2332
rect 6280 2248 11360 2288
rect 12163 2248 12172 2288
rect 12212 2248 13324 2288
rect 13364 2248 13373 2288
rect 16579 2248 16588 2288
rect 16628 2248 25132 2288
rect 25172 2248 25181 2288
rect 28960 2248 30892 2288
rect 30932 2248 30941 2288
rect 34339 2248 34348 2288
rect 34388 2248 35020 2288
rect 35060 2248 35069 2288
rect 55363 2248 55372 2288
rect 55412 2248 56620 2288
rect 56660 2248 56669 2288
rect 58051 2248 58060 2288
rect 58100 2248 59308 2288
rect 59348 2248 59357 2288
rect 75907 2248 75916 2288
rect 75956 2248 77164 2288
rect 77204 2248 77213 2288
rect 78403 2248 78412 2288
rect 78452 2248 80428 2288
rect 80468 2248 80477 2288
rect 81292 2248 90508 2288
rect 90548 2248 90557 2288
rect 11320 2204 11360 2248
rect 16579 2247 16637 2248
rect 56611 2247 56669 2248
rect 71203 2204 71261 2205
rect 7171 2164 7180 2204
rect 7220 2164 8332 2204
rect 8372 2164 8381 2204
rect 8707 2164 8716 2204
rect 8756 2164 9676 2204
rect 9716 2164 9725 2204
rect 11320 2164 21964 2204
rect 22004 2164 22013 2204
rect 57283 2164 57292 2204
rect 57332 2164 58156 2204
rect 58196 2164 58205 2204
rect 58435 2164 58444 2204
rect 58484 2164 59116 2204
rect 59156 2164 59165 2204
rect 61603 2164 61612 2204
rect 61652 2164 64396 2204
rect 64436 2164 64445 2204
rect 71203 2164 71212 2204
rect 71252 2164 75284 2204
rect 78595 2164 78604 2204
rect 78644 2164 80236 2204
rect 80276 2164 80285 2204
rect 80332 2164 83692 2204
rect 83732 2164 83741 2204
rect 71203 2163 71261 2164
rect 21379 2120 21437 2121
rect 75244 2120 75284 2164
rect 80332 2120 80372 2164
rect 2371 2080 2380 2120
rect 2420 2080 3340 2120
rect 3380 2080 3389 2120
rect 7363 2080 7372 2120
rect 7412 2080 21388 2120
rect 21428 2080 21437 2120
rect 37123 2080 37132 2120
rect 37172 2080 38284 2120
rect 38324 2080 38333 2120
rect 72451 2080 72460 2120
rect 72500 2080 74284 2120
rect 74324 2080 74333 2120
rect 75244 2080 80372 2120
rect 80995 2080 81004 2120
rect 81044 2080 90124 2120
rect 90164 2080 90173 2120
rect 21379 2079 21437 2080
rect 1699 1996 1708 2036
rect 1748 1996 1996 2036
rect 2036 1996 2045 2036
rect 5731 1996 5740 2036
rect 5780 1996 6412 2036
rect 6452 1996 6461 2036
rect 6787 1996 6796 2036
rect 6836 1996 7948 2036
rect 7988 1996 7997 2036
rect 10540 1996 22252 2036
rect 22292 1996 22301 2036
rect 31651 1996 31660 2036
rect 31700 1996 32332 2036
rect 32372 1996 32381 2036
rect 33187 1996 33196 2036
rect 33236 1996 34828 2036
rect 34868 1996 34877 2036
rect 36739 1996 36748 2036
rect 36788 1996 37708 2036
rect 37748 1996 37757 2036
rect 41347 1996 41356 2036
rect 41396 1996 42700 2036
rect 42740 1996 42749 2036
rect 50563 1996 50572 2036
rect 50612 1996 50860 2036
rect 50900 1996 50909 2036
rect 59395 1996 59404 2036
rect 59444 1996 61420 2036
rect 61460 1996 61469 2036
rect 70915 1996 70924 2036
rect 70964 1996 72556 2036
rect 72596 1996 72605 2036
rect 75619 1996 75628 2036
rect 75668 1996 81196 2036
rect 81236 1996 81245 2036
rect 83299 1996 83308 2036
rect 83348 1996 85516 2036
rect 85556 1996 85565 2036
rect 96931 1996 96940 2036
rect 96980 1996 97708 2036
rect 97748 1996 97757 2036
rect 2083 1912 2092 1952
rect 2132 1912 2380 1952
rect 2420 1912 2429 1952
rect 5539 1912 5548 1952
rect 5588 1912 5836 1952
rect 5876 1912 5885 1952
rect 6019 1912 6028 1952
rect 6068 1912 7180 1952
rect 7220 1912 7229 1952
rect 5635 1828 5644 1868
rect 5684 1828 6796 1868
rect 6836 1828 6845 1868
rect 10540 1784 10580 1996
rect 16675 1952 16733 1953
rect 86179 1952 86237 1953
rect 11779 1912 11788 1952
rect 11828 1912 12940 1952
rect 12980 1912 12989 1952
rect 16675 1912 16684 1952
rect 16724 1912 18604 1952
rect 18644 1912 18653 1952
rect 81283 1912 81292 1952
rect 81332 1912 86188 1952
rect 86228 1912 86237 1952
rect 88579 1912 88588 1952
rect 88628 1912 89932 1952
rect 89972 1912 89981 1952
rect 16675 1911 16733 1912
rect 86179 1911 86237 1912
rect 11011 1828 11020 1868
rect 11060 1828 12172 1868
rect 12212 1828 12221 1868
rect 20611 1828 20620 1868
rect 20660 1828 23020 1868
rect 23060 1828 23069 1868
rect 26371 1828 26380 1868
rect 26420 1828 28684 1868
rect 28724 1828 28733 1868
rect 60355 1828 60364 1868
rect 60404 1828 63244 1868
rect 63284 1828 63293 1868
rect 68227 1828 68236 1868
rect 68276 1828 69676 1868
rect 69716 1828 69725 1868
rect 73315 1828 73324 1868
rect 73364 1828 81332 1868
rect 4675 1744 4684 1784
rect 4724 1744 6028 1784
rect 6068 1744 6077 1784
rect 6691 1744 6700 1784
rect 6740 1744 10580 1784
rect 10627 1744 10636 1784
rect 10676 1744 11788 1784
rect 11828 1744 11837 1784
rect 22915 1744 22924 1784
rect 22964 1744 24748 1784
rect 24788 1744 24797 1784
rect 25987 1744 25996 1784
rect 26036 1744 28108 1784
rect 28148 1744 28157 1784
rect 29443 1744 29452 1784
rect 29492 1744 30220 1784
rect 30260 1744 30269 1784
rect 32803 1744 32812 1784
rect 32852 1744 34252 1784
rect 34292 1744 34301 1784
rect 38179 1744 38188 1784
rect 38228 1744 40012 1784
rect 40052 1744 40061 1784
rect 52483 1744 52492 1784
rect 52532 1744 54124 1784
rect 54164 1744 54173 1784
rect 56707 1744 56716 1784
rect 56756 1744 60556 1784
rect 60596 1744 60605 1784
rect 72835 1744 72844 1784
rect 72884 1744 75724 1784
rect 75764 1744 75773 1784
rect 4483 1660 4492 1700
rect 4532 1660 5644 1700
rect 5684 1660 5693 1700
rect 6307 1660 6316 1700
rect 6356 1660 7564 1700
rect 7604 1660 7613 1700
rect 9859 1660 9868 1700
rect 9908 1660 11020 1700
rect 11060 1660 11069 1700
rect 11395 1660 11404 1700
rect 11444 1660 12556 1700
rect 12596 1660 12605 1700
rect 12739 1660 12748 1700
rect 12788 1660 13132 1700
rect 13172 1660 13181 1700
rect 14467 1660 14476 1700
rect 14516 1660 16492 1700
rect 16532 1660 16541 1700
rect 21859 1660 21868 1700
rect 21908 1660 23692 1700
rect 23732 1660 23741 1700
rect 24835 1660 24844 1700
rect 24884 1660 26380 1700
rect 26420 1660 26429 1700
rect 35875 1660 35884 1700
rect 35924 1660 37516 1700
rect 37556 1660 37565 1700
rect 37987 1660 37996 1700
rect 38036 1660 39532 1700
rect 39572 1660 39581 1700
rect 40099 1660 40108 1700
rect 40148 1660 42508 1700
rect 42548 1660 42557 1700
rect 51907 1660 51916 1700
rect 51956 1660 53356 1700
rect 53396 1660 53405 1700
rect 55171 1660 55180 1700
rect 55220 1660 57964 1700
rect 58004 1660 58013 1700
rect 63235 1660 63244 1700
rect 63284 1660 66028 1700
rect 66068 1660 66077 1700
rect 71299 1660 71308 1700
rect 71348 1660 73804 1700
rect 73844 1660 73853 1700
rect 74179 1660 74188 1700
rect 74228 1660 77260 1700
rect 77300 1660 77309 1700
rect 81292 1616 81332 1828
rect 90700 1744 91084 1784
rect 91124 1744 91133 1784
rect 91267 1744 91276 1784
rect 91316 1744 92620 1784
rect 92660 1744 92669 1784
rect 92803 1744 92812 1784
rect 92852 1744 94156 1784
rect 94196 1744 94205 1784
rect 94723 1744 94732 1784
rect 94772 1744 96076 1784
rect 96116 1744 96125 1784
rect 90700 1700 90740 1744
rect 81859 1660 81868 1700
rect 81908 1660 82060 1700
rect 82100 1660 82109 1700
rect 82924 1660 88876 1700
rect 88916 1660 88925 1700
rect 89836 1660 90740 1700
rect 90883 1660 90892 1700
rect 90932 1660 92236 1700
rect 92276 1660 92285 1700
rect 92419 1660 92428 1700
rect 92468 1660 93772 1700
rect 93812 1660 93821 1700
rect 93955 1660 93964 1700
rect 94004 1660 95308 1700
rect 95348 1660 95357 1700
rect 95875 1660 95884 1700
rect 95924 1660 97228 1700
rect 97268 1660 97277 1700
rect 82924 1616 82964 1660
rect 89836 1616 89876 1660
rect 4099 1576 4108 1616
rect 4148 1576 5260 1616
rect 5300 1576 5309 1616
rect 9571 1576 9580 1616
rect 9620 1576 10636 1616
rect 10676 1576 10685 1616
rect 13411 1576 13420 1616
rect 13460 1576 15052 1616
rect 15092 1576 15101 1616
rect 15235 1576 15244 1616
rect 15284 1576 17740 1616
rect 17780 1576 17789 1616
rect 19075 1576 19084 1616
rect 19124 1576 21580 1616
rect 21620 1576 21629 1616
rect 23299 1576 23308 1616
rect 23348 1576 25036 1616
rect 25076 1576 25085 1616
rect 27427 1576 27436 1616
rect 27476 1576 29452 1616
rect 29492 1576 29501 1616
rect 30979 1576 30988 1616
rect 31028 1576 32716 1616
rect 32756 1576 32765 1616
rect 34531 1576 34540 1616
rect 34580 1576 36748 1616
rect 36788 1576 36797 1616
rect 37411 1576 37420 1616
rect 37460 1576 39244 1616
rect 39284 1576 39293 1616
rect 39715 1576 39724 1616
rect 39764 1576 41932 1616
rect 41972 1576 41981 1616
rect 42403 1576 42412 1616
rect 42452 1576 45580 1616
rect 45620 1576 45629 1616
rect 48163 1576 48172 1616
rect 48212 1576 49804 1616
rect 49844 1576 49853 1616
rect 51523 1576 51532 1616
rect 51572 1576 52012 1616
rect 52052 1576 52061 1616
rect 52291 1576 52300 1616
rect 52340 1576 53740 1616
rect 53780 1576 53789 1616
rect 54211 1576 54220 1616
rect 54260 1576 56620 1616
rect 56660 1576 56669 1616
rect 57475 1576 57484 1616
rect 57524 1576 60940 1616
rect 60980 1576 60989 1616
rect 64195 1576 64204 1616
rect 64244 1576 66412 1616
rect 66452 1576 66461 1616
rect 68035 1576 68044 1616
rect 68084 1576 70348 1616
rect 70388 1576 70397 1616
rect 70819 1576 70828 1616
rect 70868 1576 73036 1616
rect 73076 1576 73085 1616
rect 81292 1576 82964 1616
rect 83011 1576 83020 1616
rect 83060 1576 86860 1616
rect 86900 1576 86909 1616
rect 88003 1576 88012 1616
rect 88052 1576 89548 1616
rect 89588 1576 89597 1616
rect 89827 1576 89836 1616
rect 89876 1576 89885 1616
rect 90115 1576 90124 1616
rect 90164 1576 91468 1616
rect 91508 1576 91517 1616
rect 91651 1576 91660 1616
rect 91700 1576 93004 1616
rect 93044 1576 93053 1616
rect 93571 1576 93580 1616
rect 93620 1576 94924 1616
rect 94964 1576 94973 1616
rect 95107 1576 95116 1616
rect 95156 1576 96460 1616
rect 96500 1576 96509 1616
rect 3715 1492 3724 1532
rect 3764 1492 4876 1532
rect 4916 1492 4925 1532
rect 10243 1492 10252 1532
rect 10292 1492 11404 1532
rect 11444 1492 11453 1532
rect 13027 1492 13036 1532
rect 13076 1492 14476 1532
rect 14516 1492 14525 1532
rect 14851 1492 14860 1532
rect 14900 1492 17164 1532
rect 17204 1492 17213 1532
rect 19459 1492 19468 1532
rect 19508 1492 21964 1532
rect 22004 1492 22013 1532
rect 22147 1492 22156 1532
rect 22196 1492 23884 1532
rect 23924 1492 23933 1532
rect 24451 1492 24460 1532
rect 24500 1492 25804 1532
rect 25844 1492 25853 1532
rect 26851 1492 26860 1532
rect 26900 1492 28876 1532
rect 28916 1492 28925 1532
rect 38563 1492 38572 1532
rect 38612 1492 40204 1532
rect 40244 1492 40253 1532
rect 48547 1492 48556 1532
rect 48596 1492 49996 1532
rect 50036 1492 50045 1532
rect 54979 1492 54988 1532
rect 55028 1492 57580 1532
rect 57620 1492 57629 1532
rect 71683 1492 71692 1532
rect 71732 1492 74572 1532
rect 74612 1492 74621 1532
rect 81475 1492 81484 1532
rect 81524 1492 84556 1532
rect 84596 1492 84605 1532
rect 86083 1492 86092 1532
rect 86132 1492 88396 1532
rect 88436 1492 88445 1532
rect 88963 1492 88972 1532
rect 89012 1492 90316 1532
rect 90356 1492 90365 1532
rect 90499 1492 90508 1532
rect 90548 1492 91852 1532
rect 91892 1492 91901 1532
rect 92035 1492 92044 1532
rect 92084 1492 93388 1532
rect 93428 1492 93437 1532
rect 94339 1492 94348 1532
rect 94388 1492 95500 1532
rect 95540 1492 95549 1532
rect 96259 1492 96268 1532
rect 96308 1492 97612 1532
rect 97652 1492 97661 1532
rect 3139 1408 3148 1448
rect 3188 1408 32780 1448
rect 36643 1408 36652 1448
rect 36692 1408 38668 1448
rect 38708 1408 38717 1448
rect 40867 1408 40876 1448
rect 40916 1408 43660 1448
rect 43700 1408 43709 1448
rect 53059 1408 53068 1448
rect 53108 1408 55084 1448
rect 55124 1408 55133 1448
rect 57859 1408 57868 1448
rect 57908 1408 61324 1448
rect 61364 1408 61373 1448
rect 73795 1408 73804 1448
rect 73844 1408 76876 1448
rect 76916 1408 76925 1448
rect 80899 1408 80908 1448
rect 80948 1408 82348 1448
rect 82388 1408 82397 1448
rect 82627 1408 82636 1448
rect 82676 1408 86476 1448
rect 86516 1408 86525 1448
rect 87235 1408 87244 1448
rect 87284 1408 88492 1448
rect 88532 1408 88541 1448
rect 96451 1408 96460 1448
rect 96500 1408 97132 1448
rect 97172 1408 97181 1448
rect 32740 1364 32780 1408
rect 71779 1364 71837 1365
rect 9187 1324 9196 1364
rect 9236 1324 10252 1364
rect 10292 1324 10301 1364
rect 13987 1324 13996 1364
rect 14036 1324 14860 1364
rect 14900 1324 14909 1364
rect 15619 1324 15628 1364
rect 15668 1324 18220 1364
rect 18260 1324 18269 1364
rect 19843 1324 19852 1364
rect 19892 1324 22348 1364
rect 22388 1324 22397 1364
rect 24067 1324 24076 1364
rect 24116 1324 25420 1364
rect 25460 1324 25469 1364
rect 27139 1324 27148 1364
rect 27188 1324 29068 1364
rect 29108 1324 29117 1364
rect 29923 1324 29932 1364
rect 29972 1324 31756 1364
rect 31796 1324 31805 1364
rect 32740 1324 34924 1364
rect 34964 1324 34973 1364
rect 53827 1324 53836 1364
rect 53876 1324 56236 1364
rect 56276 1324 56285 1364
rect 66883 1324 66892 1364
rect 66932 1324 69196 1364
rect 69236 1324 69245 1364
rect 71779 1324 71788 1364
rect 71828 1324 81292 1364
rect 81332 1324 81341 1364
rect 82243 1324 82252 1364
rect 82292 1324 86188 1364
rect 86228 1324 86237 1364
rect 86659 1324 86668 1364
rect 86708 1324 87916 1364
rect 87956 1324 87965 1364
rect 88387 1324 88396 1364
rect 88436 1324 89068 1364
rect 89108 1324 89117 1364
rect 90307 1324 90316 1364
rect 90356 1324 90988 1364
rect 91028 1324 91037 1364
rect 95491 1324 95500 1364
rect 95540 1324 96844 1364
rect 96884 1324 96893 1364
rect 97603 1324 97612 1364
rect 97652 1324 98764 1364
rect 98804 1324 98813 1364
rect 71779 1323 71837 1324
rect 79939 1280 79997 1281
rect 85795 1280 85853 1281
rect 3043 1240 3052 1280
rect 3092 1240 4108 1280
rect 4148 1240 4157 1280
rect 13219 1240 13228 1280
rect 13268 1240 13708 1280
rect 13748 1240 13757 1280
rect 14755 1240 14764 1280
rect 14804 1240 15436 1280
rect 15476 1240 15485 1280
rect 16291 1240 16300 1280
rect 16340 1240 18124 1280
rect 18164 1240 18173 1280
rect 18307 1240 18316 1280
rect 18356 1240 20236 1280
rect 20276 1240 20285 1280
rect 23491 1240 23500 1280
rect 23540 1240 24652 1280
rect 24692 1240 24701 1280
rect 25507 1240 25516 1280
rect 25556 1240 25996 1280
rect 26036 1240 26045 1280
rect 28579 1240 28588 1280
rect 28628 1240 29836 1280
rect 29876 1240 29885 1280
rect 30211 1240 30220 1280
rect 30260 1240 31564 1280
rect 31604 1240 31613 1280
rect 32419 1240 32428 1280
rect 32468 1240 33484 1280
rect 33524 1240 33533 1280
rect 34723 1240 34732 1280
rect 34772 1240 35788 1280
rect 35828 1240 35837 1280
rect 36355 1240 36364 1280
rect 36404 1240 37132 1280
rect 37172 1240 37181 1280
rect 39619 1240 39628 1280
rect 39668 1240 40780 1280
rect 40820 1240 40829 1280
rect 42787 1240 42796 1280
rect 42836 1240 45964 1280
rect 46004 1240 46013 1280
rect 47683 1240 47692 1280
rect 47732 1240 48076 1280
rect 48116 1240 48125 1280
rect 51715 1240 51724 1280
rect 51764 1240 52972 1280
rect 53012 1240 53021 1280
rect 53251 1240 53260 1280
rect 53300 1240 55468 1280
rect 55508 1240 55517 1280
rect 58627 1240 58636 1280
rect 58676 1240 61708 1280
rect 61748 1240 61757 1280
rect 64003 1240 64012 1280
rect 64052 1240 65068 1280
rect 65108 1240 65117 1280
rect 65923 1240 65932 1280
rect 65972 1240 67372 1280
rect 67412 1240 67421 1280
rect 69379 1240 69388 1280
rect 69428 1240 71884 1280
rect 71924 1240 71933 1280
rect 73219 1240 73228 1280
rect 73268 1240 76012 1280
rect 76052 1240 76061 1280
rect 77443 1240 77452 1280
rect 77492 1240 79756 1280
rect 79796 1240 79805 1280
rect 79854 1240 79948 1280
rect 79988 1240 79997 1280
rect 80515 1240 80524 1280
rect 80564 1240 82732 1280
rect 82772 1240 82781 1280
rect 83971 1240 83980 1280
rect 84020 1240 85228 1280
rect 85268 1240 85277 1280
rect 85507 1240 85516 1280
rect 85556 1240 85804 1280
rect 85844 1240 85853 1280
rect 87811 1240 87820 1280
rect 87860 1240 88684 1280
rect 88724 1240 88733 1280
rect 89155 1240 89164 1280
rect 89204 1240 89644 1280
rect 89684 1240 89693 1280
rect 89923 1240 89932 1280
rect 89972 1240 90412 1280
rect 90452 1240 90461 1280
rect 79939 1239 79997 1240
rect 85795 1239 85853 1240
rect 35683 1196 35741 1197
rect 85987 1196 86045 1197
rect 2851 1156 2860 1196
rect 2900 1156 3148 1196
rect 3188 1156 3197 1196
rect 3427 1156 3436 1196
rect 3476 1156 4492 1196
rect 4532 1156 4541 1196
rect 15331 1156 15340 1196
rect 15380 1156 16588 1196
rect 16628 1156 16637 1196
rect 16867 1156 16876 1196
rect 16916 1156 17356 1196
rect 17396 1156 17405 1196
rect 20899 1156 20908 1196
rect 20948 1156 22156 1196
rect 22196 1156 22205 1196
rect 23395 1156 23404 1196
rect 23444 1156 24076 1196
rect 24116 1156 24125 1196
rect 25891 1156 25900 1196
rect 25940 1156 26572 1196
rect 26612 1156 26621 1196
rect 28963 1156 28972 1196
rect 29012 1156 30412 1196
rect 30452 1156 30461 1196
rect 31363 1156 31372 1196
rect 31412 1156 33292 1196
rect 33332 1156 33341 1196
rect 35395 1156 35404 1196
rect 35444 1156 35692 1196
rect 35732 1156 35741 1196
rect 37027 1156 37036 1196
rect 37076 1156 39052 1196
rect 39092 1156 39101 1196
rect 40291 1156 40300 1196
rect 40340 1156 41548 1196
rect 41588 1156 41597 1196
rect 45091 1156 45100 1196
rect 45140 1156 47884 1196
rect 47924 1156 47933 1196
rect 59779 1156 59788 1196
rect 59828 1156 61996 1196
rect 62036 1156 62045 1196
rect 62659 1156 62668 1196
rect 62708 1156 64684 1196
rect 64724 1156 64733 1196
rect 68611 1156 68620 1196
rect 68660 1156 70732 1196
rect 70772 1156 70781 1196
rect 73027 1156 73036 1196
rect 73076 1156 75052 1196
rect 75092 1156 75101 1196
rect 76291 1156 76300 1196
rect 76340 1156 79180 1196
rect 79220 1156 79229 1196
rect 80131 1156 80140 1196
rect 80180 1156 83404 1196
rect 83444 1156 83453 1196
rect 84163 1156 84172 1196
rect 84212 1156 85996 1196
rect 86036 1156 86045 1196
rect 35683 1155 35741 1156
rect 85987 1155 86045 1156
rect 14371 1072 14380 1112
rect 14420 1072 16204 1112
rect 16244 1072 16253 1112
rect 18787 1072 18796 1112
rect 18836 1072 20620 1112
rect 20660 1072 20669 1112
rect 22531 1072 22540 1112
rect 22580 1072 24460 1112
rect 24500 1072 24509 1112
rect 30115 1072 30124 1112
rect 30164 1072 30988 1112
rect 31028 1072 31037 1112
rect 34147 1072 34156 1112
rect 34196 1072 36556 1112
rect 36596 1072 36605 1112
rect 38947 1072 38956 1112
rect 38996 1072 40588 1112
rect 40628 1072 40637 1112
rect 47203 1072 47212 1112
rect 47252 1072 47692 1112
rect 47732 1072 47741 1112
rect 56515 1072 56524 1112
rect 56564 1072 58924 1112
rect 58964 1072 58973 1112
rect 59203 1072 59212 1112
rect 59252 1072 62092 1112
rect 62132 1072 62141 1112
rect 67459 1072 67468 1112
rect 67508 1072 69964 1112
rect 70004 1072 70013 1112
rect 74563 1072 74572 1112
rect 74612 1072 77644 1112
rect 77684 1072 77693 1112
rect 79555 1072 79564 1112
rect 79604 1072 82924 1112
rect 82964 1072 82973 1112
rect 83203 1072 83212 1112
rect 83252 1072 84844 1112
rect 84884 1072 84893 1112
rect 86851 1072 86860 1112
rect 86900 1072 88780 1112
rect 88820 1072 88829 1112
rect 9379 988 9388 1028
rect 9428 988 9676 1028
rect 9716 988 9725 1028
rect 13795 988 13804 1028
rect 13844 988 15628 1028
rect 15668 988 15677 1028
rect 18691 988 18700 1028
rect 18740 988 21004 1028
rect 21044 988 21053 1028
rect 21475 988 21484 1028
rect 21524 988 23500 1028
rect 23540 988 23549 1028
rect 26275 988 26284 1028
rect 26324 988 27148 1028
rect 27188 988 27197 1028
rect 28387 988 28396 1028
rect 28436 988 30796 1028
rect 30836 988 30845 1028
rect 33763 988 33772 1028
rect 33812 988 36364 1028
rect 36404 988 36413 1028
rect 42019 988 42028 1028
rect 42068 988 45196 1028
rect 45236 988 45245 1028
rect 56131 988 56140 1028
rect 56180 988 58540 1028
rect 58580 988 58589 1028
rect 60931 988 60940 1028
rect 60980 988 63724 1028
rect 63764 988 63773 1028
rect 69187 988 69196 1028
rect 69236 988 71500 1028
rect 71540 988 71549 1028
rect 75715 988 75724 1028
rect 75764 988 76880 1028
rect 77059 988 77068 1028
rect 77108 988 79852 1028
rect 79892 988 79901 1028
rect 81283 988 81292 1028
rect 81332 988 83500 1028
rect 83540 988 83549 1028
rect 85315 988 85324 1028
rect 85364 988 88108 1028
rect 88148 988 88157 1028
rect 16675 904 16684 944
rect 16724 904 19084 944
rect 19124 904 19133 944
rect 20707 904 20716 944
rect 20756 904 22540 944
rect 22580 904 22589 944
rect 29731 904 29740 944
rect 29780 904 30604 944
rect 30644 904 30653 944
rect 32899 904 32908 944
rect 32948 904 32957 944
rect 33379 904 33388 944
rect 33428 904 36172 944
rect 36212 904 36221 944
rect 41635 904 41644 944
rect 41684 904 44812 944
rect 44852 904 44861 944
rect 61315 904 61324 944
rect 61364 904 64108 944
rect 64148 904 64157 944
rect 69955 904 69964 944
rect 70004 904 72268 944
rect 72308 904 72317 944
rect 73603 904 73612 944
rect 73652 904 76396 944
rect 76436 904 76445 944
rect 20707 860 20765 861
rect 32908 860 32948 904
rect 76840 860 76880 988
rect 77635 904 77644 944
rect 77684 904 80332 944
rect 80372 904 80381 944
rect 85699 860 85757 861
rect 17059 820 17068 860
rect 17108 820 17932 860
rect 17972 820 17981 860
rect 20707 820 20716 860
rect 20756 820 22924 860
rect 22964 820 22973 860
rect 32908 820 35980 860
rect 36020 820 36029 860
rect 60163 820 60172 860
rect 60212 820 62380 860
rect 62420 820 62429 860
rect 67651 820 67660 860
rect 67700 820 69292 860
rect 69332 820 69341 860
rect 73987 820 73996 860
rect 74036 820 76204 860
rect 76244 820 76253 860
rect 76840 820 78796 860
rect 78836 820 78845 860
rect 82435 820 82444 860
rect 82484 820 85708 860
rect 85748 820 85757 860
rect 20707 819 20765 820
rect 85699 819 85757 820
rect 13123 736 13132 776
rect 13172 736 22828 776
rect 22868 736 22877 776
rect 32227 736 32236 776
rect 32276 736 32908 776
rect 32948 736 32957 776
rect 40483 736 40492 776
rect 40532 736 43084 776
rect 43124 736 43133 776
rect 55747 736 55756 776
rect 55796 736 58732 776
rect 58772 736 58781 776
rect 77827 736 77836 776
rect 77876 736 80044 776
rect 80084 736 80093 776
rect 80323 736 80332 776
rect 80372 736 81964 776
rect 82004 736 82013 776
rect 83587 736 83596 776
rect 83636 736 86764 776
rect 86804 736 86813 776
rect 18019 652 18028 692
rect 18068 652 19852 692
rect 19892 652 19901 692
rect 79747 652 79756 692
rect 79796 652 82156 692
rect 82196 652 82205 692
rect 84547 652 84556 692
rect 84596 652 87532 692
rect 87572 652 87581 692
rect 12835 568 12844 608
rect 12884 568 13132 608
rect 13172 568 13181 608
rect 16771 568 16780 608
rect 16820 568 19468 608
rect 19508 568 19517 608
rect 39331 568 39340 608
rect 39380 568 41356 608
rect 41396 568 41405 608
rect 82051 568 82060 608
rect 82100 568 85612 608
rect 85652 568 85661 608
rect 12451 484 12460 524
rect 12500 484 13900 524
rect 13940 484 13949 524
rect 70339 484 70348 524
rect 70388 484 72652 524
rect 72692 484 72701 524
rect 83779 484 83788 524
rect 83828 484 87340 524
rect 87380 484 87389 524
rect 16483 400 16492 440
rect 16532 400 16780 440
rect 16820 400 16829 440
rect 80707 400 80716 440
rect 80756 400 83692 440
rect 83732 400 83741 440
rect 15907 316 15916 356
rect 15956 316 18892 356
rect 18932 316 18941 356
rect 41251 316 41260 356
rect 41300 316 44236 356
rect 44276 316 44285 356
rect 86083 272 86141 273
rect 42307 232 42316 272
rect 42356 232 45004 272
rect 45044 232 45053 272
rect 55555 232 55564 272
rect 55604 232 58348 272
rect 58388 232 58397 272
rect 82819 232 82828 272
rect 82868 232 86092 272
rect 86132 232 86141 272
rect 86083 231 86141 232
rect 79843 188 79901 189
rect 36259 148 36268 188
rect 36308 148 38132 188
rect 79363 148 79372 188
rect 79412 148 79852 188
rect 79892 148 79901 188
rect 38092 104 38132 148
rect 79843 147 79901 148
rect 88780 148 89260 188
rect 89300 148 89309 188
rect 88780 104 88820 148
rect 38083 64 38092 104
rect 38132 64 38141 104
rect 88771 64 88780 104
rect 88820 64 88829 104
<< via3 >>
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 33928 11320 33968 11360
rect 34010 11320 34050 11360
rect 34092 11320 34132 11360
rect 34174 11320 34214 11360
rect 34256 11320 34296 11360
rect 49048 11320 49088 11360
rect 49130 11320 49170 11360
rect 49212 11320 49252 11360
rect 49294 11320 49334 11360
rect 49376 11320 49416 11360
rect 64168 11320 64208 11360
rect 64250 11320 64290 11360
rect 64332 11320 64372 11360
rect 64414 11320 64454 11360
rect 64496 11320 64536 11360
rect 79288 11320 79328 11360
rect 79370 11320 79410 11360
rect 79452 11320 79492 11360
rect 79534 11320 79574 11360
rect 79616 11320 79656 11360
rect 94408 11320 94448 11360
rect 94490 11320 94530 11360
rect 94572 11320 94612 11360
rect 94654 11320 94694 11360
rect 94736 11320 94776 11360
rect 17452 10900 17492 10940
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 58540 10564 58580 10604
rect 65408 10564 65448 10604
rect 65490 10564 65530 10604
rect 65572 10564 65612 10604
rect 65654 10564 65694 10604
rect 65736 10564 65776 10604
rect 80528 10564 80568 10604
rect 80610 10564 80650 10604
rect 80692 10564 80732 10604
rect 80774 10564 80814 10604
rect 80856 10564 80896 10604
rect 95648 10564 95688 10604
rect 95730 10564 95770 10604
rect 95812 10564 95852 10604
rect 95894 10564 95934 10604
rect 95976 10564 96016 10604
rect 19852 10480 19892 10520
rect 12076 10228 12116 10268
rect 35596 10228 35636 10268
rect 82444 10228 82484 10268
rect 82636 10228 82676 10268
rect 16204 10060 16244 10100
rect 37900 10060 37940 10100
rect 60364 10060 60404 10100
rect 74380 10060 74420 10100
rect 88588 10060 88628 10100
rect 32044 9976 32084 10016
rect 38668 9976 38708 10016
rect 75628 9976 75668 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 15148 9808 15188 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 64168 9808 64208 9848
rect 64250 9808 64290 9848
rect 64332 9808 64372 9848
rect 64414 9808 64454 9848
rect 64496 9808 64536 9848
rect 79288 9808 79328 9848
rect 79370 9808 79410 9848
rect 79452 9808 79492 9848
rect 79534 9808 79574 9848
rect 79616 9808 79656 9848
rect 94408 9808 94448 9848
rect 94490 9808 94530 9848
rect 94572 9808 94612 9848
rect 94654 9808 94694 9848
rect 94736 9808 94776 9848
rect 69484 9640 69524 9680
rect 75244 9556 75284 9596
rect 45292 9304 45332 9344
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 24460 9052 24500 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 65408 9052 65448 9092
rect 65490 9052 65530 9092
rect 65572 9052 65612 9092
rect 65654 9052 65694 9092
rect 65736 9052 65776 9092
rect 78412 9052 78452 9092
rect 80528 9052 80568 9092
rect 80610 9052 80650 9092
rect 80692 9052 80732 9092
rect 80774 9052 80814 9092
rect 80856 9052 80896 9092
rect 82252 9052 82292 9092
rect 89356 9052 89396 9092
rect 95648 9052 95688 9092
rect 95730 9052 95770 9092
rect 95812 9052 95852 9092
rect 95894 9052 95934 9092
rect 95976 9052 96016 9092
rect 26380 8968 26420 9008
rect 24940 8884 24980 8924
rect 81100 8884 81140 8924
rect 81580 8884 81620 8924
rect 12556 8800 12596 8840
rect 22156 8800 22196 8840
rect 31660 8800 31700 8840
rect 55084 8800 55124 8840
rect 56812 8800 56852 8840
rect 59692 8800 59732 8840
rect 70540 8800 70580 8840
rect 73036 8800 73076 8840
rect 75052 8800 75092 8840
rect 9004 8716 9044 8756
rect 15148 8716 15188 8756
rect 81868 8884 81908 8924
rect 82060 8800 82100 8840
rect 88876 8800 88916 8840
rect 33772 8716 33812 8756
rect 49996 8716 50036 8756
rect 66988 8716 67028 8756
rect 35212 8632 35252 8672
rect 54988 8632 55028 8672
rect 56812 8632 56852 8672
rect 83692 8632 83732 8672
rect 28108 8548 28148 8588
rect 49516 8548 49556 8588
rect 55852 8548 55892 8588
rect 71020 8548 71060 8588
rect 78796 8464 78836 8504
rect 35212 8380 35252 8420
rect 83788 8380 83828 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 37036 8296 37076 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 55084 8296 55124 8336
rect 64168 8296 64208 8336
rect 64250 8296 64290 8336
rect 64332 8296 64372 8336
rect 64414 8296 64454 8336
rect 64496 8296 64536 8336
rect 70636 8296 70676 8336
rect 79288 8296 79328 8336
rect 79370 8296 79410 8336
rect 79452 8296 79492 8336
rect 79534 8296 79574 8336
rect 79616 8296 79656 8336
rect 94408 8296 94448 8336
rect 94490 8296 94530 8336
rect 94572 8296 94612 8336
rect 94654 8296 94694 8336
rect 94736 8296 94776 8336
rect 83692 8212 83732 8252
rect 57964 8128 58004 8168
rect 88684 8128 88724 8168
rect 89260 8128 89300 8168
rect 31948 8044 31988 8084
rect 32428 7960 32468 8000
rect 37228 7960 37268 8000
rect 56812 8044 56852 8084
rect 59980 8044 60020 8084
rect 74860 8044 74900 8084
rect 81676 8044 81716 8084
rect 45292 7960 45332 8000
rect 45580 7960 45620 8000
rect 33004 7876 33044 7916
rect 33196 7876 33236 7916
rect 36172 7876 36212 7916
rect 42124 7876 42164 7916
rect 44044 7876 44084 7916
rect 46924 7876 46964 7916
rect 62668 7876 62708 7916
rect 66796 7876 66836 7916
rect 67660 7876 67700 7916
rect 72076 7876 72116 7916
rect 85612 7876 85652 7916
rect 17452 7792 17492 7832
rect 24652 7792 24692 7832
rect 30892 7792 30932 7832
rect 31276 7792 31316 7832
rect 31852 7792 31892 7832
rect 32044 7792 32084 7832
rect 45100 7792 45140 7832
rect 54892 7708 54932 7748
rect 59692 7708 59732 7748
rect 88876 7708 88916 7748
rect 22828 7624 22868 7664
rect 36844 7624 36884 7664
rect 44332 7624 44372 7664
rect 75820 7624 75860 7664
rect 78412 7624 78452 7664
rect 83788 7624 83828 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 19372 7540 19412 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 65408 7540 65448 7580
rect 65490 7540 65530 7580
rect 65572 7540 65612 7580
rect 65654 7540 65694 7580
rect 65736 7540 65776 7580
rect 74860 7540 74900 7580
rect 77068 7540 77108 7580
rect 80528 7540 80568 7580
rect 80610 7540 80650 7580
rect 80692 7540 80732 7580
rect 80774 7540 80814 7580
rect 80856 7540 80896 7580
rect 82924 7540 82964 7580
rect 88396 7540 88436 7580
rect 88588 7540 88628 7580
rect 89356 7540 89396 7580
rect 95648 7540 95688 7580
rect 95730 7540 95770 7580
rect 95812 7540 95852 7580
rect 95894 7540 95934 7580
rect 95976 7540 96016 7580
rect 30124 7456 30164 7496
rect 33772 7456 33812 7496
rect 37900 7456 37940 7496
rect 19276 7372 19316 7412
rect 34444 7288 34484 7328
rect 56236 7288 56276 7328
rect 59692 7288 59732 7328
rect 59884 7372 59924 7412
rect 60268 7288 60308 7328
rect 64012 7456 64052 7496
rect 88204 7456 88244 7496
rect 88684 7456 88724 7496
rect 74956 7372 74996 7412
rect 78892 7372 78932 7412
rect 71020 7288 71060 7328
rect 88204 7288 88244 7328
rect 22924 7204 22964 7244
rect 25708 7204 25748 7244
rect 30028 7204 30068 7244
rect 33772 7204 33812 7244
rect 40108 7204 40148 7244
rect 63052 7204 63092 7244
rect 64492 7204 64532 7244
rect 66796 7204 66836 7244
rect 81868 7204 81908 7244
rect 83692 7204 83732 7244
rect 36460 7120 36500 7160
rect 34540 7036 34580 7076
rect 46348 7120 46388 7160
rect 51820 7036 51860 7076
rect 88204 7036 88244 7076
rect 23500 6952 23540 6992
rect 34828 6952 34868 6992
rect 37516 6952 37556 6992
rect 48940 6952 48980 6992
rect 59980 6952 60020 6992
rect 74092 6952 74132 6992
rect 12556 6868 12596 6908
rect 36460 6868 36500 6908
rect 55756 6868 55796 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 26956 6784 26996 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34732 6784 34772 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 56140 6868 56180 6908
rect 75052 6868 75092 6908
rect 55564 6784 55604 6824
rect 64168 6784 64208 6824
rect 64250 6784 64290 6824
rect 64332 6784 64372 6824
rect 64414 6784 64454 6824
rect 64496 6784 64536 6824
rect 79288 6784 79328 6824
rect 79370 6784 79410 6824
rect 79452 6784 79492 6824
rect 79534 6784 79574 6824
rect 79616 6784 79656 6824
rect 94408 6784 94448 6824
rect 94490 6784 94530 6824
rect 94572 6784 94612 6824
rect 94654 6784 94694 6824
rect 94736 6784 94776 6824
rect 16204 6700 16244 6740
rect 23404 6700 23444 6740
rect 24556 6700 24596 6740
rect 48940 6616 48980 6656
rect 71980 6616 72020 6656
rect 76300 6616 76340 6656
rect 77548 6616 77588 6656
rect 80428 6616 80468 6656
rect 84268 6616 84308 6656
rect 35692 6532 35732 6572
rect 38476 6532 38516 6572
rect 56908 6532 56948 6572
rect 57388 6532 57428 6572
rect 60748 6532 60788 6572
rect 66988 6532 67028 6572
rect 67180 6532 67220 6572
rect 79852 6532 79892 6572
rect 82348 6532 82388 6572
rect 19948 6364 19988 6404
rect 30124 6364 30164 6404
rect 35788 6364 35828 6404
rect 45676 6364 45716 6404
rect 19756 6280 19796 6320
rect 32908 6280 32948 6320
rect 33772 6280 33812 6320
rect 34348 6280 34388 6320
rect 36172 6280 36212 6320
rect 37900 6280 37940 6320
rect 55660 6448 55700 6488
rect 54988 6364 55028 6404
rect 60076 6364 60116 6404
rect 69388 6364 69428 6404
rect 81964 6448 82004 6488
rect 82252 6448 82292 6488
rect 82156 6364 82196 6404
rect 34252 6196 34292 6236
rect 37324 6196 37364 6236
rect 14476 6112 14516 6152
rect 24652 6112 24692 6152
rect 57292 6280 57332 6320
rect 57580 6280 57620 6320
rect 71020 6280 71060 6320
rect 71308 6280 71348 6320
rect 71980 6280 72020 6320
rect 73036 6280 73076 6320
rect 77836 6280 77876 6320
rect 79948 6280 79988 6320
rect 82828 6280 82868 6320
rect 83788 6280 83828 6320
rect 32140 6112 32180 6152
rect 34924 6112 34964 6152
rect 57004 6196 57044 6236
rect 57196 6196 57236 6236
rect 58060 6196 58100 6236
rect 72748 6196 72788 6236
rect 74956 6196 74996 6236
rect 76876 6196 76916 6236
rect 37708 6112 37748 6152
rect 41548 6112 41588 6152
rect 45100 6112 45140 6152
rect 55756 6112 55796 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 23020 6028 23060 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 38188 6028 38228 6068
rect 57868 6112 57908 6152
rect 38476 6028 38516 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 65408 6028 65448 6068
rect 65490 6028 65530 6068
rect 65572 6028 65612 6068
rect 65654 6028 65694 6068
rect 65736 6028 65776 6068
rect 24556 5944 24596 5984
rect 73804 6028 73844 6068
rect 80528 6028 80568 6068
rect 80610 6028 80650 6068
rect 80692 6028 80732 6068
rect 80774 6028 80814 6068
rect 80856 6028 80896 6068
rect 36172 5944 36212 5984
rect 60268 5944 60308 5984
rect 68332 5944 68372 5984
rect 72940 5944 72980 5984
rect 81676 5944 81716 5984
rect 19180 5860 19220 5900
rect 23884 5860 23924 5900
rect 26956 5860 26996 5900
rect 30028 5860 30068 5900
rect 33100 5860 33140 5900
rect 34444 5860 34484 5900
rect 36076 5860 36116 5900
rect 82540 5944 82580 5984
rect 95648 6028 95688 6068
rect 95730 6028 95770 6068
rect 95812 6028 95852 6068
rect 95894 6028 95934 6068
rect 95976 6028 96016 6068
rect 61996 5860 62036 5900
rect 83884 5860 83924 5900
rect 15628 5692 15668 5732
rect 31276 5776 31316 5816
rect 15820 5692 15860 5732
rect 23308 5692 23348 5732
rect 1708 5608 1748 5648
rect 34924 5608 34964 5648
rect 35980 5608 36020 5648
rect 55852 5776 55892 5816
rect 57484 5776 57524 5816
rect 67852 5776 67892 5816
rect 72940 5776 72980 5816
rect 58252 5692 58292 5732
rect 61228 5692 61268 5732
rect 64588 5692 64628 5732
rect 76588 5692 76628 5732
rect 81868 5692 81908 5732
rect 84364 5692 84404 5732
rect 88396 5692 88436 5732
rect 19948 5524 19988 5564
rect 33772 5524 33812 5564
rect 43660 5608 43700 5648
rect 18700 5440 18740 5480
rect 20620 5440 20660 5480
rect 21580 5440 21620 5480
rect 33676 5440 33716 5480
rect 36556 5440 36596 5480
rect 37324 5440 37364 5480
rect 37708 5440 37748 5480
rect 55660 5524 55700 5564
rect 56524 5524 56564 5564
rect 56716 5608 56756 5648
rect 66796 5608 66836 5648
rect 81772 5608 81812 5648
rect 82156 5608 82196 5648
rect 97516 5608 97556 5648
rect 57676 5524 57716 5564
rect 60460 5524 60500 5564
rect 74476 5524 74516 5564
rect 75052 5524 75092 5564
rect 41740 5440 41780 5480
rect 58252 5440 58292 5480
rect 61900 5440 61940 5480
rect 17356 5356 17396 5396
rect 19468 5356 19508 5396
rect 20716 5356 20756 5396
rect 39916 5356 39956 5396
rect 41068 5356 41108 5396
rect 52204 5356 52244 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 22924 5272 22964 5312
rect 28396 5272 28436 5312
rect 56140 5356 56180 5396
rect 57676 5356 57716 5396
rect 61708 5356 61748 5396
rect 71980 5440 72020 5480
rect 72556 5440 72596 5480
rect 72940 5440 72980 5480
rect 70348 5356 70388 5396
rect 70828 5356 70868 5396
rect 72652 5356 72692 5396
rect 80140 5524 80180 5564
rect 75916 5440 75956 5480
rect 77836 5440 77876 5480
rect 79756 5440 79796 5480
rect 80620 5440 80660 5480
rect 81868 5440 81908 5480
rect 28588 5272 28628 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 49900 5272 49940 5312
rect 20812 5188 20852 5228
rect 23980 5188 24020 5228
rect 24364 5188 24404 5228
rect 40300 5188 40340 5228
rect 41644 5188 41684 5228
rect 56620 5188 56660 5228
rect 57100 5188 57140 5228
rect 57292 5272 57332 5312
rect 58156 5272 58196 5312
rect 64168 5272 64208 5312
rect 64250 5272 64290 5312
rect 64332 5272 64372 5312
rect 64414 5272 64454 5312
rect 64496 5272 64536 5312
rect 81484 5356 81524 5396
rect 76108 5272 76148 5312
rect 79288 5272 79328 5312
rect 79370 5272 79410 5312
rect 79452 5272 79492 5312
rect 79534 5272 79574 5312
rect 79616 5272 79656 5312
rect 81676 5272 81716 5312
rect 94408 5272 94448 5312
rect 94490 5272 94530 5312
rect 94572 5272 94612 5312
rect 94654 5272 94694 5312
rect 94736 5272 94776 5312
rect 64012 5188 64052 5228
rect 67852 5188 67892 5228
rect 69004 5188 69044 5228
rect 38092 5104 38132 5144
rect 68620 5104 68660 5144
rect 73708 5104 73748 5144
rect 76684 5104 76724 5144
rect 19660 5020 19700 5060
rect 21388 5020 21428 5060
rect 21964 5020 22004 5060
rect 28588 5020 28628 5060
rect 44236 5020 44276 5060
rect 57484 5020 57524 5060
rect 2092 4936 2132 4976
rect 2476 4936 2516 4976
rect 24844 4936 24884 4976
rect 28780 4936 28820 4976
rect 57868 5020 57908 5060
rect 68716 5020 68756 5060
rect 71884 5020 71924 5060
rect 34540 4936 34580 4976
rect 38188 4936 38228 4976
rect 47308 4936 47348 4976
rect 48364 4936 48404 4976
rect 15628 4684 15668 4724
rect 17548 4852 17588 4892
rect 19948 4852 19988 4892
rect 21292 4852 21332 4892
rect 27628 4852 27668 4892
rect 23308 4768 23348 4808
rect 18508 4684 18548 4724
rect 19372 4684 19412 4724
rect 21196 4684 21236 4724
rect 25516 4768 25556 4808
rect 31468 4768 31508 4808
rect 22348 4684 22388 4724
rect 24844 4684 24884 4724
rect 25036 4684 25076 4724
rect 30604 4684 30644 4724
rect 17164 4600 17204 4640
rect 35500 4852 35540 4892
rect 37036 4852 37076 4892
rect 37228 4852 37268 4892
rect 38860 4768 38900 4808
rect 17356 4600 17396 4640
rect 23212 4600 23252 4640
rect 33484 4600 33524 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20716 4516 20756 4556
rect 28780 4516 28820 4556
rect 34252 4516 34292 4556
rect 49516 4852 49556 4892
rect 56620 4936 56660 4976
rect 58252 4936 58292 4976
rect 57484 4852 57524 4892
rect 39052 4768 39092 4808
rect 35500 4684 35540 4724
rect 35980 4684 36020 4724
rect 67948 4936 67988 4976
rect 76012 4936 76052 4976
rect 76780 4936 76820 4976
rect 87052 4936 87092 4976
rect 87724 4936 87764 4976
rect 88492 4936 88532 4976
rect 97708 4936 97748 4976
rect 98092 4936 98132 4976
rect 63244 4852 63284 4892
rect 56236 4684 56276 4724
rect 56812 4684 56852 4724
rect 68236 4768 68276 4808
rect 72076 4768 72116 4808
rect 72652 4852 72692 4892
rect 73420 4852 73460 4892
rect 77260 4852 77300 4892
rect 77548 4852 77588 4892
rect 85804 4852 85844 4892
rect 85612 4768 85652 4808
rect 56524 4600 56564 4640
rect 67564 4600 67604 4640
rect 68620 4600 68660 4640
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 61708 4516 61748 4556
rect 65408 4516 65448 4556
rect 65490 4516 65530 4556
rect 65572 4516 65612 4556
rect 65654 4516 65694 4556
rect 65736 4516 65776 4556
rect 68716 4516 68756 4556
rect 70732 4684 70772 4724
rect 71212 4684 71252 4724
rect 72652 4684 72692 4724
rect 72844 4684 72884 4724
rect 76780 4684 76820 4724
rect 81292 4684 81332 4724
rect 88972 4684 89012 4724
rect 69964 4600 70004 4640
rect 74092 4600 74132 4640
rect 75148 4600 75188 4640
rect 71884 4516 71924 4556
rect 80428 4516 80468 4556
rect 80528 4516 80568 4556
rect 80610 4516 80650 4556
rect 80692 4516 80732 4556
rect 80774 4516 80814 4556
rect 80856 4516 80896 4556
rect 95648 4516 95688 4556
rect 95730 4516 95770 4556
rect 95812 4516 95852 4556
rect 95894 4516 95934 4556
rect 95976 4516 96016 4556
rect 17356 4432 17396 4472
rect 19372 4432 19412 4472
rect 21196 4432 21236 4472
rect 36556 4432 36596 4472
rect 39052 4432 39092 4472
rect 55564 4432 55604 4472
rect 56716 4432 56756 4472
rect 73036 4432 73076 4472
rect 77260 4432 77300 4472
rect 24652 4348 24692 4388
rect 35020 4348 35060 4388
rect 35788 4348 35828 4388
rect 37804 4348 37844 4388
rect 50380 4348 50420 4388
rect 55276 4348 55316 4388
rect 55852 4348 55892 4388
rect 61804 4348 61844 4388
rect 70444 4348 70484 4388
rect 22732 4264 22772 4304
rect 23404 4264 23444 4304
rect 31468 4264 31508 4304
rect 31660 4264 31700 4304
rect 65452 4264 65492 4304
rect 66892 4264 66932 4304
rect 67084 4264 67124 4304
rect 19564 4180 19604 4220
rect 20236 4180 20276 4220
rect 23788 4180 23828 4220
rect 24940 4180 24980 4220
rect 28396 4180 28436 4220
rect 29932 4180 29972 4220
rect 49132 4180 49172 4220
rect 49612 4180 49652 4220
rect 7084 4096 7124 4136
rect 12076 4096 12116 4136
rect 25708 4096 25748 4136
rect 17164 4012 17204 4052
rect 23980 4012 24020 4052
rect 19756 3928 19796 3968
rect 19948 3928 19988 3968
rect 30604 4096 30644 4136
rect 32908 4096 32948 4136
rect 34060 4096 34100 4136
rect 39052 4096 39092 4136
rect 41452 4096 41492 4136
rect 42604 4096 42644 4136
rect 42988 4096 43028 4136
rect 43372 4096 43412 4136
rect 54124 4096 54164 4136
rect 81772 4348 81812 4388
rect 85900 4348 85940 4388
rect 57964 4180 58004 4220
rect 64780 4180 64820 4220
rect 73420 4180 73460 4220
rect 77548 4180 77588 4220
rect 56812 4096 56852 4136
rect 47308 4012 47348 4052
rect 60460 4012 60500 4052
rect 29068 3928 29108 3968
rect 31276 3928 31316 3968
rect 49516 3928 49556 3968
rect 49708 3928 49748 3968
rect 49900 3844 49940 3884
rect 55852 3844 55892 3884
rect 61996 4096 62036 4136
rect 66220 4096 66260 4136
rect 68620 4096 68660 4136
rect 69004 4096 69044 4136
rect 69484 4096 69524 4136
rect 70444 4096 70484 4136
rect 75244 4096 75284 4136
rect 75628 4096 75668 4136
rect 79756 4096 79796 4136
rect 86284 4096 86324 4136
rect 64780 4012 64820 4052
rect 66412 4012 66452 4052
rect 73516 4012 73556 4052
rect 75724 4012 75764 4052
rect 77260 4012 77300 4052
rect 60556 3928 60596 3968
rect 66892 3928 66932 3968
rect 70540 3928 70580 3968
rect 71788 3928 71828 3968
rect 84268 3928 84308 3968
rect 58540 3844 58580 3884
rect 62092 3844 62132 3884
rect 66796 3844 66836 3884
rect 68236 3844 68276 3884
rect 70732 3844 70772 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 23884 3760 23924 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 35596 3760 35636 3800
rect 38092 3760 38132 3800
rect 40300 3760 40340 3800
rect 41068 3760 41108 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 57100 3760 57140 3800
rect 64168 3760 64208 3800
rect 64250 3760 64290 3800
rect 64332 3760 64372 3800
rect 64414 3760 64454 3800
rect 64496 3760 64536 3800
rect 67084 3760 67124 3800
rect 67852 3760 67892 3800
rect 14476 3676 14516 3716
rect 16396 3676 16436 3716
rect 20140 3676 20180 3716
rect 20332 3676 20372 3716
rect 20620 3676 20660 3716
rect 24460 3676 24500 3716
rect 25420 3592 25460 3632
rect 26380 3592 26420 3632
rect 75148 3844 75188 3884
rect 86860 3844 86900 3884
rect 68332 3760 68372 3800
rect 75340 3760 75380 3800
rect 77068 3760 77108 3800
rect 79288 3760 79328 3800
rect 79370 3760 79410 3800
rect 79452 3760 79492 3800
rect 79534 3760 79574 3800
rect 79616 3760 79656 3800
rect 79756 3760 79796 3800
rect 81484 3760 81524 3800
rect 94408 3760 94448 3800
rect 94490 3760 94530 3800
rect 94572 3760 94612 3800
rect 94654 3760 94694 3800
rect 94736 3760 94776 3800
rect 63436 3592 63476 3632
rect 19852 3508 19892 3548
rect 20908 3508 20948 3548
rect 21580 3508 21620 3548
rect 60268 3508 60308 3548
rect 1228 3424 1268 3464
rect 1612 3424 1652 3464
rect 1996 3424 2036 3464
rect 2380 3424 2420 3464
rect 6220 3424 6260 3464
rect 6988 3424 7028 3464
rect 16204 3424 16244 3464
rect 17164 3424 17204 3464
rect 17452 3424 17492 3464
rect 18508 3424 18548 3464
rect 19276 3424 19316 3464
rect 21964 3424 22004 3464
rect 22156 3424 22196 3464
rect 23500 3424 23540 3464
rect 28108 3424 28148 3464
rect 31948 3424 31988 3464
rect 18700 3340 18740 3380
rect 32140 3424 32180 3464
rect 36076 3424 36116 3464
rect 36556 3424 36596 3464
rect 43372 3424 43412 3464
rect 47980 3424 48020 3464
rect 56908 3424 56948 3464
rect 30028 3340 30068 3380
rect 34348 3340 34388 3380
rect 20332 3256 20372 3296
rect 20812 3256 20852 3296
rect 20716 3172 20756 3212
rect 20908 3088 20948 3128
rect 63820 3676 63860 3716
rect 80620 3676 80660 3716
rect 63724 3592 63764 3632
rect 76588 3592 76628 3632
rect 81868 3592 81908 3632
rect 57388 3424 57428 3464
rect 58156 3424 58196 3464
rect 60748 3424 60788 3464
rect 67468 3424 67508 3464
rect 69388 3424 69428 3464
rect 70348 3424 70388 3464
rect 76300 3424 76340 3464
rect 76780 3424 76820 3464
rect 80140 3424 80180 3464
rect 89260 3424 89300 3464
rect 94732 3424 94772 3464
rect 95116 3424 95156 3464
rect 95500 3424 95540 3464
rect 95884 3424 95924 3464
rect 96652 3424 96692 3464
rect 97420 3424 97460 3464
rect 97804 3424 97844 3464
rect 97996 3424 98036 3464
rect 70828 3340 70868 3380
rect 85708 3340 85748 3380
rect 86092 3340 86132 3380
rect 37804 3256 37844 3296
rect 39724 3256 39764 3296
rect 49228 3256 49268 3296
rect 49612 3256 49652 3296
rect 63148 3256 63188 3296
rect 63820 3256 63860 3296
rect 34732 3088 34772 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 68236 3256 68276 3296
rect 70636 3256 70676 3296
rect 72748 3256 72788 3296
rect 75820 3256 75860 3296
rect 41548 3172 41588 3212
rect 59500 3172 59540 3212
rect 60556 3172 60596 3212
rect 55276 3088 55316 3128
rect 78796 3172 78836 3212
rect 87052 3172 87092 3212
rect 19660 3004 19700 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 54124 3004 54164 3044
rect 63148 3004 63188 3044
rect 65408 3004 65448 3044
rect 65490 3004 65530 3044
rect 65572 3004 65612 3044
rect 65654 3004 65694 3044
rect 65736 3004 65776 3044
rect 80528 3004 80568 3044
rect 80610 3004 80650 3044
rect 80692 3004 80732 3044
rect 80774 3004 80814 3044
rect 80856 3004 80896 3044
rect 17164 2920 17204 2960
rect 54892 2920 54932 2960
rect 19468 2836 19508 2876
rect 33676 2836 33716 2876
rect 34540 2836 34580 2876
rect 41548 2836 41588 2876
rect 57196 2836 57236 2876
rect 61900 2836 61940 2876
rect 19372 2752 19412 2792
rect 46636 2752 46676 2792
rect 73804 2920 73844 2960
rect 81676 3088 81716 3128
rect 81292 3004 81332 3044
rect 95648 3004 95688 3044
rect 95730 3004 95770 3044
rect 95812 3004 95852 3044
rect 95894 3004 95934 3044
rect 95976 3004 96016 3044
rect 81868 2836 81908 2876
rect 46828 2752 46868 2792
rect 60364 2752 60404 2792
rect 16588 2668 16628 2708
rect 38860 2668 38900 2708
rect 16684 2584 16724 2624
rect 75916 2584 75956 2624
rect 85996 2584 86036 2624
rect 21388 2500 21428 2540
rect 76108 2500 76148 2540
rect 87628 2500 87668 2540
rect 15628 2416 15668 2456
rect 85900 2416 85940 2456
rect 86188 2416 86228 2456
rect 62092 2332 62132 2372
rect 87628 2332 87668 2372
rect 16588 2248 16628 2288
rect 56620 2248 56660 2288
rect 71212 2164 71252 2204
rect 21388 2080 21428 2120
rect 16684 1912 16724 1952
rect 86188 1912 86228 1952
rect 71788 1324 71828 1364
rect 79948 1240 79988 1280
rect 85804 1240 85844 1280
rect 35692 1156 35732 1196
rect 85996 1156 86036 1196
rect 20716 820 20756 860
rect 85708 820 85748 860
rect 86092 232 86132 272
rect 79852 148 79892 188
<< metal4 >>
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 18808 11360 19176 11369
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 18808 11311 19176 11320
rect 33928 11360 34296 11369
rect 33968 11320 34010 11360
rect 34050 11320 34092 11360
rect 34132 11320 34174 11360
rect 34214 11320 34256 11360
rect 33928 11311 34296 11320
rect 49048 11360 49416 11369
rect 49088 11320 49130 11360
rect 49170 11320 49212 11360
rect 49252 11320 49294 11360
rect 49334 11320 49376 11360
rect 49048 11311 49416 11320
rect 64168 11360 64536 11369
rect 64208 11320 64250 11360
rect 64290 11320 64332 11360
rect 64372 11320 64414 11360
rect 64454 11320 64496 11360
rect 64168 11311 64536 11320
rect 79288 11360 79656 11369
rect 79328 11320 79370 11360
rect 79410 11320 79452 11360
rect 79492 11320 79534 11360
rect 79574 11320 79616 11360
rect 79288 11311 79656 11320
rect 94408 11360 94776 11369
rect 94448 11320 94490 11360
rect 94530 11320 94572 11360
rect 94612 11320 94654 11360
rect 94694 11320 94736 11360
rect 94408 11311 94776 11320
rect 17452 10940 17492 10949
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 12076 10268 12116 10277
rect 9003 10016 9045 10025
rect 9003 9976 9004 10016
rect 9044 9976 9045 10016
rect 9003 9967 9045 9976
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 9004 8756 9044 9967
rect 9004 8707 9044 8716
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 7083 8168 7125 8177
rect 7083 8128 7084 8168
rect 7124 8128 7125 8168
rect 7083 8119 7125 8128
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 6219 6320 6261 6329
rect 6219 6280 6220 6320
rect 6260 6280 6261 6320
rect 6219 6271 6261 6280
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 1707 5648 1749 5657
rect 1707 5608 1708 5648
rect 1748 5608 1749 5648
rect 1707 5599 1749 5608
rect 1708 5514 1748 5599
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 2091 4976 2133 4985
rect 2091 4936 2092 4976
rect 2132 4936 2133 4976
rect 2091 4927 2133 4936
rect 2476 4976 2516 4985
rect 2092 4842 2132 4927
rect 2476 4481 2516 4936
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 2475 4472 2517 4481
rect 2475 4432 2476 4472
rect 2516 4432 2517 4472
rect 2475 4423 2517 4432
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 1228 3464 1268 3473
rect 1228 3305 1268 3424
rect 1611 3464 1653 3473
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 1995 3464 2037 3473
rect 1995 3424 1996 3464
rect 2036 3424 2037 3464
rect 1995 3415 2037 3424
rect 2379 3464 2421 3473
rect 2379 3424 2380 3464
rect 2420 3424 2421 3464
rect 2379 3415 2421 3424
rect 6220 3464 6260 6271
rect 7084 4136 7124 8119
rect 7084 4087 7124 4096
rect 12076 4136 12116 10228
rect 16204 10100 16244 10109
rect 15148 9848 15188 9857
rect 12556 8840 12596 8849
rect 12556 6908 12596 8800
rect 15148 8756 15188 9808
rect 15148 8707 15188 8716
rect 16204 8177 16244 10060
rect 17452 9437 17492 10900
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 50288 10604 50656 10613
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50288 10555 50656 10564
rect 58540 10604 58580 10613
rect 19852 10520 19892 10529
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 17451 9428 17493 9437
rect 17451 9388 17452 9428
rect 17492 9388 17493 9428
rect 17451 9379 17493 9388
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 16203 8168 16245 8177
rect 16203 8128 16204 8168
rect 16244 8128 16245 8168
rect 16203 8119 16245 8128
rect 12556 6859 12596 6868
rect 17452 7832 17492 7841
rect 16204 6740 16244 6749
rect 12076 4087 12116 4096
rect 14476 6152 14516 6161
rect 14476 3716 14516 6112
rect 15628 5732 15668 5741
rect 15820 5732 15860 5741
rect 15668 5692 15820 5732
rect 15628 5683 15668 5692
rect 15820 5683 15860 5692
rect 14476 3667 14516 3676
rect 15628 4724 15668 4733
rect 6987 3632 7029 3641
rect 6987 3592 6988 3632
rect 7028 3592 7029 3632
rect 6987 3583 7029 3592
rect 6220 3415 6260 3424
rect 6988 3464 7028 3583
rect 6988 3415 7028 3424
rect 1612 3330 1652 3415
rect 1996 3330 2036 3415
rect 2380 3330 2420 3415
rect 1227 3296 1269 3305
rect 1227 3256 1228 3296
rect 1268 3256 1269 3296
rect 1227 3247 1269 3256
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 15628 2456 15668 4684
rect 16204 3464 16244 6700
rect 17356 5396 17396 5405
rect 17164 4640 17204 4649
rect 17164 4052 17204 4600
rect 17356 4640 17396 5356
rect 17356 4591 17396 4600
rect 17356 4472 17396 4481
rect 17356 4313 17396 4432
rect 17355 4304 17397 4313
rect 17355 4264 17356 4304
rect 17396 4264 17397 4304
rect 17355 4255 17397 4264
rect 17164 4003 17204 4012
rect 16204 3415 16244 3424
rect 16396 3716 16436 3725
rect 16396 3389 16436 3676
rect 17164 3464 17204 3473
rect 16395 3380 16437 3389
rect 16395 3340 16396 3380
rect 16436 3340 16437 3380
rect 16395 3331 16437 3340
rect 17164 2960 17204 3424
rect 17452 3464 17492 7792
rect 19372 7580 19412 7589
rect 19276 7412 19316 7421
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19179 5900 19221 5909
rect 19179 5860 19180 5900
rect 19220 5860 19221 5900
rect 19179 5851 19221 5860
rect 19180 5766 19220 5851
rect 18700 5480 18740 5489
rect 17547 4892 17589 4901
rect 17547 4852 17548 4892
rect 17588 4852 17589 4892
rect 17547 4843 17589 4852
rect 17548 4758 17588 4843
rect 18507 4724 18549 4733
rect 18507 4684 18508 4724
rect 18548 4684 18549 4724
rect 18507 4675 18549 4684
rect 18508 4590 18548 4675
rect 17452 3415 17492 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18508 3330 18548 3415
rect 18700 3380 18740 5440
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3464 19316 7372
rect 19372 4724 19412 7540
rect 19755 6320 19797 6329
rect 19755 6280 19756 6320
rect 19796 6280 19797 6320
rect 19755 6271 19797 6280
rect 19756 6186 19796 6271
rect 19372 4675 19412 4684
rect 19468 5396 19508 5405
rect 19276 3415 19316 3424
rect 19372 4472 19412 4481
rect 18700 3331 18740 3340
rect 17164 2911 17204 2920
rect 19372 2792 19412 4432
rect 19468 2876 19508 5356
rect 19660 5060 19700 5069
rect 19563 4220 19605 4229
rect 19563 4180 19564 4220
rect 19604 4180 19605 4220
rect 19563 4171 19605 4180
rect 19564 4086 19604 4171
rect 19660 3044 19700 5020
rect 19756 3968 19796 3977
rect 19756 3557 19796 3928
rect 19755 3548 19797 3557
rect 19755 3508 19756 3548
rect 19796 3508 19797 3548
rect 19755 3499 19797 3508
rect 19852 3548 19892 10480
rect 35596 10268 35636 10277
rect 32043 10016 32085 10025
rect 32043 9976 32044 10016
rect 32084 9976 32085 10016
rect 32043 9967 32085 9976
rect 32044 9882 32084 9967
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 24460 9092 24500 9101
rect 22156 8840 22196 8849
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19948 6404 19988 6413
rect 19948 5564 19988 6364
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19948 5515 19988 5524
rect 20620 5480 20660 5489
rect 19948 4892 19988 4901
rect 19948 4229 19988 4852
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19947 4220 19989 4229
rect 19947 4180 19948 4220
rect 19988 4180 19989 4220
rect 19947 4171 19989 4180
rect 20235 4220 20277 4229
rect 20235 4180 20236 4220
rect 20276 4180 20277 4220
rect 20235 4171 20277 4180
rect 20236 4086 20276 4171
rect 19852 3499 19892 3508
rect 19948 3968 19988 3977
rect 19948 3305 19988 3928
rect 20139 3716 20181 3725
rect 20139 3676 20140 3716
rect 20180 3676 20181 3716
rect 20139 3667 20181 3676
rect 20332 3716 20372 3725
rect 20140 3582 20180 3667
rect 19947 3296 19989 3305
rect 19947 3256 19948 3296
rect 19988 3256 19989 3296
rect 19947 3247 19989 3256
rect 20332 3296 20372 3676
rect 20620 3716 20660 5440
rect 21580 5480 21620 5489
rect 20716 5396 20756 5405
rect 20716 4556 20756 5356
rect 20716 4507 20756 4516
rect 20812 5228 20852 5237
rect 20620 3667 20660 3676
rect 20332 3247 20372 3256
rect 20812 3296 20852 5188
rect 21387 5060 21429 5069
rect 21387 5020 21388 5060
rect 21428 5020 21429 5060
rect 21387 5011 21429 5020
rect 21388 4926 21428 5011
rect 21292 4892 21332 4903
rect 21292 4817 21332 4852
rect 21291 4808 21333 4817
rect 21291 4768 21292 4808
rect 21332 4768 21333 4808
rect 21291 4759 21333 4768
rect 21196 4724 21236 4733
rect 21196 4472 21236 4684
rect 21196 4423 21236 4432
rect 21292 4229 21332 4759
rect 21291 4220 21333 4229
rect 21291 4180 21292 4220
rect 21332 4180 21333 4220
rect 21291 4171 21333 4180
rect 20812 3247 20852 3256
rect 20908 3548 20948 3557
rect 20716 3212 20756 3221
rect 19660 2995 19700 3004
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19468 2827 19508 2836
rect 19372 2743 19412 2752
rect 15628 2407 15668 2416
rect 16588 2708 16628 2717
rect 16588 2288 16628 2668
rect 16588 2239 16628 2248
rect 16684 2624 16724 2633
rect 16684 1952 16724 2584
rect 16684 1903 16724 1912
rect 20716 860 20756 3172
rect 20908 3128 20948 3508
rect 21580 3548 21620 5440
rect 21580 3499 21620 3508
rect 21964 5060 22004 5069
rect 21964 3464 22004 5020
rect 21964 3415 22004 3424
rect 22156 3464 22196 8800
rect 22828 7664 22868 7673
rect 22828 6488 22868 7624
rect 22923 7244 22965 7253
rect 22923 7204 22924 7244
rect 22964 7204 22965 7244
rect 22923 7195 22965 7204
rect 23307 7244 23349 7253
rect 23307 7204 23308 7244
rect 23348 7204 23349 7244
rect 23307 7195 23349 7204
rect 22924 7110 22964 7195
rect 22923 6488 22965 6497
rect 22828 6448 22924 6488
rect 22964 6448 22965 6488
rect 22923 6439 22965 6448
rect 22924 5312 22964 6439
rect 23020 6068 23060 6077
rect 23020 5909 23060 6028
rect 23019 5900 23061 5909
rect 23019 5860 23020 5900
rect 23060 5860 23061 5900
rect 23019 5851 23061 5860
rect 23308 5732 23348 7195
rect 23500 6992 23540 7001
rect 23308 5683 23348 5692
rect 23404 6740 23444 6749
rect 22924 5263 22964 5272
rect 23308 4808 23348 4817
rect 23212 4768 23308 4808
rect 22348 4724 22388 4733
rect 22348 3641 22388 4684
rect 23212 4640 23252 4768
rect 23308 4759 23348 4768
rect 23212 4591 23252 4600
rect 22731 4304 22773 4313
rect 22731 4264 22732 4304
rect 22772 4264 22773 4304
rect 22731 4255 22773 4264
rect 23404 4304 23444 6700
rect 23404 4255 23444 4264
rect 22732 4170 22772 4255
rect 22347 3632 22389 3641
rect 22347 3592 22348 3632
rect 22388 3592 22389 3632
rect 22347 3583 22389 3592
rect 22156 3415 22196 3424
rect 23500 3464 23540 6952
rect 23884 5900 23924 5909
rect 23788 4220 23828 4231
rect 23788 4145 23828 4180
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 23884 3800 23924 5860
rect 23980 5228 24020 5237
rect 23980 4052 24020 5188
rect 24364 5228 24404 5237
rect 24364 4901 24404 5188
rect 24363 4892 24405 4901
rect 24363 4852 24364 4892
rect 24404 4852 24405 4892
rect 24363 4843 24405 4852
rect 23980 4003 24020 4012
rect 23884 3751 23924 3760
rect 24460 3716 24500 9052
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 26380 9008 26420 9017
rect 24940 8924 24980 8933
rect 24652 7832 24692 7841
rect 24556 6740 24596 6749
rect 24556 5984 24596 6700
rect 24652 6581 24692 7792
rect 24651 6572 24693 6581
rect 24651 6532 24652 6572
rect 24692 6532 24693 6572
rect 24651 6523 24693 6532
rect 24652 6152 24692 6523
rect 24652 6103 24692 6112
rect 24556 5935 24596 5944
rect 24651 5060 24693 5069
rect 24651 5020 24652 5060
rect 24692 5020 24693 5060
rect 24651 5011 24693 5020
rect 24652 4388 24692 5011
rect 24844 4976 24884 4985
rect 24844 4724 24884 4936
rect 24844 4675 24884 4684
rect 24652 4339 24692 4348
rect 24940 4220 24980 8884
rect 25708 7244 25748 7253
rect 25515 4808 25557 4817
rect 25515 4768 25516 4808
rect 25556 4768 25557 4808
rect 25515 4759 25557 4768
rect 25035 4724 25077 4733
rect 25035 4684 25036 4724
rect 25076 4684 25077 4724
rect 25035 4675 25077 4684
rect 25036 4590 25076 4675
rect 25516 4674 25556 4759
rect 24940 4171 24980 4180
rect 25708 4136 25748 7204
rect 25708 4087 25748 4096
rect 24460 3667 24500 3676
rect 25420 3632 25460 3641
rect 25420 3473 25460 3592
rect 26380 3632 26420 8968
rect 31660 8840 31700 8849
rect 28108 8588 28148 8597
rect 26956 6824 26996 6833
rect 26956 5909 26996 6784
rect 26955 5900 26997 5909
rect 26955 5860 26956 5900
rect 26996 5860 26997 5900
rect 26955 5851 26997 5860
rect 26956 5766 26996 5851
rect 27627 4892 27669 4901
rect 27627 4852 27628 4892
rect 27668 4852 27669 4892
rect 27627 4843 27669 4852
rect 27628 4145 27668 4843
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 26380 3583 26420 3592
rect 23500 3415 23540 3424
rect 25419 3464 25461 3473
rect 25419 3424 25420 3464
rect 25460 3424 25461 3464
rect 25419 3415 25461 3424
rect 28108 3464 28148 8548
rect 30892 7832 30932 7841
rect 30124 7496 30164 7505
rect 30124 7253 30164 7456
rect 30028 7244 30068 7253
rect 30028 6329 30068 7204
rect 30123 7244 30165 7253
rect 30123 7204 30124 7244
rect 30164 7204 30165 7244
rect 30123 7195 30165 7204
rect 30124 6413 30164 7195
rect 30123 6404 30165 6413
rect 30123 6364 30124 6404
rect 30164 6364 30165 6404
rect 30123 6355 30165 6364
rect 30027 6320 30069 6329
rect 30027 6280 30028 6320
rect 30068 6280 30069 6320
rect 30027 6271 30069 6280
rect 30124 6270 30164 6355
rect 30028 5900 30068 5909
rect 28396 5312 28436 5321
rect 28396 4220 28436 5272
rect 28588 5312 28628 5321
rect 28588 5060 28628 5272
rect 28588 4229 28628 5020
rect 28780 4976 28820 4985
rect 28780 4556 28820 4936
rect 28780 4507 28820 4516
rect 28396 4171 28436 4180
rect 28587 4220 28629 4229
rect 28587 4180 28588 4220
rect 28628 4180 28629 4220
rect 28587 4171 28629 4180
rect 29932 4220 29972 4231
rect 29932 4145 29972 4180
rect 29931 4136 29973 4145
rect 29931 4096 29932 4136
rect 29972 4096 29973 4136
rect 29931 4087 29973 4096
rect 29067 3968 29109 3977
rect 29067 3928 29068 3968
rect 29108 3928 29109 3968
rect 29067 3919 29109 3928
rect 29068 3834 29108 3919
rect 28108 3415 28148 3424
rect 30028 3380 30068 5860
rect 30892 5657 30932 7792
rect 31275 7832 31317 7841
rect 31275 7792 31276 7832
rect 31316 7792 31317 7832
rect 31275 7783 31317 7792
rect 31276 7698 31316 7783
rect 31276 5816 31316 5825
rect 30891 5648 30933 5657
rect 30891 5608 30892 5648
rect 30932 5608 30933 5648
rect 30891 5599 30933 5608
rect 30604 4724 30644 4733
rect 30604 4136 30644 4684
rect 30604 4087 30644 4096
rect 31276 3968 31316 5776
rect 31468 4808 31508 4817
rect 31468 4304 31508 4768
rect 31468 4255 31508 4264
rect 31660 4304 31700 8800
rect 33772 8756 33812 8765
rect 31948 8084 31988 8093
rect 31852 7832 31892 7841
rect 31852 5825 31892 7792
rect 31851 5816 31893 5825
rect 31851 5776 31852 5816
rect 31892 5776 31893 5816
rect 31851 5767 31893 5776
rect 31660 4255 31700 4264
rect 31276 3919 31316 3928
rect 31948 3464 31988 8044
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 32428 7866 32468 7951
rect 33004 7916 33044 7925
rect 32043 7832 32085 7841
rect 32043 7792 32044 7832
rect 32084 7792 32085 7832
rect 32043 7783 32085 7792
rect 32044 7698 32084 7783
rect 32908 6320 32948 6329
rect 31948 3415 31988 3424
rect 32140 6152 32180 6161
rect 32140 3464 32180 6112
rect 32715 5564 32757 5573
rect 32715 5524 32716 5564
rect 32756 5524 32757 5564
rect 32715 5515 32757 5524
rect 32716 4733 32756 5515
rect 32715 4724 32757 4733
rect 32715 4684 32716 4724
rect 32756 4684 32757 4724
rect 32715 4675 32757 4684
rect 32908 4136 32948 6280
rect 32908 4087 32948 4096
rect 33004 3557 33044 7876
rect 33195 7916 33237 7925
rect 33195 7876 33196 7916
rect 33236 7876 33237 7916
rect 33195 7867 33237 7876
rect 33196 7782 33236 7867
rect 33772 7496 33812 8716
rect 35212 8672 35252 8681
rect 35212 8420 35252 8632
rect 35212 8371 35252 8380
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 33772 7447 33812 7456
rect 34444 7328 34484 7337
rect 33772 7244 33812 7253
rect 33772 6320 33812 7204
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 33099 5900 33141 5909
rect 33099 5860 33100 5900
rect 33140 5860 33141 5900
rect 33099 5851 33141 5860
rect 33100 5766 33140 5851
rect 33772 5564 33812 6280
rect 34348 6320 34388 6329
rect 34252 6236 34292 6245
rect 34252 5741 34292 6196
rect 34251 5732 34293 5741
rect 34251 5692 34252 5732
rect 34292 5692 34293 5732
rect 34251 5683 34293 5692
rect 33772 5515 33812 5524
rect 33676 5480 33716 5489
rect 33484 4640 33524 4649
rect 33484 3725 33524 4600
rect 33483 3716 33525 3725
rect 33483 3676 33484 3716
rect 33524 3676 33525 3716
rect 33483 3667 33525 3676
rect 33003 3548 33045 3557
rect 33003 3508 33004 3548
rect 33044 3508 33045 3548
rect 33003 3499 33045 3508
rect 32140 3415 32180 3424
rect 30028 3331 30068 3340
rect 20908 3079 20948 3088
rect 33676 2876 33716 5440
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34251 4976 34293 4985
rect 34251 4936 34252 4976
rect 34292 4936 34293 4976
rect 34251 4927 34293 4936
rect 34252 4556 34292 4927
rect 34252 4507 34292 4516
rect 34059 4136 34101 4145
rect 34059 4096 34060 4136
rect 34100 4096 34101 4136
rect 34059 4087 34101 4096
rect 34060 4002 34100 4087
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34348 3380 34388 6280
rect 34444 5900 34484 7288
rect 34444 5851 34484 5860
rect 34540 7076 34580 7085
rect 34540 4976 34580 7036
rect 34828 6992 34868 7001
rect 34540 4927 34580 4936
rect 34732 6824 34772 6833
rect 34539 4136 34581 4145
rect 34539 4096 34540 4136
rect 34580 4096 34581 4136
rect 34539 4087 34581 4096
rect 34348 3331 34388 3340
rect 33676 2827 33716 2836
rect 34540 2876 34580 4087
rect 34732 3128 34772 6784
rect 34828 4901 34868 6952
rect 34924 6152 34964 6161
rect 34924 5909 34964 6112
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 34923 5900 34965 5909
rect 34923 5860 34924 5900
rect 34964 5860 34965 5900
rect 34923 5851 34965 5860
rect 34924 5648 34964 5657
rect 34827 4892 34869 4901
rect 34827 4852 34828 4892
rect 34868 4852 34869 4892
rect 34827 4843 34869 4852
rect 34924 4145 34964 5608
rect 35500 4892 35540 4901
rect 35500 4724 35540 4852
rect 35500 4675 35540 4684
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35019 4388 35061 4397
rect 35019 4348 35020 4388
rect 35060 4348 35061 4388
rect 35019 4339 35061 4348
rect 35020 4254 35060 4339
rect 34923 4136 34965 4145
rect 34923 4096 34924 4136
rect 34964 4096 34965 4136
rect 34923 4087 34965 4096
rect 35596 3800 35636 10228
rect 37899 10100 37941 10109
rect 37899 10060 37900 10100
rect 37940 10060 37941 10100
rect 37899 10051 37941 10060
rect 48363 10100 48405 10109
rect 48363 10060 48364 10100
rect 48404 10060 48405 10100
rect 48363 10051 48405 10060
rect 37900 9966 37940 10051
rect 38668 10016 38708 10025
rect 37036 8336 37076 8345
rect 36172 7916 36212 7925
rect 36172 7085 36212 7876
rect 36844 7664 36884 7673
rect 36460 7160 36500 7169
rect 36171 7076 36213 7085
rect 36171 7036 36172 7076
rect 36212 7036 36213 7076
rect 36171 7027 36213 7036
rect 36460 6908 36500 7120
rect 35596 3751 35636 3760
rect 35692 6572 35732 6581
rect 34732 3079 34772 3088
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 34540 2827 34580 2836
rect 21388 2540 21428 2549
rect 21388 2120 21428 2500
rect 21388 2071 21428 2080
rect 35692 1196 35732 6532
rect 35787 6488 35829 6497
rect 35787 6448 35788 6488
rect 35828 6448 35829 6488
rect 35787 6439 35829 6448
rect 35788 6404 35828 6439
rect 35788 6353 35828 6364
rect 36460 6329 36500 6868
rect 36844 6497 36884 7624
rect 36843 6488 36885 6497
rect 36843 6448 36844 6488
rect 36884 6448 36885 6488
rect 36843 6439 36885 6448
rect 36172 6320 36212 6329
rect 36172 5984 36212 6280
rect 36459 6320 36501 6329
rect 36459 6280 36460 6320
rect 36500 6280 36501 6320
rect 36459 6271 36501 6280
rect 36172 5935 36212 5944
rect 36076 5900 36116 5909
rect 35980 5648 36020 5657
rect 35787 4724 35829 4733
rect 35787 4684 35788 4724
rect 35828 4684 35829 4724
rect 35787 4675 35829 4684
rect 35980 4724 36020 5608
rect 35980 4675 36020 4684
rect 35788 4388 35828 4675
rect 35788 4339 35828 4348
rect 36076 3464 36116 5860
rect 36651 5816 36693 5825
rect 36651 5776 36652 5816
rect 36692 5776 36693 5816
rect 36651 5767 36693 5776
rect 36555 5480 36597 5489
rect 36555 5440 36556 5480
rect 36596 5440 36597 5480
rect 36555 5431 36597 5440
rect 36556 5346 36596 5431
rect 36076 3415 36116 3424
rect 36556 4472 36596 4481
rect 36556 3464 36596 4432
rect 36652 4145 36692 5767
rect 37036 4892 37076 8296
rect 37036 4843 37076 4852
rect 37228 8000 37268 8009
rect 37228 4892 37268 7960
rect 37900 7496 37940 7505
rect 37515 6992 37557 7001
rect 37515 6952 37516 6992
rect 37556 6952 37557 6992
rect 37515 6943 37557 6952
rect 37516 6858 37556 6943
rect 37900 6581 37940 7456
rect 37899 6572 37941 6581
rect 37899 6532 37900 6572
rect 37940 6532 37941 6572
rect 37899 6523 37941 6532
rect 38476 6572 38516 6581
rect 37707 6404 37749 6413
rect 37707 6364 37708 6404
rect 37748 6364 37749 6404
rect 37707 6355 37749 6364
rect 37324 6236 37364 6245
rect 37324 5480 37364 6196
rect 37708 6152 37748 6355
rect 37900 6320 37940 6523
rect 37900 6271 37940 6280
rect 37708 6103 37748 6112
rect 38188 6068 38228 6077
rect 37324 5431 37364 5440
rect 37708 5480 37748 5489
rect 37228 4843 37268 4852
rect 36651 4136 36693 4145
rect 36651 4096 36652 4136
rect 36692 4096 36693 4136
rect 36651 4087 36693 4096
rect 37708 3473 37748 5440
rect 38092 5144 38132 5153
rect 37804 4388 37844 4397
rect 36556 3415 36596 3424
rect 37707 3464 37749 3473
rect 37707 3424 37708 3464
rect 37748 3424 37749 3464
rect 37707 3415 37749 3424
rect 37804 3296 37844 4348
rect 38092 3800 38132 5104
rect 38188 4976 38228 6028
rect 38476 6068 38516 6532
rect 38476 6019 38516 6028
rect 38188 4927 38228 4936
rect 38668 3809 38708 9976
rect 45292 9344 45332 9353
rect 45292 8009 45332 9304
rect 45579 8084 45621 8093
rect 45579 8044 45580 8084
rect 45620 8044 45621 8084
rect 45579 8035 45621 8044
rect 42603 8000 42645 8009
rect 42603 7960 42604 8000
rect 42644 7960 42645 8000
rect 42603 7951 42645 7960
rect 45291 8000 45333 8009
rect 45291 7960 45292 8000
rect 45332 7960 45333 8000
rect 45291 7951 45333 7960
rect 45580 8000 45620 8035
rect 42123 7916 42165 7925
rect 42123 7876 42124 7916
rect 42164 7876 42165 7916
rect 42123 7867 42165 7876
rect 42124 7782 42164 7867
rect 41451 7748 41493 7757
rect 41451 7708 41452 7748
rect 41492 7708 41493 7748
rect 41451 7699 41493 7708
rect 40107 7244 40149 7253
rect 40107 7204 40108 7244
rect 40148 7204 40149 7244
rect 40107 7195 40149 7204
rect 40108 7110 40148 7195
rect 39915 5900 39957 5909
rect 39915 5860 39916 5900
rect 39956 5860 39957 5900
rect 39915 5851 39957 5860
rect 39916 5396 39956 5851
rect 40299 5732 40341 5741
rect 40299 5692 40300 5732
rect 40340 5692 40341 5732
rect 40299 5683 40341 5692
rect 39916 5347 39956 5356
rect 40300 5228 40340 5683
rect 40300 5179 40340 5188
rect 41068 5396 41108 5405
rect 39723 4892 39765 4901
rect 39723 4852 39724 4892
rect 39764 4852 39765 4892
rect 39723 4843 39765 4852
rect 38860 4808 38900 4817
rect 38092 3751 38132 3760
rect 38667 3800 38709 3809
rect 38667 3760 38668 3800
rect 38708 3760 38709 3800
rect 38667 3751 38709 3760
rect 37804 3247 37844 3256
rect 38860 2708 38900 4768
rect 39052 4808 39092 4817
rect 39052 4472 39092 4768
rect 39052 4136 39092 4432
rect 39052 4087 39092 4096
rect 39724 3296 39764 4843
rect 40299 3800 40341 3809
rect 40299 3760 40300 3800
rect 40340 3760 40341 3800
rect 40299 3751 40341 3760
rect 41068 3800 41108 5356
rect 41452 4136 41492 7699
rect 41643 6992 41685 7001
rect 41643 6952 41644 6992
rect 41684 6952 41685 6992
rect 41643 6943 41685 6952
rect 41547 6320 41589 6329
rect 41547 6280 41548 6320
rect 41588 6280 41589 6320
rect 41547 6271 41589 6280
rect 41548 6152 41588 6271
rect 41548 6103 41588 6112
rect 41644 5228 41684 6943
rect 41739 5480 41781 5489
rect 41739 5440 41740 5480
rect 41780 5440 41781 5480
rect 41739 5431 41781 5440
rect 41740 5346 41780 5431
rect 41644 5179 41684 5188
rect 41452 4087 41492 4096
rect 42604 4136 42644 7951
rect 44043 7916 44085 7925
rect 44043 7876 44044 7916
rect 44084 7876 44085 7916
rect 44043 7867 44085 7876
rect 43371 7832 43413 7841
rect 43371 7792 43372 7832
rect 43412 7792 43413 7832
rect 43371 7783 43413 7792
rect 42604 4087 42644 4096
rect 42987 4136 43029 4145
rect 42987 4096 42988 4136
rect 43028 4096 43029 4136
rect 42987 4087 43029 4096
rect 43372 4136 43412 7783
rect 44044 7782 44084 7867
rect 45292 7866 45332 7951
rect 45580 7949 45620 7960
rect 46924 7916 46964 7925
rect 45100 7832 45140 7841
rect 44331 7664 44373 7673
rect 44331 7624 44332 7664
rect 44372 7624 44373 7664
rect 44331 7615 44373 7624
rect 44332 7530 44372 7615
rect 45100 6152 45140 7792
rect 46924 7757 46964 7876
rect 46923 7748 46965 7757
rect 46923 7708 46924 7748
rect 46964 7708 46965 7748
rect 46923 7699 46965 7708
rect 46348 7160 46388 7200
rect 46348 7085 46388 7120
rect 46347 7076 46389 7085
rect 46347 7036 46348 7076
rect 46388 7036 46389 7076
rect 46347 7027 46389 7036
rect 45675 6572 45717 6581
rect 45675 6532 45676 6572
rect 45716 6532 45717 6572
rect 45675 6523 45717 6532
rect 45676 6404 45716 6523
rect 45676 6355 45716 6364
rect 45100 6103 45140 6112
rect 46348 5909 46388 7027
rect 46347 5900 46389 5909
rect 46347 5860 46348 5900
rect 46388 5860 46389 5900
rect 46347 5851 46389 5860
rect 43659 5648 43701 5657
rect 43659 5608 43660 5648
rect 43700 5608 43701 5648
rect 43659 5599 43701 5608
rect 43660 5514 43700 5599
rect 44236 5060 44276 5069
rect 44236 4901 44276 5020
rect 47308 4976 47348 4985
rect 44235 4892 44277 4901
rect 44235 4852 44236 4892
rect 44276 4852 44277 4892
rect 44235 4843 44277 4852
rect 43372 4087 43412 4096
rect 42988 4002 43028 4087
rect 47308 4052 47348 4936
rect 48364 4976 48404 10051
rect 49048 9848 49416 9857
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49048 9799 49416 9808
rect 49995 9428 50037 9437
rect 49995 9388 49996 9428
rect 50036 9388 50037 9428
rect 49995 9379 50037 9388
rect 49996 8756 50036 9379
rect 50288 9092 50656 9101
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50288 9043 50656 9052
rect 49996 8707 50036 8716
rect 55084 8840 55124 8849
rect 54988 8672 55028 8681
rect 49516 8588 49556 8597
rect 49048 8336 49416 8345
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49048 8287 49416 8296
rect 48940 6992 48980 7001
rect 48940 6656 48980 6952
rect 49048 6824 49416 6833
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49048 6775 49416 6784
rect 48940 6245 48980 6616
rect 48939 6236 48981 6245
rect 48939 6196 48940 6236
rect 48980 6196 48981 6236
rect 48939 6187 48981 6196
rect 49048 5312 49416 5321
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49048 5263 49416 5272
rect 48364 4927 48404 4936
rect 49516 4892 49556 8548
rect 54892 7748 54932 7757
rect 50288 7580 50656 7589
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50288 7531 50656 7540
rect 51819 7244 51861 7253
rect 51819 7204 51820 7244
rect 51860 7204 51861 7244
rect 51819 7195 51861 7204
rect 51820 7076 51860 7195
rect 51820 7027 51860 7036
rect 50288 6068 50656 6077
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50288 6019 50656 6028
rect 52203 5396 52245 5405
rect 52203 5356 52204 5396
rect 52244 5356 52245 5396
rect 52203 5347 52245 5356
rect 49516 4843 49556 4852
rect 49900 5312 49940 5321
rect 49131 4220 49173 4229
rect 49131 4180 49132 4220
rect 49172 4180 49173 4220
rect 49131 4171 49173 4180
rect 49612 4220 49652 4229
rect 49132 4086 49172 4171
rect 47308 4003 47348 4012
rect 49516 3968 49556 3977
rect 41068 3751 41108 3760
rect 49048 3800 49416 3809
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49048 3751 49416 3760
rect 40300 3666 40340 3751
rect 49516 3557 49556 3928
rect 49515 3548 49557 3557
rect 49515 3508 49516 3548
rect 49556 3508 49557 3548
rect 49515 3499 49557 3508
rect 43371 3464 43413 3473
rect 43371 3424 43372 3464
rect 43412 3424 43413 3464
rect 43371 3415 43413 3424
rect 47979 3464 48021 3473
rect 47979 3424 47980 3464
rect 48020 3424 48021 3464
rect 47979 3415 48021 3424
rect 43372 3330 43412 3415
rect 47980 3330 48020 3415
rect 39724 3247 39764 3256
rect 49227 3296 49269 3305
rect 49227 3256 49228 3296
rect 49268 3256 49269 3296
rect 49227 3247 49269 3256
rect 49612 3296 49652 4180
rect 49707 3968 49749 3977
rect 49707 3928 49708 3968
rect 49748 3928 49749 3968
rect 49707 3919 49749 3928
rect 49708 3834 49748 3919
rect 49900 3884 49940 5272
rect 52204 5262 52244 5347
rect 50288 4556 50656 4565
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50288 4507 50656 4516
rect 50379 4388 50421 4397
rect 50379 4348 50380 4388
rect 50420 4348 50421 4388
rect 50379 4339 50421 4348
rect 50380 4254 50420 4339
rect 49900 3835 49940 3844
rect 54124 4136 54164 4145
rect 49612 3247 49652 3256
rect 41548 3212 41588 3221
rect 41548 2876 41588 3172
rect 49228 3162 49268 3247
rect 50288 3044 50656 3053
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50288 2995 50656 3004
rect 54124 3044 54164 4096
rect 54124 2995 54164 3004
rect 54892 2960 54932 7708
rect 54988 6404 55028 8632
rect 55084 8336 55124 8800
rect 56812 8840 56852 8849
rect 56812 8672 56852 8800
rect 55084 8287 55124 8296
rect 55852 8588 55892 8597
rect 55756 6908 55796 6917
rect 55564 6824 55604 6833
rect 54988 6355 55028 6364
rect 55467 6404 55509 6413
rect 55467 6364 55468 6404
rect 55508 6364 55509 6404
rect 55467 6355 55509 6364
rect 55371 6320 55413 6329
rect 55371 6280 55372 6320
rect 55412 6280 55413 6320
rect 55371 6271 55413 6280
rect 55372 6161 55412 6271
rect 55468 6161 55508 6355
rect 55371 6152 55413 6161
rect 55371 6112 55372 6152
rect 55412 6112 55413 6152
rect 55371 6103 55413 6112
rect 55467 6152 55509 6161
rect 55467 6112 55468 6152
rect 55508 6112 55509 6152
rect 55467 6103 55509 6112
rect 55564 4472 55604 6784
rect 55660 6488 55700 6497
rect 55660 5564 55700 6448
rect 55756 6152 55796 6868
rect 55756 6103 55796 6112
rect 55852 5816 55892 8548
rect 56812 8084 56852 8632
rect 56812 8035 56852 8044
rect 57964 8168 58004 8177
rect 56236 7328 56276 7337
rect 55852 5767 55892 5776
rect 56140 6908 56180 6917
rect 55660 5515 55700 5524
rect 56140 5396 56180 6868
rect 56140 5347 56180 5356
rect 56236 4724 56276 7288
rect 56908 6572 56948 6581
rect 56716 5648 56756 5657
rect 56236 4675 56276 4684
rect 56524 5564 56564 5573
rect 56524 4640 56564 5524
rect 56619 5564 56661 5573
rect 56619 5524 56620 5564
rect 56660 5524 56661 5564
rect 56619 5515 56661 5524
rect 56620 5228 56660 5515
rect 56620 5179 56660 5188
rect 56524 4591 56564 4600
rect 56620 4976 56660 4985
rect 55564 4423 55604 4432
rect 55276 4388 55316 4397
rect 55276 3128 55316 4348
rect 55852 4388 55892 4397
rect 55852 3884 55892 4348
rect 55852 3835 55892 3844
rect 55276 3079 55316 3088
rect 54892 2911 54932 2920
rect 41548 2827 41588 2836
rect 46636 2792 46676 2801
rect 46828 2792 46868 2801
rect 46676 2752 46828 2792
rect 46636 2743 46676 2752
rect 46828 2743 46868 2752
rect 38860 2659 38900 2668
rect 56620 2288 56660 4936
rect 56716 4472 56756 5608
rect 56716 4423 56756 4432
rect 56812 4724 56852 4733
rect 56812 4136 56852 4684
rect 56812 4087 56852 4096
rect 56908 3464 56948 6532
rect 57388 6572 57428 6581
rect 57003 6320 57045 6329
rect 57003 6280 57004 6320
rect 57044 6280 57045 6320
rect 57003 6271 57045 6280
rect 57292 6320 57332 6329
rect 57004 6236 57044 6271
rect 57004 6185 57044 6196
rect 57196 6236 57236 6245
rect 57100 5228 57140 5237
rect 57100 3800 57140 5188
rect 57100 3751 57140 3760
rect 56908 3415 56948 3424
rect 57196 2876 57236 6196
rect 57292 5312 57332 6280
rect 57292 5263 57332 5272
rect 57388 3464 57428 6532
rect 57579 6320 57621 6329
rect 57579 6280 57580 6320
rect 57620 6280 57621 6320
rect 57579 6271 57621 6280
rect 57580 6186 57620 6271
rect 57868 6152 57908 6161
rect 57484 5816 57524 5825
rect 57484 5060 57524 5776
rect 57676 5564 57716 5573
rect 57676 5396 57716 5524
rect 57676 5347 57716 5356
rect 57484 5011 57524 5020
rect 57868 5060 57908 6112
rect 57868 5011 57908 5020
rect 57484 4892 57524 4901
rect 57964 4892 58004 8128
rect 57524 4852 58004 4892
rect 58060 6236 58100 6245
rect 57484 4843 57524 4852
rect 57963 4220 58005 4229
rect 57963 4180 57964 4220
rect 58004 4180 58005 4220
rect 57963 4171 58005 4180
rect 57964 4086 58004 4171
rect 57388 3415 57428 3424
rect 58060 3305 58100 6196
rect 58252 5732 58292 5741
rect 58252 5480 58292 5692
rect 58252 5431 58292 5440
rect 58156 5312 58196 5321
rect 58156 3464 58196 5272
rect 58252 4976 58292 4985
rect 58252 3977 58292 4936
rect 58251 3968 58293 3977
rect 58251 3928 58252 3968
rect 58292 3928 58293 3968
rect 58251 3919 58293 3928
rect 58540 3884 58580 10564
rect 65408 10604 65776 10613
rect 65448 10564 65490 10604
rect 65530 10564 65572 10604
rect 65612 10564 65654 10604
rect 65694 10564 65736 10604
rect 65408 10555 65776 10564
rect 80528 10604 80896 10613
rect 80568 10564 80610 10604
rect 80650 10564 80692 10604
rect 80732 10564 80774 10604
rect 80814 10564 80856 10604
rect 80528 10555 80896 10564
rect 95648 10604 96016 10613
rect 95688 10564 95730 10604
rect 95770 10564 95812 10604
rect 95852 10564 95894 10604
rect 95934 10564 95976 10604
rect 95648 10555 96016 10564
rect 82444 10268 82484 10277
rect 82636 10268 82676 10277
rect 82484 10228 82636 10268
rect 82444 10219 82484 10228
rect 82636 10219 82676 10228
rect 60364 10100 60404 10109
rect 59692 8840 59732 8849
rect 59692 7748 59732 8800
rect 59692 7699 59732 7708
rect 59980 8084 60020 8093
rect 59884 7412 59924 7421
rect 59692 7328 59732 7337
rect 59884 7328 59924 7372
rect 59732 7288 59924 7328
rect 59692 7279 59732 7288
rect 59980 6992 60020 8044
rect 59980 6943 60020 6952
rect 60268 7328 60308 7337
rect 60075 6404 60117 6413
rect 60075 6364 60076 6404
rect 60116 6364 60117 6404
rect 60075 6355 60117 6364
rect 60076 6270 60116 6355
rect 60268 5984 60308 7288
rect 60268 5935 60308 5944
rect 58540 3835 58580 3844
rect 58156 3415 58196 3424
rect 60268 3548 60308 3557
rect 60268 3305 60308 3508
rect 58059 3296 58101 3305
rect 58059 3256 58060 3296
rect 58100 3256 58101 3296
rect 58059 3247 58101 3256
rect 60267 3296 60309 3305
rect 60267 3256 60268 3296
rect 60308 3256 60309 3296
rect 60267 3247 60309 3256
rect 59499 3212 59541 3221
rect 59499 3172 59500 3212
rect 59540 3172 59541 3212
rect 59499 3163 59541 3172
rect 59500 3078 59540 3163
rect 57196 2827 57236 2836
rect 60364 2792 60404 10060
rect 74380 10100 74420 10109
rect 64168 9848 64536 9857
rect 64208 9808 64250 9848
rect 64290 9808 64332 9848
rect 64372 9808 64414 9848
rect 64454 9808 64496 9848
rect 64168 9799 64536 9808
rect 69484 9680 69524 9689
rect 65408 9092 65776 9101
rect 65448 9052 65490 9092
rect 65530 9052 65572 9092
rect 65612 9052 65654 9092
rect 65694 9052 65736 9092
rect 65408 9043 65776 9052
rect 66988 8756 67028 8765
rect 64168 8336 64536 8345
rect 64208 8296 64250 8336
rect 64290 8296 64332 8336
rect 64372 8296 64414 8336
rect 64454 8296 64496 8336
rect 64168 8287 64536 8296
rect 62667 8084 62709 8093
rect 62667 8044 62668 8084
rect 62708 8044 62709 8084
rect 62667 8035 62709 8044
rect 62668 7916 62708 8035
rect 66988 8009 67028 8716
rect 67467 8756 67509 8765
rect 67467 8716 67468 8756
rect 67508 8716 67509 8756
rect 67467 8707 67509 8716
rect 66987 8000 67029 8009
rect 66987 7960 66988 8000
rect 67028 7960 67029 8000
rect 66987 7951 67029 7960
rect 62668 7867 62708 7876
rect 66796 7916 66836 7925
rect 66699 7832 66741 7841
rect 66796 7832 66836 7876
rect 66699 7792 66700 7832
rect 66740 7792 66836 7832
rect 66699 7783 66741 7792
rect 64491 7748 64533 7757
rect 64491 7708 64492 7748
rect 64532 7708 64533 7748
rect 64491 7699 64533 7708
rect 64012 7496 64052 7505
rect 63052 7244 63092 7253
rect 60747 6572 60789 6581
rect 60747 6532 60748 6572
rect 60788 6532 60789 6572
rect 60747 6523 60789 6532
rect 60748 6438 60788 6523
rect 63052 5909 63092 7204
rect 61996 5900 62036 5909
rect 61227 5732 61269 5741
rect 61227 5692 61228 5732
rect 61268 5692 61269 5732
rect 61227 5683 61269 5692
rect 61228 5598 61268 5683
rect 60459 5564 60501 5573
rect 60459 5524 60460 5564
rect 60500 5524 60501 5564
rect 60459 5515 60501 5524
rect 60460 5430 60500 5515
rect 61900 5480 61940 5489
rect 61708 5396 61748 5405
rect 61708 4556 61748 5356
rect 61708 4507 61748 4516
rect 61803 4388 61845 4397
rect 61803 4348 61804 4388
rect 61844 4348 61845 4388
rect 61803 4339 61845 4348
rect 61804 4254 61844 4339
rect 60460 4052 60500 4061
rect 60460 3557 60500 4012
rect 60556 3968 60596 3977
rect 60459 3548 60501 3557
rect 60459 3508 60460 3548
rect 60500 3508 60501 3548
rect 60459 3499 60501 3508
rect 60556 3212 60596 3928
rect 60747 3464 60789 3473
rect 60747 3424 60748 3464
rect 60788 3424 60789 3464
rect 60747 3415 60789 3424
rect 60748 3330 60788 3415
rect 60556 3163 60596 3172
rect 61900 2876 61940 5440
rect 61996 4136 62036 5860
rect 63051 5900 63093 5909
rect 63051 5860 63052 5900
rect 63092 5860 63093 5900
rect 63051 5851 63093 5860
rect 64012 5228 64052 7456
rect 64492 7244 64532 7699
rect 65408 7580 65776 7589
rect 65448 7540 65490 7580
rect 65530 7540 65572 7580
rect 65612 7540 65654 7580
rect 65694 7540 65736 7580
rect 65408 7531 65776 7540
rect 64492 7195 64532 7204
rect 66796 7244 66836 7253
rect 64168 6824 64536 6833
rect 64208 6784 64250 6824
rect 64290 6784 64332 6824
rect 64372 6784 64414 6824
rect 64454 6784 64496 6824
rect 64168 6775 64536 6784
rect 66796 6245 66836 7204
rect 66987 6572 67029 6581
rect 66987 6532 66988 6572
rect 67028 6532 67029 6572
rect 66987 6523 67029 6532
rect 67180 6572 67220 6583
rect 66988 6438 67028 6523
rect 67180 6497 67220 6532
rect 67179 6488 67221 6497
rect 67179 6448 67180 6488
rect 67220 6448 67221 6488
rect 67179 6439 67221 6448
rect 66795 6236 66837 6245
rect 66795 6196 66796 6236
rect 66836 6196 66837 6236
rect 66795 6187 66837 6196
rect 65408 6068 65776 6077
rect 65448 6028 65490 6068
rect 65530 6028 65572 6068
rect 65612 6028 65654 6068
rect 65694 6028 65736 6068
rect 65408 6019 65776 6028
rect 64588 5732 64628 5741
rect 64588 5489 64628 5692
rect 66796 5648 66836 5657
rect 64587 5480 64629 5489
rect 64587 5440 64588 5480
rect 64628 5440 64629 5480
rect 64587 5431 64629 5440
rect 64168 5312 64536 5321
rect 64208 5272 64250 5312
rect 64290 5272 64332 5312
rect 64372 5272 64414 5312
rect 64454 5272 64496 5312
rect 64168 5263 64536 5272
rect 64012 5179 64052 5188
rect 63243 4892 63285 4901
rect 63243 4852 63244 4892
rect 63284 4852 63285 4892
rect 63243 4843 63285 4852
rect 63244 4758 63284 4843
rect 65408 4556 65776 4565
rect 65448 4516 65490 4556
rect 65530 4516 65572 4556
rect 65612 4516 65654 4556
rect 65694 4516 65736 4556
rect 65408 4507 65776 4516
rect 64780 4229 64820 4314
rect 65451 4304 65493 4313
rect 65451 4264 65452 4304
rect 65492 4264 65493 4304
rect 65451 4255 65493 4264
rect 64779 4220 64821 4229
rect 64779 4180 64780 4220
rect 64820 4180 64821 4220
rect 64779 4171 64821 4180
rect 65452 4170 65492 4255
rect 61996 4087 62036 4096
rect 66220 4136 66260 4145
rect 64780 4052 64820 4061
rect 66220 4052 66260 4096
rect 66412 4052 66452 4061
rect 66220 4012 66412 4052
rect 61900 2827 61940 2836
rect 62092 3884 62132 3893
rect 60364 2743 60404 2752
rect 62092 2372 62132 3844
rect 64168 3800 64536 3809
rect 64208 3760 64250 3800
rect 64290 3760 64332 3800
rect 64372 3760 64414 3800
rect 64454 3760 64496 3800
rect 64168 3751 64536 3760
rect 63820 3716 63860 3725
rect 63436 3632 63476 3641
rect 63724 3632 63764 3641
rect 63476 3592 63724 3632
rect 63436 3583 63476 3592
rect 63724 3583 63764 3592
rect 63148 3296 63188 3305
rect 63148 3044 63188 3256
rect 63820 3296 63860 3676
rect 64780 3557 64820 4012
rect 66412 4003 66452 4012
rect 66796 3884 66836 5608
rect 66892 4304 66932 4313
rect 66892 3968 66932 4264
rect 67084 4304 67124 4315
rect 67084 4229 67124 4264
rect 67083 4220 67125 4229
rect 67083 4180 67084 4220
rect 67124 4180 67125 4220
rect 67083 4171 67125 4180
rect 66892 3919 66932 3928
rect 66796 3835 66836 3844
rect 67084 3800 67124 3809
rect 67084 3641 67124 3760
rect 67083 3632 67125 3641
rect 67083 3592 67084 3632
rect 67124 3592 67125 3632
rect 67083 3583 67125 3592
rect 64779 3548 64821 3557
rect 64779 3508 64780 3548
rect 64820 3508 64821 3548
rect 64779 3499 64821 3508
rect 67468 3464 67508 8707
rect 67659 7916 67701 7925
rect 67659 7876 67660 7916
rect 67700 7876 67701 7916
rect 67659 7867 67701 7876
rect 67660 7782 67700 7867
rect 69388 6404 69428 6413
rect 68332 5984 68372 5993
rect 67851 5816 67893 5825
rect 67851 5776 67852 5816
rect 67892 5776 67893 5816
rect 67851 5767 67893 5776
rect 67852 5682 67892 5767
rect 67852 5228 67892 5237
rect 67563 4640 67605 4649
rect 67563 4600 67564 4640
rect 67604 4600 67605 4640
rect 67563 4591 67605 4600
rect 67564 4506 67604 4591
rect 67852 3800 67892 5188
rect 67948 4976 67988 4985
rect 67948 4313 67988 4936
rect 68236 4808 68276 4817
rect 67947 4304 67989 4313
rect 67947 4264 67948 4304
rect 67988 4264 67989 4304
rect 67947 4255 67989 4264
rect 67852 3751 67892 3760
rect 68236 3884 68276 4768
rect 67468 3415 67508 3424
rect 63820 3247 63860 3256
rect 68236 3296 68276 3844
rect 68332 3800 68372 5944
rect 69004 5228 69044 5237
rect 68620 5144 68660 5153
rect 68620 4640 68660 5104
rect 68620 4136 68660 4600
rect 68716 5060 68756 5069
rect 68716 4556 68756 5020
rect 68716 4507 68756 4516
rect 68620 4087 68660 4096
rect 69004 4136 69044 5188
rect 69004 4087 69044 4096
rect 68332 3751 68372 3760
rect 69388 3464 69428 6364
rect 69484 4136 69524 9640
rect 70539 8840 70581 8849
rect 70539 8800 70540 8840
rect 70580 8800 70581 8840
rect 70539 8791 70581 8800
rect 73035 8840 73077 8849
rect 73035 8800 73036 8840
rect 73076 8800 73077 8840
rect 73035 8791 73077 8800
rect 70540 8706 70580 8791
rect 73036 8706 73076 8791
rect 71020 8588 71060 8597
rect 70636 8336 70676 8345
rect 70348 5396 70388 5405
rect 69963 4640 70005 4649
rect 69963 4600 69964 4640
rect 70004 4600 70005 4640
rect 69963 4591 70005 4600
rect 69964 4506 70004 4591
rect 69484 4087 69524 4096
rect 69388 3415 69428 3424
rect 70348 3464 70388 5356
rect 70444 4388 70484 4397
rect 70444 4136 70484 4348
rect 70539 4304 70581 4313
rect 70539 4264 70540 4304
rect 70580 4264 70581 4304
rect 70539 4255 70581 4264
rect 70444 4087 70484 4096
rect 70540 3968 70580 4255
rect 70540 3919 70580 3928
rect 70348 3415 70388 3424
rect 68236 3247 68276 3256
rect 70636 3296 70676 8296
rect 71020 7589 71060 8548
rect 72076 7916 72116 7925
rect 71019 7580 71061 7589
rect 71019 7540 71020 7580
rect 71060 7540 71061 7580
rect 71019 7531 71061 7540
rect 71020 7328 71060 7531
rect 71020 7279 71060 7288
rect 71979 6656 72021 6665
rect 71979 6616 71980 6656
rect 72020 6616 72021 6656
rect 71979 6607 72021 6616
rect 71019 6572 71061 6581
rect 71019 6532 71020 6572
rect 71060 6532 71061 6572
rect 71019 6523 71061 6532
rect 71020 6320 71060 6523
rect 71980 6522 72020 6607
rect 71307 6488 71349 6497
rect 71307 6448 71308 6488
rect 71348 6448 71349 6488
rect 71307 6439 71349 6448
rect 71883 6488 71925 6497
rect 71883 6448 71884 6488
rect 71924 6448 71925 6488
rect 71883 6439 71925 6448
rect 71020 6271 71060 6280
rect 71308 6320 71348 6439
rect 71308 6271 71348 6280
rect 70828 5396 70868 5405
rect 70732 4724 70772 4733
rect 70732 3884 70772 4684
rect 70732 3835 70772 3844
rect 70828 3380 70868 5356
rect 71884 5060 71924 6439
rect 71980 6320 72020 6329
rect 72076 6320 72116 7876
rect 74092 6992 74132 7001
rect 72020 6280 72116 6320
rect 73036 6320 73076 6329
rect 71980 5657 72020 6280
rect 72748 6236 72788 6245
rect 71979 5648 72021 5657
rect 71979 5608 71980 5648
rect 72020 5608 72021 5648
rect 71979 5599 72021 5608
rect 71884 5011 71924 5020
rect 71980 5480 72020 5489
rect 70828 3331 70868 3340
rect 71212 4724 71252 4733
rect 70636 3247 70676 3256
rect 63148 2995 63188 3004
rect 65408 3044 65776 3053
rect 65448 3004 65490 3044
rect 65530 3004 65572 3044
rect 65612 3004 65654 3044
rect 65694 3004 65736 3044
rect 65408 2995 65776 3004
rect 62092 2323 62132 2332
rect 56620 2239 56660 2248
rect 71212 2204 71252 4684
rect 71883 4640 71925 4649
rect 71980 4640 72020 5440
rect 72556 5480 72596 5489
rect 72075 4808 72117 4817
rect 72075 4768 72076 4808
rect 72116 4768 72117 4808
rect 72075 4759 72117 4768
rect 72076 4674 72116 4759
rect 71883 4600 71884 4640
rect 71924 4600 72020 4640
rect 71883 4591 71925 4600
rect 71884 4556 71924 4591
rect 71884 4505 71924 4516
rect 72556 4313 72596 5440
rect 72652 5396 72692 5405
rect 72652 4892 72692 5356
rect 72652 4724 72692 4852
rect 72652 4675 72692 4684
rect 72555 4304 72597 4313
rect 72555 4264 72556 4304
rect 72596 4264 72597 4304
rect 72555 4255 72597 4264
rect 71212 2155 71252 2164
rect 71788 3968 71828 3977
rect 71788 1364 71828 3928
rect 72748 3296 72788 6196
rect 72940 5984 72980 5993
rect 72940 5816 72980 5944
rect 72940 5767 72980 5776
rect 72939 5480 72981 5489
rect 72939 5440 72940 5480
rect 72980 5440 72981 5480
rect 72939 5431 72981 5440
rect 72940 5346 72980 5431
rect 72843 4724 72885 4733
rect 72843 4684 72844 4724
rect 72884 4684 72885 4724
rect 72843 4675 72885 4684
rect 72844 4590 72884 4675
rect 73036 4472 73076 6280
rect 73804 6068 73844 6077
rect 73708 5144 73748 5153
rect 73036 4423 73076 4432
rect 73420 4892 73460 4901
rect 73420 4220 73460 4852
rect 73515 4640 73557 4649
rect 73515 4600 73516 4640
rect 73556 4600 73557 4640
rect 73515 4591 73557 4600
rect 73420 4171 73460 4180
rect 73516 4052 73556 4591
rect 73708 4145 73748 5104
rect 73707 4136 73749 4145
rect 73707 4096 73708 4136
rect 73748 4096 73749 4136
rect 73707 4087 73749 4096
rect 73516 4003 73556 4012
rect 72748 3247 72788 3256
rect 73804 2960 73844 6028
rect 74092 4640 74132 6952
rect 74380 5825 74420 10060
rect 88588 10100 88628 10109
rect 75628 10016 75668 10025
rect 75244 9596 75284 9605
rect 75052 8840 75092 8849
rect 75052 8765 75092 8800
rect 75051 8756 75093 8765
rect 75051 8716 75052 8756
rect 75092 8716 75093 8756
rect 75051 8707 75093 8716
rect 75052 8705 75092 8707
rect 74860 8084 74900 8093
rect 74860 7589 74900 8044
rect 74859 7580 74901 7589
rect 74859 7540 74860 7580
rect 74900 7540 74901 7580
rect 74859 7531 74901 7540
rect 74860 7446 74900 7531
rect 74955 7412 74997 7421
rect 74955 7372 74956 7412
rect 74996 7372 74997 7412
rect 74955 7363 74997 7372
rect 74956 6665 74996 7363
rect 75052 6908 75092 6917
rect 74955 6656 74997 6665
rect 74955 6616 74956 6656
rect 74996 6616 74997 6656
rect 74955 6607 74997 6616
rect 74956 6236 74996 6607
rect 74956 6187 74996 6196
rect 74379 5816 74421 5825
rect 74379 5776 74380 5816
rect 74420 5776 74421 5816
rect 74379 5767 74421 5776
rect 74475 5564 74517 5573
rect 74475 5524 74476 5564
rect 74516 5524 74517 5564
rect 74475 5515 74517 5524
rect 75052 5564 75092 6868
rect 75052 5515 75092 5524
rect 74476 5430 74516 5515
rect 75147 5060 75189 5069
rect 75147 5020 75148 5060
rect 75188 5020 75189 5060
rect 75147 5011 75189 5020
rect 74092 4591 74132 4600
rect 75148 4640 75188 5011
rect 75148 4229 75188 4600
rect 75147 4220 75189 4229
rect 75147 4180 75148 4220
rect 75188 4180 75189 4220
rect 75147 4171 75189 4180
rect 75148 3884 75188 4171
rect 75244 4136 75284 9556
rect 75244 4087 75284 4096
rect 75628 4136 75668 9976
rect 79288 9848 79656 9857
rect 79328 9808 79370 9848
rect 79410 9808 79452 9848
rect 79492 9808 79534 9848
rect 79574 9808 79616 9848
rect 79288 9799 79656 9808
rect 78412 9092 78452 9101
rect 75628 4087 75668 4096
rect 75820 7664 75860 7673
rect 75724 4052 75764 4061
rect 75724 3968 75764 4012
rect 75148 3835 75188 3844
rect 75340 3928 75764 3968
rect 75340 3800 75380 3928
rect 75340 3751 75380 3760
rect 75820 3296 75860 7624
rect 78412 7664 78452 9052
rect 80528 9092 80896 9101
rect 80568 9052 80610 9092
rect 80650 9052 80692 9092
rect 80732 9052 80774 9092
rect 80814 9052 80856 9092
rect 80528 9043 80896 9052
rect 82252 9092 82292 9101
rect 81099 9008 81141 9017
rect 81099 8968 81100 9008
rect 81140 8968 81141 9008
rect 81099 8959 81141 8968
rect 82059 9008 82101 9017
rect 82059 8968 82060 9008
rect 82100 8968 82101 9008
rect 82059 8959 82101 8968
rect 81100 8924 81140 8959
rect 81100 8873 81140 8884
rect 81580 8924 81620 8933
rect 81868 8924 81908 8933
rect 81620 8884 81868 8924
rect 81580 8875 81620 8884
rect 81868 8875 81908 8884
rect 82060 8840 82100 8959
rect 82060 8791 82100 8800
rect 78412 7615 78452 7624
rect 78796 8504 78836 8513
rect 77068 7580 77108 7589
rect 76300 6656 76340 6665
rect 75820 3247 75860 3256
rect 75916 5480 75956 5489
rect 73804 2911 73844 2920
rect 75916 2624 75956 5440
rect 76108 5312 76148 5321
rect 76011 4976 76053 4985
rect 76011 4936 76012 4976
rect 76052 4936 76053 4976
rect 76011 4927 76053 4936
rect 76012 4842 76052 4927
rect 75916 2575 75956 2584
rect 76108 2540 76148 5272
rect 76300 3464 76340 6616
rect 76876 6236 76916 6245
rect 76876 5741 76916 6196
rect 76588 5732 76628 5741
rect 76588 3632 76628 5692
rect 76875 5732 76917 5741
rect 76875 5692 76876 5732
rect 76916 5692 76917 5732
rect 76875 5683 76917 5692
rect 76684 5144 76724 5155
rect 76684 5069 76724 5104
rect 76683 5060 76725 5069
rect 76683 5020 76684 5060
rect 76724 5020 76725 5060
rect 76683 5011 76725 5020
rect 76780 4985 76820 5070
rect 76779 4976 76821 4985
rect 76779 4936 76780 4976
rect 76820 4936 76821 4976
rect 76779 4927 76821 4936
rect 76588 3583 76628 3592
rect 76780 4724 76820 4733
rect 76300 3415 76340 3424
rect 76780 3464 76820 4684
rect 77068 3800 77108 7540
rect 77548 6656 77588 6665
rect 77260 4892 77300 4901
rect 77260 4472 77300 4852
rect 77260 4052 77300 4432
rect 77548 4892 77588 6616
rect 77836 6320 77876 6329
rect 77836 5741 77876 6280
rect 77835 5732 77877 5741
rect 77835 5692 77836 5732
rect 77876 5692 77877 5732
rect 77835 5683 77877 5692
rect 77836 5480 77876 5683
rect 77836 5431 77876 5440
rect 77548 4220 77588 4852
rect 77548 4171 77588 4180
rect 77260 4003 77300 4012
rect 77068 3751 77108 3760
rect 76780 3415 76820 3424
rect 78796 3212 78836 8464
rect 79288 8336 79656 8345
rect 79328 8296 79370 8336
rect 79410 8296 79452 8336
rect 79492 8296 79534 8336
rect 79574 8296 79616 8336
rect 79288 8287 79656 8296
rect 81675 8252 81717 8261
rect 81675 8212 81676 8252
rect 81716 8212 81717 8252
rect 81675 8203 81717 8212
rect 81676 8084 81716 8203
rect 81676 8035 81716 8044
rect 80528 7580 80896 7589
rect 80568 7540 80610 7580
rect 80650 7540 80692 7580
rect 80732 7540 80774 7580
rect 80814 7540 80856 7580
rect 80528 7531 80896 7540
rect 78891 7412 78933 7421
rect 78891 7372 78892 7412
rect 78932 7372 78933 7412
rect 78891 7363 78933 7372
rect 78892 7278 78932 7363
rect 81868 7244 81908 7253
rect 79288 6824 79656 6833
rect 79328 6784 79370 6824
rect 79410 6784 79452 6824
rect 79492 6784 79534 6824
rect 79574 6784 79616 6824
rect 79288 6775 79656 6784
rect 80428 6656 80468 6665
rect 79852 6572 79892 6581
rect 79755 5480 79797 5489
rect 79755 5440 79756 5480
rect 79796 5440 79797 5480
rect 79755 5431 79797 5440
rect 79756 5346 79796 5431
rect 79288 5312 79656 5321
rect 79328 5272 79370 5312
rect 79410 5272 79452 5312
rect 79492 5272 79534 5312
rect 79574 5272 79616 5312
rect 79288 5263 79656 5272
rect 79756 4136 79796 4145
rect 79288 3800 79656 3809
rect 79328 3760 79370 3800
rect 79410 3760 79452 3800
rect 79492 3760 79534 3800
rect 79574 3760 79616 3800
rect 79288 3751 79656 3760
rect 79756 3800 79796 4096
rect 79756 3751 79796 3760
rect 78796 3163 78836 3172
rect 76108 2491 76148 2500
rect 71788 1315 71828 1324
rect 35692 1147 35732 1156
rect 20716 811 20756 820
rect 79852 188 79892 6532
rect 79948 6320 79988 6329
rect 79948 1280 79988 6280
rect 80140 5564 80180 5573
rect 80140 3464 80180 5524
rect 80428 4556 80468 6616
rect 80528 6068 80896 6077
rect 80568 6028 80610 6068
rect 80650 6028 80692 6068
rect 80732 6028 80774 6068
rect 80814 6028 80856 6068
rect 80528 6019 80896 6028
rect 81676 5984 81716 5993
rect 81868 5984 81908 7204
rect 81963 6488 82005 6497
rect 81963 6448 81964 6488
rect 82004 6448 82005 6488
rect 81963 6439 82005 6448
rect 82252 6488 82292 9052
rect 83692 8672 83732 8681
rect 83692 8252 83732 8632
rect 82923 7580 82965 7589
rect 82923 7540 82924 7580
rect 82964 7540 82965 7580
rect 82923 7531 82965 7540
rect 82924 7446 82964 7531
rect 83692 7244 83732 8212
rect 83788 8420 83828 8429
rect 83788 7664 83828 8380
rect 85611 8252 85653 8261
rect 85611 8212 85612 8252
rect 85652 8212 85653 8252
rect 85611 8203 85653 8212
rect 85612 7916 85652 8203
rect 85612 7867 85652 7876
rect 83788 7615 83828 7624
rect 86859 7580 86901 7589
rect 86859 7540 86860 7580
rect 86900 7540 86901 7580
rect 86859 7531 86901 7540
rect 88396 7580 88436 7589
rect 83692 7195 83732 7204
rect 84268 6656 84308 6665
rect 82252 6439 82292 6448
rect 82348 6572 82388 6581
rect 81964 6354 82004 6439
rect 82348 6413 82388 6532
rect 82156 6404 82196 6413
rect 81716 5944 81908 5984
rect 81676 5935 81716 5944
rect 81868 5732 81908 5944
rect 81868 5683 81908 5692
rect 81772 5648 81812 5657
rect 80620 5480 80660 5489
rect 80620 4985 80660 5440
rect 81484 5396 81524 5405
rect 80619 4976 80661 4985
rect 80619 4936 80620 4976
rect 80660 4936 80661 4976
rect 80619 4927 80661 4936
rect 81292 4724 81332 4733
rect 80428 4507 80468 4516
rect 80528 4556 80896 4565
rect 80568 4516 80610 4556
rect 80650 4516 80692 4556
rect 80732 4516 80774 4556
rect 80814 4516 80856 4556
rect 80528 4507 80896 4516
rect 80140 3415 80180 3424
rect 80620 3716 80660 3725
rect 80620 3389 80660 3676
rect 80619 3380 80661 3389
rect 80619 3340 80620 3380
rect 80660 3340 80661 3380
rect 80619 3331 80661 3340
rect 80528 3044 80896 3053
rect 80568 3004 80610 3044
rect 80650 3004 80692 3044
rect 80732 3004 80774 3044
rect 80814 3004 80856 3044
rect 80528 2995 80896 3004
rect 81292 3044 81332 4684
rect 81484 3800 81524 5356
rect 81484 3751 81524 3760
rect 81676 5312 81716 5321
rect 81676 3128 81716 5272
rect 81772 4388 81812 5608
rect 82156 5648 82196 6364
rect 82347 6404 82389 6413
rect 82347 6364 82348 6404
rect 82388 6364 82389 6404
rect 82347 6355 82389 6364
rect 82827 6320 82869 6329
rect 82827 6280 82828 6320
rect 82868 6280 82869 6320
rect 82827 6271 82869 6280
rect 83788 6320 83828 6329
rect 83828 6280 83924 6320
rect 83788 6271 83828 6280
rect 82828 6186 82868 6271
rect 82156 5599 82196 5608
rect 82540 5984 82580 5993
rect 81868 5480 81908 5489
rect 81868 4901 81908 5440
rect 82540 5069 82580 5944
rect 83884 5900 83924 6280
rect 83884 5851 83924 5860
rect 82539 5060 82581 5069
rect 82539 5020 82540 5060
rect 82580 5020 82581 5060
rect 82539 5011 82581 5020
rect 81867 4892 81909 4901
rect 81867 4852 81868 4892
rect 81908 4852 81909 4892
rect 81867 4843 81909 4852
rect 81772 4339 81812 4348
rect 84268 3968 84308 6616
rect 84364 5732 84404 5743
rect 84364 5657 84404 5692
rect 84363 5648 84405 5657
rect 84363 5608 84364 5648
rect 84404 5608 84405 5648
rect 84363 5599 84405 5608
rect 85611 5060 85653 5069
rect 85611 5020 85612 5060
rect 85652 5020 85653 5060
rect 85611 5011 85653 5020
rect 85612 4808 85652 5011
rect 85612 4759 85652 4768
rect 85804 4892 85844 4901
rect 84268 3919 84308 3928
rect 81676 3079 81716 3088
rect 81868 3632 81908 3641
rect 81292 2995 81332 3004
rect 81868 2876 81908 3592
rect 81868 2827 81908 2836
rect 85708 3380 85748 3389
rect 79948 1231 79988 1240
rect 85708 860 85748 3340
rect 85804 1280 85844 4852
rect 85900 4388 85940 4397
rect 85900 2456 85940 4348
rect 86283 4136 86325 4145
rect 86283 4096 86284 4136
rect 86324 4096 86325 4136
rect 86283 4087 86325 4096
rect 86284 4002 86324 4087
rect 86860 3884 86900 7531
rect 88204 7496 88244 7505
rect 88204 7328 88244 7456
rect 88204 7076 88244 7288
rect 88204 7027 88244 7036
rect 88396 5732 88436 7540
rect 88588 7580 88628 10060
rect 94408 9848 94776 9857
rect 94448 9808 94490 9848
rect 94530 9808 94572 9848
rect 94612 9808 94654 9848
rect 94694 9808 94736 9848
rect 94408 9799 94776 9808
rect 89356 9092 89396 9101
rect 88876 8840 88916 8849
rect 88588 7531 88628 7540
rect 88684 8168 88724 8177
rect 88684 7496 88724 8128
rect 88876 7748 88916 8800
rect 88876 7699 88916 7708
rect 89260 8168 89300 8177
rect 88684 7447 88724 7456
rect 88396 5683 88436 5692
rect 86860 3835 86900 3844
rect 87052 4976 87092 4985
rect 86092 3380 86132 3389
rect 85900 2407 85940 2416
rect 85996 2624 86036 2633
rect 85804 1231 85844 1240
rect 85996 1196 86036 2584
rect 85996 1147 86036 1156
rect 85708 811 85748 820
rect 86092 272 86132 3340
rect 87052 3212 87092 4936
rect 87724 4976 87764 4985
rect 87724 4313 87764 4936
rect 88492 4976 88532 4985
rect 88492 4817 88532 4936
rect 88491 4808 88533 4817
rect 88491 4768 88492 4808
rect 88532 4768 88533 4808
rect 88491 4759 88533 4768
rect 88971 4724 89013 4733
rect 88971 4684 88972 4724
rect 89012 4684 89013 4724
rect 88971 4675 89013 4684
rect 88972 4590 89012 4675
rect 87723 4304 87765 4313
rect 87723 4264 87724 4304
rect 87764 4264 87765 4304
rect 87723 4255 87765 4264
rect 89260 3464 89300 8128
rect 89356 7580 89396 9052
rect 95648 9092 96016 9101
rect 95688 9052 95730 9092
rect 95770 9052 95812 9092
rect 95852 9052 95894 9092
rect 95934 9052 95976 9092
rect 95648 9043 96016 9052
rect 94408 8336 94776 8345
rect 94448 8296 94490 8336
rect 94530 8296 94572 8336
rect 94612 8296 94654 8336
rect 94694 8296 94736 8336
rect 94408 8287 94776 8296
rect 89356 7531 89396 7540
rect 95648 7580 96016 7589
rect 95688 7540 95730 7580
rect 95770 7540 95812 7580
rect 95852 7540 95894 7580
rect 95934 7540 95976 7580
rect 95648 7531 96016 7540
rect 94408 6824 94776 6833
rect 94448 6784 94490 6824
rect 94530 6784 94572 6824
rect 94612 6784 94654 6824
rect 94694 6784 94736 6824
rect 94408 6775 94776 6784
rect 97995 6404 98037 6413
rect 97995 6364 97996 6404
rect 98036 6364 98037 6404
rect 97995 6355 98037 6364
rect 97803 6320 97845 6329
rect 97803 6280 97804 6320
rect 97844 6280 97845 6320
rect 97803 6271 97845 6280
rect 95648 6068 96016 6077
rect 95688 6028 95730 6068
rect 95770 6028 95812 6068
rect 95852 6028 95894 6068
rect 95934 6028 95976 6068
rect 95648 6019 96016 6028
rect 97515 5648 97557 5657
rect 97515 5608 97516 5648
rect 97556 5608 97557 5648
rect 97515 5599 97557 5608
rect 97516 5514 97556 5599
rect 94408 5312 94776 5321
rect 94448 5272 94490 5312
rect 94530 5272 94572 5312
rect 94612 5272 94654 5312
rect 94694 5272 94736 5312
rect 94408 5263 94776 5272
rect 97707 4976 97749 4985
rect 97707 4936 97708 4976
rect 97748 4936 97749 4976
rect 97707 4927 97749 4936
rect 97708 4842 97748 4927
rect 95648 4556 96016 4565
rect 95688 4516 95730 4556
rect 95770 4516 95812 4556
rect 95852 4516 95894 4556
rect 95934 4516 95976 4556
rect 95648 4507 96016 4516
rect 94408 3800 94776 3809
rect 94448 3760 94490 3800
rect 94530 3760 94572 3800
rect 94612 3760 94654 3800
rect 94694 3760 94736 3800
rect 94408 3751 94776 3760
rect 95883 3632 95925 3641
rect 95883 3592 95884 3632
rect 95924 3592 95925 3632
rect 95883 3583 95925 3592
rect 89260 3415 89300 3424
rect 94732 3464 94772 3473
rect 91947 3380 91989 3389
rect 91947 3340 91948 3380
rect 91988 3340 92084 3380
rect 91947 3331 91989 3340
rect 92044 3221 92084 3340
rect 94732 3305 94772 3424
rect 95116 3464 95156 3473
rect 94731 3296 94773 3305
rect 94731 3256 94732 3296
rect 94772 3256 94773 3296
rect 94731 3247 94773 3256
rect 87052 3163 87092 3172
rect 92043 3212 92085 3221
rect 92043 3172 92044 3212
rect 92084 3172 92085 3212
rect 92043 3163 92085 3172
rect 95116 3137 95156 3424
rect 95499 3464 95541 3473
rect 95499 3424 95500 3464
rect 95540 3424 95541 3464
rect 95499 3415 95541 3424
rect 95884 3464 95924 3583
rect 95884 3415 95924 3424
rect 96651 3464 96693 3473
rect 96651 3424 96652 3464
rect 96692 3424 96693 3464
rect 96651 3415 96693 3424
rect 97420 3464 97460 3473
rect 95500 3330 95540 3415
rect 96652 3330 96692 3415
rect 97420 3221 97460 3424
rect 97804 3464 97844 6271
rect 97804 3415 97844 3424
rect 97996 3464 98036 6355
rect 98091 4976 98133 4985
rect 98091 4936 98092 4976
rect 98132 4936 98133 4976
rect 98091 4927 98133 4936
rect 98092 4842 98132 4927
rect 97996 3415 98036 3424
rect 97419 3212 97461 3221
rect 97419 3172 97420 3212
rect 97460 3172 97461 3212
rect 97419 3163 97461 3172
rect 95115 3128 95157 3137
rect 95115 3088 95116 3128
rect 95156 3088 95157 3128
rect 95115 3079 95157 3088
rect 95648 3044 96016 3053
rect 95688 3004 95730 3044
rect 95770 3004 95812 3044
rect 95852 3004 95894 3044
rect 95934 3004 95976 3044
rect 95648 2995 96016 3004
rect 87628 2540 87668 2549
rect 86188 2456 86228 2465
rect 86188 1952 86228 2416
rect 87628 2372 87668 2500
rect 87628 2323 87668 2332
rect 86188 1903 86228 1912
rect 86092 223 86132 232
rect 79852 139 79892 148
<< via4 >>
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 33928 11320 33968 11360
rect 34010 11320 34050 11360
rect 34092 11320 34132 11360
rect 34174 11320 34214 11360
rect 34256 11320 34296 11360
rect 49048 11320 49088 11360
rect 49130 11320 49170 11360
rect 49212 11320 49252 11360
rect 49294 11320 49334 11360
rect 49376 11320 49416 11360
rect 64168 11320 64208 11360
rect 64250 11320 64290 11360
rect 64332 11320 64372 11360
rect 64414 11320 64454 11360
rect 64496 11320 64536 11360
rect 79288 11320 79328 11360
rect 79370 11320 79410 11360
rect 79452 11320 79492 11360
rect 79534 11320 79574 11360
rect 79616 11320 79656 11360
rect 94408 11320 94448 11360
rect 94490 11320 94530 11360
rect 94572 11320 94612 11360
rect 94654 11320 94694 11360
rect 94736 11320 94776 11360
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 9004 9976 9044 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 7084 8128 7124 8168
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 6220 6280 6260 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 1708 5608 1748 5648
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 2092 4936 2132 4976
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 2476 4432 2516 4472
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1612 3424 1652 3464
rect 1996 3424 2036 3464
rect 2380 3424 2420 3464
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 17452 9388 17492 9428
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 16204 8128 16244 8168
rect 6988 3592 7028 3632
rect 1228 3256 1268 3296
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 17356 4264 17396 4304
rect 16396 3340 16436 3380
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19180 5860 19220 5900
rect 17548 4852 17588 4892
rect 18508 4684 18548 4724
rect 18508 3424 18548 3464
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19756 6280 19796 6320
rect 19564 4180 19604 4220
rect 19756 3508 19796 3548
rect 32044 9976 32084 10016
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 19948 4180 19988 4220
rect 20236 4180 20276 4220
rect 20140 3676 20180 3716
rect 19948 3256 19988 3296
rect 21388 5020 21428 5060
rect 21292 4768 21332 4808
rect 21292 4180 21332 4220
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 22924 7204 22964 7244
rect 23308 7204 23348 7244
rect 22924 6448 22964 6488
rect 23020 5860 23060 5900
rect 22732 4264 22772 4304
rect 22348 3592 22388 3632
rect 23788 4096 23828 4136
rect 24364 4852 24404 4892
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 24652 6532 24692 6572
rect 24652 5020 24692 5060
rect 25516 4768 25556 4808
rect 25036 4684 25076 4724
rect 26956 5860 26996 5900
rect 27628 4852 27668 4892
rect 27628 4096 27668 4136
rect 25420 3424 25460 3464
rect 30124 7204 30164 7244
rect 30124 6364 30164 6404
rect 30028 6280 30068 6320
rect 28588 4180 28628 4220
rect 29932 4096 29972 4136
rect 29068 3928 29108 3968
rect 31276 7792 31316 7832
rect 30892 5608 30932 5648
rect 31852 5776 31892 5816
rect 32428 7960 32468 8000
rect 32044 7792 32084 7832
rect 32716 5524 32756 5564
rect 32716 4684 32756 4724
rect 33196 7876 33236 7916
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33100 5860 33140 5900
rect 34252 5692 34292 5732
rect 33484 3676 33524 3716
rect 33004 3508 33044 3548
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 34252 4936 34292 4976
rect 34060 4096 34100 4136
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 34540 4096 34580 4136
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 34924 5860 34964 5900
rect 34828 4852 34868 4892
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35020 4348 35060 4388
rect 34924 4096 34964 4136
rect 37900 10060 37940 10100
rect 48364 10060 48404 10100
rect 36172 7036 36212 7076
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35788 6448 35828 6488
rect 36844 6448 36884 6488
rect 36460 6280 36500 6320
rect 35788 4684 35828 4724
rect 36652 5776 36692 5816
rect 36556 5440 36596 5480
rect 37516 6952 37556 6992
rect 37900 6532 37940 6572
rect 37708 6364 37748 6404
rect 36652 4096 36692 4136
rect 37708 3424 37748 3464
rect 45580 8044 45620 8084
rect 42604 7960 42644 8000
rect 45292 7960 45332 8000
rect 42124 7876 42164 7916
rect 41452 7708 41492 7748
rect 40108 7204 40148 7244
rect 39916 5860 39956 5900
rect 40300 5692 40340 5732
rect 39724 4852 39764 4892
rect 38668 3760 38708 3800
rect 40300 3760 40340 3800
rect 41644 6952 41684 6992
rect 41548 6280 41588 6320
rect 41740 5440 41780 5480
rect 44044 7876 44084 7916
rect 43372 7792 43412 7832
rect 42988 4096 43028 4136
rect 44332 7624 44372 7664
rect 46924 7708 46964 7748
rect 46348 7036 46388 7076
rect 45676 6532 45716 6572
rect 46348 5860 46388 5900
rect 43660 5608 43700 5648
rect 44236 4852 44276 4892
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 49996 9388 50036 9428
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 48940 6196 48980 6236
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 51820 7204 51860 7244
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 52204 5356 52244 5396
rect 49132 4180 49172 4220
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 49516 3508 49556 3548
rect 43372 3424 43412 3464
rect 47980 3424 48020 3464
rect 49228 3256 49268 3296
rect 49708 3928 49748 3968
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 50380 4348 50420 4388
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 55468 6364 55508 6404
rect 55372 6280 55412 6320
rect 55372 6112 55412 6152
rect 55468 6112 55508 6152
rect 56620 5524 56660 5564
rect 57004 6280 57044 6320
rect 57580 6280 57620 6320
rect 57964 4180 58004 4220
rect 58252 3928 58292 3968
rect 65408 10564 65448 10604
rect 65490 10564 65530 10604
rect 65572 10564 65612 10604
rect 65654 10564 65694 10604
rect 65736 10564 65776 10604
rect 80528 10564 80568 10604
rect 80610 10564 80650 10604
rect 80692 10564 80732 10604
rect 80774 10564 80814 10604
rect 80856 10564 80896 10604
rect 95648 10564 95688 10604
rect 95730 10564 95770 10604
rect 95812 10564 95852 10604
rect 95894 10564 95934 10604
rect 95976 10564 96016 10604
rect 60076 6364 60116 6404
rect 58060 3256 58100 3296
rect 60268 3256 60308 3296
rect 59500 3172 59540 3212
rect 64168 9808 64208 9848
rect 64250 9808 64290 9848
rect 64332 9808 64372 9848
rect 64414 9808 64454 9848
rect 64496 9808 64536 9848
rect 65408 9052 65448 9092
rect 65490 9052 65530 9092
rect 65572 9052 65612 9092
rect 65654 9052 65694 9092
rect 65736 9052 65776 9092
rect 64168 8296 64208 8336
rect 64250 8296 64290 8336
rect 64332 8296 64372 8336
rect 64414 8296 64454 8336
rect 64496 8296 64536 8336
rect 62668 8044 62708 8084
rect 67468 8716 67508 8756
rect 66988 7960 67028 8000
rect 66700 7792 66740 7832
rect 64492 7708 64532 7748
rect 60748 6532 60788 6572
rect 61228 5692 61268 5732
rect 60460 5524 60500 5564
rect 61804 4348 61844 4388
rect 60460 3508 60500 3548
rect 60748 3424 60788 3464
rect 63052 5860 63092 5900
rect 65408 7540 65448 7580
rect 65490 7540 65530 7580
rect 65572 7540 65612 7580
rect 65654 7540 65694 7580
rect 65736 7540 65776 7580
rect 64168 6784 64208 6824
rect 64250 6784 64290 6824
rect 64332 6784 64372 6824
rect 64414 6784 64454 6824
rect 64496 6784 64536 6824
rect 66988 6532 67028 6572
rect 67180 6448 67220 6488
rect 66796 6196 66836 6236
rect 65408 6028 65448 6068
rect 65490 6028 65530 6068
rect 65572 6028 65612 6068
rect 65654 6028 65694 6068
rect 65736 6028 65776 6068
rect 64588 5440 64628 5480
rect 64168 5272 64208 5312
rect 64250 5272 64290 5312
rect 64332 5272 64372 5312
rect 64414 5272 64454 5312
rect 64496 5272 64536 5312
rect 63244 4852 63284 4892
rect 65408 4516 65448 4556
rect 65490 4516 65530 4556
rect 65572 4516 65612 4556
rect 65654 4516 65694 4556
rect 65736 4516 65776 4556
rect 65452 4264 65492 4304
rect 64780 4180 64820 4220
rect 64168 3760 64208 3800
rect 64250 3760 64290 3800
rect 64332 3760 64372 3800
rect 64414 3760 64454 3800
rect 64496 3760 64536 3800
rect 67084 4180 67124 4220
rect 67084 3592 67124 3632
rect 64780 3508 64820 3548
rect 67660 7876 67700 7916
rect 67852 5776 67892 5816
rect 67564 4600 67604 4640
rect 67948 4264 67988 4304
rect 70540 8800 70580 8840
rect 73036 8800 73076 8840
rect 69964 4600 70004 4640
rect 70540 4264 70580 4304
rect 71020 7540 71060 7580
rect 71980 6616 72020 6656
rect 71020 6532 71060 6572
rect 71308 6448 71348 6488
rect 71884 6448 71924 6488
rect 71980 5608 72020 5648
rect 65408 3004 65448 3044
rect 65490 3004 65530 3044
rect 65572 3004 65612 3044
rect 65654 3004 65694 3044
rect 65736 3004 65776 3044
rect 72076 4768 72116 4808
rect 71884 4600 71924 4640
rect 72556 4264 72596 4304
rect 72940 5440 72980 5480
rect 72844 4684 72884 4724
rect 73516 4600 73556 4640
rect 73708 4096 73748 4136
rect 75052 8716 75092 8756
rect 74860 7540 74900 7580
rect 74956 7372 74996 7412
rect 74956 6616 74996 6656
rect 74380 5776 74420 5816
rect 74476 5524 74516 5564
rect 75148 5020 75188 5060
rect 75148 4180 75188 4220
rect 79288 9808 79328 9848
rect 79370 9808 79410 9848
rect 79452 9808 79492 9848
rect 79534 9808 79574 9848
rect 79616 9808 79656 9848
rect 80528 9052 80568 9092
rect 80610 9052 80650 9092
rect 80692 9052 80732 9092
rect 80774 9052 80814 9092
rect 80856 9052 80896 9092
rect 81100 8968 81140 9008
rect 82060 8968 82100 9008
rect 76012 4936 76052 4976
rect 76876 5692 76916 5732
rect 76684 5020 76724 5060
rect 76780 4936 76820 4976
rect 77836 5692 77876 5732
rect 79288 8296 79328 8336
rect 79370 8296 79410 8336
rect 79452 8296 79492 8336
rect 79534 8296 79574 8336
rect 79616 8296 79656 8336
rect 81676 8212 81716 8252
rect 80528 7540 80568 7580
rect 80610 7540 80650 7580
rect 80692 7540 80732 7580
rect 80774 7540 80814 7580
rect 80856 7540 80896 7580
rect 78892 7372 78932 7412
rect 79288 6784 79328 6824
rect 79370 6784 79410 6824
rect 79452 6784 79492 6824
rect 79534 6784 79574 6824
rect 79616 6784 79656 6824
rect 79756 5440 79796 5480
rect 79288 5272 79328 5312
rect 79370 5272 79410 5312
rect 79452 5272 79492 5312
rect 79534 5272 79574 5312
rect 79616 5272 79656 5312
rect 79288 3760 79328 3800
rect 79370 3760 79410 3800
rect 79452 3760 79492 3800
rect 79534 3760 79574 3800
rect 79616 3760 79656 3800
rect 80528 6028 80568 6068
rect 80610 6028 80650 6068
rect 80692 6028 80732 6068
rect 80774 6028 80814 6068
rect 80856 6028 80896 6068
rect 81964 6448 82004 6488
rect 82924 7540 82964 7580
rect 85612 8212 85652 8252
rect 86860 7540 86900 7580
rect 80620 4936 80660 4976
rect 80528 4516 80568 4556
rect 80610 4516 80650 4556
rect 80692 4516 80732 4556
rect 80774 4516 80814 4556
rect 80856 4516 80896 4556
rect 80620 3340 80660 3380
rect 80528 3004 80568 3044
rect 80610 3004 80650 3044
rect 80692 3004 80732 3044
rect 80774 3004 80814 3044
rect 80856 3004 80896 3044
rect 82348 6364 82388 6404
rect 82828 6280 82868 6320
rect 82540 5020 82580 5060
rect 81868 4852 81908 4892
rect 84364 5608 84404 5648
rect 85612 5020 85652 5060
rect 86284 4096 86324 4136
rect 94408 9808 94448 9848
rect 94490 9808 94530 9848
rect 94572 9808 94612 9848
rect 94654 9808 94694 9848
rect 94736 9808 94776 9848
rect 88492 4768 88532 4808
rect 88972 4684 89012 4724
rect 87724 4264 87764 4304
rect 95648 9052 95688 9092
rect 95730 9052 95770 9092
rect 95812 9052 95852 9092
rect 95894 9052 95934 9092
rect 95976 9052 96016 9092
rect 94408 8296 94448 8336
rect 94490 8296 94530 8336
rect 94572 8296 94612 8336
rect 94654 8296 94694 8336
rect 94736 8296 94776 8336
rect 95648 7540 95688 7580
rect 95730 7540 95770 7580
rect 95812 7540 95852 7580
rect 95894 7540 95934 7580
rect 95976 7540 96016 7580
rect 94408 6784 94448 6824
rect 94490 6784 94530 6824
rect 94572 6784 94612 6824
rect 94654 6784 94694 6824
rect 94736 6784 94776 6824
rect 97996 6364 98036 6404
rect 97804 6280 97844 6320
rect 95648 6028 95688 6068
rect 95730 6028 95770 6068
rect 95812 6028 95852 6068
rect 95894 6028 95934 6068
rect 95976 6028 96016 6068
rect 97516 5608 97556 5648
rect 94408 5272 94448 5312
rect 94490 5272 94530 5312
rect 94572 5272 94612 5312
rect 94654 5272 94694 5312
rect 94736 5272 94776 5312
rect 97708 4936 97748 4976
rect 95648 4516 95688 4556
rect 95730 4516 95770 4556
rect 95812 4516 95852 4556
rect 95894 4516 95934 4556
rect 95976 4516 96016 4556
rect 94408 3760 94448 3800
rect 94490 3760 94530 3800
rect 94572 3760 94612 3800
rect 94654 3760 94694 3800
rect 94736 3760 94776 3800
rect 95884 3592 95924 3632
rect 91948 3340 91988 3380
rect 94732 3256 94772 3296
rect 92044 3172 92084 3212
rect 95500 3424 95540 3464
rect 96652 3424 96692 3464
rect 98092 4936 98132 4976
rect 97420 3172 97460 3212
rect 95116 3088 95156 3128
rect 95648 3004 95688 3044
rect 95730 3004 95770 3044
rect 95812 3004 95852 3044
rect 95894 3004 95934 3044
rect 95976 3004 96016 3044
<< metal5 >>
rect 3679 11383 4065 11402
rect 3679 11360 3745 11383
rect 3831 11360 3913 11383
rect 3999 11360 4065 11383
rect 3679 11320 3688 11360
rect 3728 11320 3745 11360
rect 3831 11320 3852 11360
rect 3892 11320 3913 11360
rect 3999 11320 4016 11360
rect 4056 11320 4065 11360
rect 3679 11297 3745 11320
rect 3831 11297 3913 11320
rect 3999 11297 4065 11320
rect 3679 11278 4065 11297
rect 18799 11383 19185 11402
rect 18799 11360 18865 11383
rect 18951 11360 19033 11383
rect 19119 11360 19185 11383
rect 18799 11320 18808 11360
rect 18848 11320 18865 11360
rect 18951 11320 18972 11360
rect 19012 11320 19033 11360
rect 19119 11320 19136 11360
rect 19176 11320 19185 11360
rect 18799 11297 18865 11320
rect 18951 11297 19033 11320
rect 19119 11297 19185 11320
rect 18799 11278 19185 11297
rect 33919 11383 34305 11402
rect 33919 11360 33985 11383
rect 34071 11360 34153 11383
rect 34239 11360 34305 11383
rect 33919 11320 33928 11360
rect 33968 11320 33985 11360
rect 34071 11320 34092 11360
rect 34132 11320 34153 11360
rect 34239 11320 34256 11360
rect 34296 11320 34305 11360
rect 33919 11297 33985 11320
rect 34071 11297 34153 11320
rect 34239 11297 34305 11320
rect 33919 11278 34305 11297
rect 49039 11383 49425 11402
rect 49039 11360 49105 11383
rect 49191 11360 49273 11383
rect 49359 11360 49425 11383
rect 49039 11320 49048 11360
rect 49088 11320 49105 11360
rect 49191 11320 49212 11360
rect 49252 11320 49273 11360
rect 49359 11320 49376 11360
rect 49416 11320 49425 11360
rect 49039 11297 49105 11320
rect 49191 11297 49273 11320
rect 49359 11297 49425 11320
rect 49039 11278 49425 11297
rect 64159 11383 64545 11402
rect 64159 11360 64225 11383
rect 64311 11360 64393 11383
rect 64479 11360 64545 11383
rect 64159 11320 64168 11360
rect 64208 11320 64225 11360
rect 64311 11320 64332 11360
rect 64372 11320 64393 11360
rect 64479 11320 64496 11360
rect 64536 11320 64545 11360
rect 64159 11297 64225 11320
rect 64311 11297 64393 11320
rect 64479 11297 64545 11320
rect 64159 11278 64545 11297
rect 79279 11383 79665 11402
rect 79279 11360 79345 11383
rect 79431 11360 79513 11383
rect 79599 11360 79665 11383
rect 79279 11320 79288 11360
rect 79328 11320 79345 11360
rect 79431 11320 79452 11360
rect 79492 11320 79513 11360
rect 79599 11320 79616 11360
rect 79656 11320 79665 11360
rect 79279 11297 79345 11320
rect 79431 11297 79513 11320
rect 79599 11297 79665 11320
rect 79279 11278 79665 11297
rect 94399 11383 94785 11402
rect 94399 11360 94465 11383
rect 94551 11360 94633 11383
rect 94719 11360 94785 11383
rect 94399 11320 94408 11360
rect 94448 11320 94465 11360
rect 94551 11320 94572 11360
rect 94612 11320 94633 11360
rect 94719 11320 94736 11360
rect 94776 11320 94785 11360
rect 94399 11297 94465 11320
rect 94551 11297 94633 11320
rect 94719 11297 94785 11320
rect 94399 11278 94785 11297
rect 4919 10627 5305 10646
rect 4919 10604 4985 10627
rect 5071 10604 5153 10627
rect 5239 10604 5305 10627
rect 4919 10564 4928 10604
rect 4968 10564 4985 10604
rect 5071 10564 5092 10604
rect 5132 10564 5153 10604
rect 5239 10564 5256 10604
rect 5296 10564 5305 10604
rect 4919 10541 4985 10564
rect 5071 10541 5153 10564
rect 5239 10541 5305 10564
rect 4919 10522 5305 10541
rect 20039 10627 20425 10646
rect 20039 10604 20105 10627
rect 20191 10604 20273 10627
rect 20359 10604 20425 10627
rect 20039 10564 20048 10604
rect 20088 10564 20105 10604
rect 20191 10564 20212 10604
rect 20252 10564 20273 10604
rect 20359 10564 20376 10604
rect 20416 10564 20425 10604
rect 20039 10541 20105 10564
rect 20191 10541 20273 10564
rect 20359 10541 20425 10564
rect 20039 10522 20425 10541
rect 35159 10627 35545 10646
rect 35159 10604 35225 10627
rect 35311 10604 35393 10627
rect 35479 10604 35545 10627
rect 35159 10564 35168 10604
rect 35208 10564 35225 10604
rect 35311 10564 35332 10604
rect 35372 10564 35393 10604
rect 35479 10564 35496 10604
rect 35536 10564 35545 10604
rect 35159 10541 35225 10564
rect 35311 10541 35393 10564
rect 35479 10541 35545 10564
rect 35159 10522 35545 10541
rect 50279 10627 50665 10646
rect 50279 10604 50345 10627
rect 50431 10604 50513 10627
rect 50599 10604 50665 10627
rect 50279 10564 50288 10604
rect 50328 10564 50345 10604
rect 50431 10564 50452 10604
rect 50492 10564 50513 10604
rect 50599 10564 50616 10604
rect 50656 10564 50665 10604
rect 50279 10541 50345 10564
rect 50431 10541 50513 10564
rect 50599 10541 50665 10564
rect 50279 10522 50665 10541
rect 65399 10627 65785 10646
rect 65399 10604 65465 10627
rect 65551 10604 65633 10627
rect 65719 10604 65785 10627
rect 65399 10564 65408 10604
rect 65448 10564 65465 10604
rect 65551 10564 65572 10604
rect 65612 10564 65633 10604
rect 65719 10564 65736 10604
rect 65776 10564 65785 10604
rect 65399 10541 65465 10564
rect 65551 10541 65633 10564
rect 65719 10541 65785 10564
rect 65399 10522 65785 10541
rect 80519 10627 80905 10646
rect 80519 10604 80585 10627
rect 80671 10604 80753 10627
rect 80839 10604 80905 10627
rect 80519 10564 80528 10604
rect 80568 10564 80585 10604
rect 80671 10564 80692 10604
rect 80732 10564 80753 10604
rect 80839 10564 80856 10604
rect 80896 10564 80905 10604
rect 80519 10541 80585 10564
rect 80671 10541 80753 10564
rect 80839 10541 80905 10564
rect 80519 10522 80905 10541
rect 95639 10627 96025 10646
rect 95639 10604 95705 10627
rect 95791 10604 95873 10627
rect 95959 10604 96025 10627
rect 95639 10564 95648 10604
rect 95688 10564 95705 10604
rect 95791 10564 95812 10604
rect 95852 10564 95873 10604
rect 95959 10564 95976 10604
rect 96016 10564 96025 10604
rect 95639 10541 95705 10564
rect 95791 10541 95873 10564
rect 95959 10541 96025 10564
rect 95639 10522 96025 10541
rect 37891 10060 37900 10100
rect 37940 10060 48364 10100
rect 48404 10060 48413 10100
rect 8995 9976 9004 10016
rect 9044 9976 32044 10016
rect 32084 9976 32093 10016
rect 3679 9871 4065 9890
rect 3679 9848 3745 9871
rect 3831 9848 3913 9871
rect 3999 9848 4065 9871
rect 3679 9808 3688 9848
rect 3728 9808 3745 9848
rect 3831 9808 3852 9848
rect 3892 9808 3913 9848
rect 3999 9808 4016 9848
rect 4056 9808 4065 9848
rect 3679 9785 3745 9808
rect 3831 9785 3913 9808
rect 3999 9785 4065 9808
rect 3679 9766 4065 9785
rect 18799 9871 19185 9890
rect 18799 9848 18865 9871
rect 18951 9848 19033 9871
rect 19119 9848 19185 9871
rect 18799 9808 18808 9848
rect 18848 9808 18865 9848
rect 18951 9808 18972 9848
rect 19012 9808 19033 9848
rect 19119 9808 19136 9848
rect 19176 9808 19185 9848
rect 18799 9785 18865 9808
rect 18951 9785 19033 9808
rect 19119 9785 19185 9808
rect 18799 9766 19185 9785
rect 33919 9871 34305 9890
rect 33919 9848 33985 9871
rect 34071 9848 34153 9871
rect 34239 9848 34305 9871
rect 33919 9808 33928 9848
rect 33968 9808 33985 9848
rect 34071 9808 34092 9848
rect 34132 9808 34153 9848
rect 34239 9808 34256 9848
rect 34296 9808 34305 9848
rect 33919 9785 33985 9808
rect 34071 9785 34153 9808
rect 34239 9785 34305 9808
rect 33919 9766 34305 9785
rect 49039 9871 49425 9890
rect 49039 9848 49105 9871
rect 49191 9848 49273 9871
rect 49359 9848 49425 9871
rect 49039 9808 49048 9848
rect 49088 9808 49105 9848
rect 49191 9808 49212 9848
rect 49252 9808 49273 9848
rect 49359 9808 49376 9848
rect 49416 9808 49425 9848
rect 49039 9785 49105 9808
rect 49191 9785 49273 9808
rect 49359 9785 49425 9808
rect 49039 9766 49425 9785
rect 64159 9871 64545 9890
rect 64159 9848 64225 9871
rect 64311 9848 64393 9871
rect 64479 9848 64545 9871
rect 64159 9808 64168 9848
rect 64208 9808 64225 9848
rect 64311 9808 64332 9848
rect 64372 9808 64393 9848
rect 64479 9808 64496 9848
rect 64536 9808 64545 9848
rect 64159 9785 64225 9808
rect 64311 9785 64393 9808
rect 64479 9785 64545 9808
rect 64159 9766 64545 9785
rect 79279 9871 79665 9890
rect 79279 9848 79345 9871
rect 79431 9848 79513 9871
rect 79599 9848 79665 9871
rect 79279 9808 79288 9848
rect 79328 9808 79345 9848
rect 79431 9808 79452 9848
rect 79492 9808 79513 9848
rect 79599 9808 79616 9848
rect 79656 9808 79665 9848
rect 79279 9785 79345 9808
rect 79431 9785 79513 9808
rect 79599 9785 79665 9808
rect 79279 9766 79665 9785
rect 94399 9871 94785 9890
rect 94399 9848 94465 9871
rect 94551 9848 94633 9871
rect 94719 9848 94785 9871
rect 94399 9808 94408 9848
rect 94448 9808 94465 9848
rect 94551 9808 94572 9848
rect 94612 9808 94633 9848
rect 94719 9808 94736 9848
rect 94776 9808 94785 9848
rect 94399 9785 94465 9808
rect 94551 9785 94633 9808
rect 94719 9785 94785 9808
rect 94399 9766 94785 9785
rect 17443 9388 17452 9428
rect 17492 9388 49996 9428
rect 50036 9388 50045 9428
rect 4919 9115 5305 9134
rect 4919 9092 4985 9115
rect 5071 9092 5153 9115
rect 5239 9092 5305 9115
rect 4919 9052 4928 9092
rect 4968 9052 4985 9092
rect 5071 9052 5092 9092
rect 5132 9052 5153 9092
rect 5239 9052 5256 9092
rect 5296 9052 5305 9092
rect 4919 9029 4985 9052
rect 5071 9029 5153 9052
rect 5239 9029 5305 9052
rect 4919 9010 5305 9029
rect 20039 9115 20425 9134
rect 20039 9092 20105 9115
rect 20191 9092 20273 9115
rect 20359 9092 20425 9115
rect 20039 9052 20048 9092
rect 20088 9052 20105 9092
rect 20191 9052 20212 9092
rect 20252 9052 20273 9092
rect 20359 9052 20376 9092
rect 20416 9052 20425 9092
rect 20039 9029 20105 9052
rect 20191 9029 20273 9052
rect 20359 9029 20425 9052
rect 20039 9010 20425 9029
rect 35159 9115 35545 9134
rect 35159 9092 35225 9115
rect 35311 9092 35393 9115
rect 35479 9092 35545 9115
rect 35159 9052 35168 9092
rect 35208 9052 35225 9092
rect 35311 9052 35332 9092
rect 35372 9052 35393 9092
rect 35479 9052 35496 9092
rect 35536 9052 35545 9092
rect 35159 9029 35225 9052
rect 35311 9029 35393 9052
rect 35479 9029 35545 9052
rect 35159 9010 35545 9029
rect 50279 9115 50665 9134
rect 50279 9092 50345 9115
rect 50431 9092 50513 9115
rect 50599 9092 50665 9115
rect 50279 9052 50288 9092
rect 50328 9052 50345 9092
rect 50431 9052 50452 9092
rect 50492 9052 50513 9092
rect 50599 9052 50616 9092
rect 50656 9052 50665 9092
rect 50279 9029 50345 9052
rect 50431 9029 50513 9052
rect 50599 9029 50665 9052
rect 50279 9010 50665 9029
rect 65399 9115 65785 9134
rect 65399 9092 65465 9115
rect 65551 9092 65633 9115
rect 65719 9092 65785 9115
rect 65399 9052 65408 9092
rect 65448 9052 65465 9092
rect 65551 9052 65572 9092
rect 65612 9052 65633 9092
rect 65719 9052 65736 9092
rect 65776 9052 65785 9092
rect 65399 9029 65465 9052
rect 65551 9029 65633 9052
rect 65719 9029 65785 9052
rect 65399 9010 65785 9029
rect 80519 9115 80905 9134
rect 80519 9092 80585 9115
rect 80671 9092 80753 9115
rect 80839 9092 80905 9115
rect 80519 9052 80528 9092
rect 80568 9052 80585 9092
rect 80671 9052 80692 9092
rect 80732 9052 80753 9092
rect 80839 9052 80856 9092
rect 80896 9052 80905 9092
rect 80519 9029 80585 9052
rect 80671 9029 80753 9052
rect 80839 9029 80905 9052
rect 80519 9010 80905 9029
rect 95639 9115 96025 9134
rect 95639 9092 95705 9115
rect 95791 9092 95873 9115
rect 95959 9092 96025 9115
rect 95639 9052 95648 9092
rect 95688 9052 95705 9092
rect 95791 9052 95812 9092
rect 95852 9052 95873 9092
rect 95959 9052 95976 9092
rect 96016 9052 96025 9092
rect 95639 9029 95705 9052
rect 95791 9029 95873 9052
rect 95959 9029 96025 9052
rect 95639 9010 96025 9029
rect 81091 8968 81100 9008
rect 81140 8968 82060 9008
rect 82100 8968 82109 9008
rect 70531 8800 70540 8840
rect 70580 8800 70589 8840
rect 73027 8800 73036 8840
rect 73076 8800 73085 8840
rect 70540 8756 70580 8800
rect 67459 8716 67468 8756
rect 67508 8716 70580 8756
rect 73036 8756 73076 8800
rect 73036 8716 75052 8756
rect 75092 8716 75101 8756
rect 3679 8359 4065 8378
rect 3679 8336 3745 8359
rect 3831 8336 3913 8359
rect 3999 8336 4065 8359
rect 3679 8296 3688 8336
rect 3728 8296 3745 8336
rect 3831 8296 3852 8336
rect 3892 8296 3913 8336
rect 3999 8296 4016 8336
rect 4056 8296 4065 8336
rect 3679 8273 3745 8296
rect 3831 8273 3913 8296
rect 3999 8273 4065 8296
rect 3679 8254 4065 8273
rect 18799 8359 19185 8378
rect 18799 8336 18865 8359
rect 18951 8336 19033 8359
rect 19119 8336 19185 8359
rect 18799 8296 18808 8336
rect 18848 8296 18865 8336
rect 18951 8296 18972 8336
rect 19012 8296 19033 8336
rect 19119 8296 19136 8336
rect 19176 8296 19185 8336
rect 18799 8273 18865 8296
rect 18951 8273 19033 8296
rect 19119 8273 19185 8296
rect 18799 8254 19185 8273
rect 33919 8359 34305 8378
rect 33919 8336 33985 8359
rect 34071 8336 34153 8359
rect 34239 8336 34305 8359
rect 33919 8296 33928 8336
rect 33968 8296 33985 8336
rect 34071 8296 34092 8336
rect 34132 8296 34153 8336
rect 34239 8296 34256 8336
rect 34296 8296 34305 8336
rect 33919 8273 33985 8296
rect 34071 8273 34153 8296
rect 34239 8273 34305 8296
rect 33919 8254 34305 8273
rect 49039 8359 49425 8378
rect 49039 8336 49105 8359
rect 49191 8336 49273 8359
rect 49359 8336 49425 8359
rect 49039 8296 49048 8336
rect 49088 8296 49105 8336
rect 49191 8296 49212 8336
rect 49252 8296 49273 8336
rect 49359 8296 49376 8336
rect 49416 8296 49425 8336
rect 49039 8273 49105 8296
rect 49191 8273 49273 8296
rect 49359 8273 49425 8296
rect 49039 8254 49425 8273
rect 64159 8359 64545 8378
rect 64159 8336 64225 8359
rect 64311 8336 64393 8359
rect 64479 8336 64545 8359
rect 64159 8296 64168 8336
rect 64208 8296 64225 8336
rect 64311 8296 64332 8336
rect 64372 8296 64393 8336
rect 64479 8296 64496 8336
rect 64536 8296 64545 8336
rect 64159 8273 64225 8296
rect 64311 8273 64393 8296
rect 64479 8273 64545 8296
rect 64159 8254 64545 8273
rect 79279 8359 79665 8378
rect 79279 8336 79345 8359
rect 79431 8336 79513 8359
rect 79599 8336 79665 8359
rect 79279 8296 79288 8336
rect 79328 8296 79345 8336
rect 79431 8296 79452 8336
rect 79492 8296 79513 8336
rect 79599 8296 79616 8336
rect 79656 8296 79665 8336
rect 79279 8273 79345 8296
rect 79431 8273 79513 8296
rect 79599 8273 79665 8296
rect 79279 8254 79665 8273
rect 94399 8359 94785 8378
rect 94399 8336 94465 8359
rect 94551 8336 94633 8359
rect 94719 8336 94785 8359
rect 94399 8296 94408 8336
rect 94448 8296 94465 8336
rect 94551 8296 94572 8336
rect 94612 8296 94633 8336
rect 94719 8296 94736 8336
rect 94776 8296 94785 8336
rect 94399 8273 94465 8296
rect 94551 8273 94633 8296
rect 94719 8273 94785 8296
rect 94399 8254 94785 8273
rect 81667 8212 81676 8252
rect 81716 8212 85612 8252
rect 85652 8212 85661 8252
rect 7075 8128 7084 8168
rect 7124 8128 16204 8168
rect 16244 8128 16253 8168
rect 45571 8044 45580 8084
rect 45620 8044 62668 8084
rect 62708 8044 62717 8084
rect 32419 7960 32428 8000
rect 32468 7960 42604 8000
rect 42644 7960 42653 8000
rect 45283 7960 45292 8000
rect 45332 7960 66988 8000
rect 67028 7960 67037 8000
rect 33187 7876 33196 7916
rect 33236 7876 42124 7916
rect 42164 7876 42173 7916
rect 44035 7876 44044 7916
rect 44084 7876 67660 7916
rect 67700 7876 67709 7916
rect 31267 7792 31276 7832
rect 31316 7792 31812 7832
rect 32035 7792 32044 7832
rect 32084 7792 43372 7832
rect 43412 7792 43421 7832
rect 46600 7792 66700 7832
rect 66740 7792 66749 7832
rect 31772 7748 31812 7792
rect 31772 7708 41452 7748
rect 41492 7708 41501 7748
rect 46600 7664 46640 7792
rect 46915 7708 46924 7748
rect 46964 7708 64492 7748
rect 64532 7708 64541 7748
rect 44323 7624 44332 7664
rect 44372 7624 46640 7664
rect 4919 7603 5305 7622
rect 4919 7580 4985 7603
rect 5071 7580 5153 7603
rect 5239 7580 5305 7603
rect 4919 7540 4928 7580
rect 4968 7540 4985 7580
rect 5071 7540 5092 7580
rect 5132 7540 5153 7580
rect 5239 7540 5256 7580
rect 5296 7540 5305 7580
rect 4919 7517 4985 7540
rect 5071 7517 5153 7540
rect 5239 7517 5305 7540
rect 4919 7498 5305 7517
rect 20039 7603 20425 7622
rect 20039 7580 20105 7603
rect 20191 7580 20273 7603
rect 20359 7580 20425 7603
rect 20039 7540 20048 7580
rect 20088 7540 20105 7580
rect 20191 7540 20212 7580
rect 20252 7540 20273 7580
rect 20359 7540 20376 7580
rect 20416 7540 20425 7580
rect 20039 7517 20105 7540
rect 20191 7517 20273 7540
rect 20359 7517 20425 7540
rect 20039 7498 20425 7517
rect 35159 7603 35545 7622
rect 35159 7580 35225 7603
rect 35311 7580 35393 7603
rect 35479 7580 35545 7603
rect 35159 7540 35168 7580
rect 35208 7540 35225 7580
rect 35311 7540 35332 7580
rect 35372 7540 35393 7580
rect 35479 7540 35496 7580
rect 35536 7540 35545 7580
rect 35159 7517 35225 7540
rect 35311 7517 35393 7540
rect 35479 7517 35545 7540
rect 35159 7498 35545 7517
rect 50279 7603 50665 7622
rect 50279 7580 50345 7603
rect 50431 7580 50513 7603
rect 50599 7580 50665 7603
rect 50279 7540 50288 7580
rect 50328 7540 50345 7580
rect 50431 7540 50452 7580
rect 50492 7540 50513 7580
rect 50599 7540 50616 7580
rect 50656 7540 50665 7580
rect 50279 7517 50345 7540
rect 50431 7517 50513 7540
rect 50599 7517 50665 7540
rect 50279 7498 50665 7517
rect 65399 7603 65785 7622
rect 65399 7580 65465 7603
rect 65551 7580 65633 7603
rect 65719 7580 65785 7603
rect 80519 7603 80905 7622
rect 80519 7580 80585 7603
rect 80671 7580 80753 7603
rect 80839 7580 80905 7603
rect 95639 7603 96025 7622
rect 95639 7580 95705 7603
rect 95791 7580 95873 7603
rect 95959 7580 96025 7603
rect 65399 7540 65408 7580
rect 65448 7540 65465 7580
rect 65551 7540 65572 7580
rect 65612 7540 65633 7580
rect 65719 7540 65736 7580
rect 65776 7540 65785 7580
rect 71011 7540 71020 7580
rect 71060 7540 74860 7580
rect 74900 7540 74909 7580
rect 80519 7540 80528 7580
rect 80568 7540 80585 7580
rect 80671 7540 80692 7580
rect 80732 7540 80753 7580
rect 80839 7540 80856 7580
rect 80896 7540 80905 7580
rect 82915 7540 82924 7580
rect 82964 7540 86860 7580
rect 86900 7540 86909 7580
rect 95639 7540 95648 7580
rect 95688 7540 95705 7580
rect 95791 7540 95812 7580
rect 95852 7540 95873 7580
rect 95959 7540 95976 7580
rect 96016 7540 96025 7580
rect 65399 7517 65465 7540
rect 65551 7517 65633 7540
rect 65719 7517 65785 7540
rect 65399 7498 65785 7517
rect 80519 7517 80585 7540
rect 80671 7517 80753 7540
rect 80839 7517 80905 7540
rect 80519 7498 80905 7517
rect 95639 7517 95705 7540
rect 95791 7517 95873 7540
rect 95959 7517 96025 7540
rect 95639 7498 96025 7517
rect 74947 7372 74956 7412
rect 74996 7372 78892 7412
rect 78932 7372 78941 7412
rect 22915 7204 22924 7244
rect 22964 7204 23308 7244
rect 23348 7204 30124 7244
rect 30164 7204 30173 7244
rect 40099 7204 40108 7244
rect 40148 7204 51820 7244
rect 51860 7204 51869 7244
rect 36163 7036 36172 7076
rect 36212 7036 46348 7076
rect 46388 7036 46397 7076
rect 37507 6952 37516 6992
rect 37556 6952 41644 6992
rect 41684 6952 41693 6992
rect 3679 6847 4065 6866
rect 3679 6824 3745 6847
rect 3831 6824 3913 6847
rect 3999 6824 4065 6847
rect 3679 6784 3688 6824
rect 3728 6784 3745 6824
rect 3831 6784 3852 6824
rect 3892 6784 3913 6824
rect 3999 6784 4016 6824
rect 4056 6784 4065 6824
rect 3679 6761 3745 6784
rect 3831 6761 3913 6784
rect 3999 6761 4065 6784
rect 3679 6742 4065 6761
rect 18799 6847 19185 6866
rect 18799 6824 18865 6847
rect 18951 6824 19033 6847
rect 19119 6824 19185 6847
rect 18799 6784 18808 6824
rect 18848 6784 18865 6824
rect 18951 6784 18972 6824
rect 19012 6784 19033 6824
rect 19119 6784 19136 6824
rect 19176 6784 19185 6824
rect 18799 6761 18865 6784
rect 18951 6761 19033 6784
rect 19119 6761 19185 6784
rect 18799 6742 19185 6761
rect 33919 6847 34305 6866
rect 33919 6824 33985 6847
rect 34071 6824 34153 6847
rect 34239 6824 34305 6847
rect 33919 6784 33928 6824
rect 33968 6784 33985 6824
rect 34071 6784 34092 6824
rect 34132 6784 34153 6824
rect 34239 6784 34256 6824
rect 34296 6784 34305 6824
rect 33919 6761 33985 6784
rect 34071 6761 34153 6784
rect 34239 6761 34305 6784
rect 33919 6742 34305 6761
rect 49039 6847 49425 6866
rect 49039 6824 49105 6847
rect 49191 6824 49273 6847
rect 49359 6824 49425 6847
rect 49039 6784 49048 6824
rect 49088 6784 49105 6824
rect 49191 6784 49212 6824
rect 49252 6784 49273 6824
rect 49359 6784 49376 6824
rect 49416 6784 49425 6824
rect 49039 6761 49105 6784
rect 49191 6761 49273 6784
rect 49359 6761 49425 6784
rect 49039 6742 49425 6761
rect 64159 6847 64545 6866
rect 64159 6824 64225 6847
rect 64311 6824 64393 6847
rect 64479 6824 64545 6847
rect 64159 6784 64168 6824
rect 64208 6784 64225 6824
rect 64311 6784 64332 6824
rect 64372 6784 64393 6824
rect 64479 6784 64496 6824
rect 64536 6784 64545 6824
rect 64159 6761 64225 6784
rect 64311 6761 64393 6784
rect 64479 6761 64545 6784
rect 64159 6742 64545 6761
rect 79279 6847 79665 6866
rect 79279 6824 79345 6847
rect 79431 6824 79513 6847
rect 79599 6824 79665 6847
rect 79279 6784 79288 6824
rect 79328 6784 79345 6824
rect 79431 6784 79452 6824
rect 79492 6784 79513 6824
rect 79599 6784 79616 6824
rect 79656 6784 79665 6824
rect 79279 6761 79345 6784
rect 79431 6761 79513 6784
rect 79599 6761 79665 6784
rect 79279 6742 79665 6761
rect 94399 6847 94785 6866
rect 94399 6824 94465 6847
rect 94551 6824 94633 6847
rect 94719 6824 94785 6847
rect 94399 6784 94408 6824
rect 94448 6784 94465 6824
rect 94551 6784 94572 6824
rect 94612 6784 94633 6824
rect 94719 6784 94736 6824
rect 94776 6784 94785 6824
rect 94399 6761 94465 6784
rect 94551 6761 94633 6784
rect 94719 6761 94785 6784
rect 94399 6742 94785 6761
rect 41560 6616 71980 6656
rect 72020 6616 74956 6656
rect 74996 6616 75005 6656
rect 41560 6572 41600 6616
rect 24643 6532 24652 6572
rect 24692 6532 37900 6572
rect 37940 6532 41600 6572
rect 45667 6532 45676 6572
rect 45716 6532 60748 6572
rect 60788 6532 60797 6572
rect 66979 6532 66988 6572
rect 67028 6532 71020 6572
rect 71060 6532 71069 6572
rect 22915 6448 22924 6488
rect 22964 6448 35788 6488
rect 35828 6448 36844 6488
rect 36884 6448 67180 6488
rect 67220 6448 71308 6488
rect 71348 6448 71357 6488
rect 71875 6448 71884 6488
rect 71924 6448 81964 6488
rect 82004 6448 82013 6488
rect 30115 6364 30124 6404
rect 30164 6364 37708 6404
rect 37748 6364 37757 6404
rect 55459 6364 55468 6404
rect 55508 6364 60076 6404
rect 60116 6364 60125 6404
rect 82339 6364 82348 6404
rect 82388 6364 97996 6404
rect 98036 6364 98045 6404
rect 6211 6280 6220 6320
rect 6260 6280 19756 6320
rect 19796 6280 19805 6320
rect 30019 6280 30028 6320
rect 30068 6280 36460 6320
rect 36500 6280 36509 6320
rect 41539 6280 41548 6320
rect 41588 6280 41600 6320
rect 41560 6236 41600 6280
rect 46600 6280 55372 6320
rect 55412 6280 55421 6320
rect 56995 6280 57004 6320
rect 57044 6280 57580 6320
rect 57620 6280 57629 6320
rect 82819 6280 82828 6320
rect 82868 6280 97804 6320
rect 97844 6280 97853 6320
rect 46600 6236 46640 6280
rect 41560 6196 46640 6236
rect 48931 6196 48940 6236
rect 48980 6196 66796 6236
rect 66836 6196 66845 6236
rect 55363 6112 55372 6152
rect 55412 6112 55468 6152
rect 55508 6112 55536 6152
rect 4919 6091 5305 6110
rect 4919 6068 4985 6091
rect 5071 6068 5153 6091
rect 5239 6068 5305 6091
rect 4919 6028 4928 6068
rect 4968 6028 4985 6068
rect 5071 6028 5092 6068
rect 5132 6028 5153 6068
rect 5239 6028 5256 6068
rect 5296 6028 5305 6068
rect 4919 6005 4985 6028
rect 5071 6005 5153 6028
rect 5239 6005 5305 6028
rect 4919 5986 5305 6005
rect 20039 6091 20425 6110
rect 20039 6068 20105 6091
rect 20191 6068 20273 6091
rect 20359 6068 20425 6091
rect 20039 6028 20048 6068
rect 20088 6028 20105 6068
rect 20191 6028 20212 6068
rect 20252 6028 20273 6068
rect 20359 6028 20376 6068
rect 20416 6028 20425 6068
rect 20039 6005 20105 6028
rect 20191 6005 20273 6028
rect 20359 6005 20425 6028
rect 20039 5986 20425 6005
rect 35159 6091 35545 6110
rect 35159 6068 35225 6091
rect 35311 6068 35393 6091
rect 35479 6068 35545 6091
rect 35159 6028 35168 6068
rect 35208 6028 35225 6068
rect 35311 6028 35332 6068
rect 35372 6028 35393 6068
rect 35479 6028 35496 6068
rect 35536 6028 35545 6068
rect 35159 6005 35225 6028
rect 35311 6005 35393 6028
rect 35479 6005 35545 6028
rect 35159 5986 35545 6005
rect 50279 6091 50665 6110
rect 50279 6068 50345 6091
rect 50431 6068 50513 6091
rect 50599 6068 50665 6091
rect 50279 6028 50288 6068
rect 50328 6028 50345 6068
rect 50431 6028 50452 6068
rect 50492 6028 50513 6068
rect 50599 6028 50616 6068
rect 50656 6028 50665 6068
rect 50279 6005 50345 6028
rect 50431 6005 50513 6028
rect 50599 6005 50665 6028
rect 50279 5986 50665 6005
rect 65399 6091 65785 6110
rect 65399 6068 65465 6091
rect 65551 6068 65633 6091
rect 65719 6068 65785 6091
rect 65399 6028 65408 6068
rect 65448 6028 65465 6068
rect 65551 6028 65572 6068
rect 65612 6028 65633 6068
rect 65719 6028 65736 6068
rect 65776 6028 65785 6068
rect 65399 6005 65465 6028
rect 65551 6005 65633 6028
rect 65719 6005 65785 6028
rect 65399 5986 65785 6005
rect 80519 6091 80905 6110
rect 80519 6068 80585 6091
rect 80671 6068 80753 6091
rect 80839 6068 80905 6091
rect 80519 6028 80528 6068
rect 80568 6028 80585 6068
rect 80671 6028 80692 6068
rect 80732 6028 80753 6068
rect 80839 6028 80856 6068
rect 80896 6028 80905 6068
rect 80519 6005 80585 6028
rect 80671 6005 80753 6028
rect 80839 6005 80905 6028
rect 80519 5986 80905 6005
rect 95639 6091 96025 6110
rect 95639 6068 95705 6091
rect 95791 6068 95873 6091
rect 95959 6068 96025 6091
rect 95639 6028 95648 6068
rect 95688 6028 95705 6068
rect 95791 6028 95812 6068
rect 95852 6028 95873 6068
rect 95959 6028 95976 6068
rect 96016 6028 96025 6068
rect 95639 6005 95705 6028
rect 95791 6005 95873 6028
rect 95959 6005 96025 6028
rect 95639 5986 96025 6005
rect 19171 5860 19180 5900
rect 19220 5860 23020 5900
rect 23060 5860 23069 5900
rect 26947 5860 26956 5900
rect 26996 5860 33100 5900
rect 33140 5860 33149 5900
rect 34915 5860 34924 5900
rect 34964 5860 39916 5900
rect 39956 5860 39965 5900
rect 46339 5860 46348 5900
rect 46388 5860 63052 5900
rect 63092 5860 63101 5900
rect 31843 5776 31852 5816
rect 31892 5776 36652 5816
rect 36692 5776 36701 5816
rect 67843 5776 67852 5816
rect 67892 5776 74380 5816
rect 74420 5776 74429 5816
rect 34243 5692 34252 5732
rect 34292 5692 40300 5732
rect 40340 5692 40349 5732
rect 61219 5692 61228 5732
rect 61268 5692 76876 5732
rect 76916 5692 77836 5732
rect 77876 5692 77885 5732
rect 1699 5608 1708 5648
rect 1748 5608 2540 5648
rect 30883 5608 30892 5648
rect 30932 5608 43660 5648
rect 43700 5608 43709 5648
rect 71971 5608 71980 5648
rect 72020 5608 84364 5648
rect 84404 5608 84413 5648
rect 90700 5608 97516 5648
rect 97556 5608 97565 5648
rect 2500 5564 2540 5608
rect 90700 5564 90740 5608
rect 2500 5524 32716 5564
rect 32756 5524 32765 5564
rect 56611 5524 56620 5564
rect 56660 5524 60460 5564
rect 60500 5524 60509 5564
rect 74467 5524 74476 5564
rect 74516 5524 90740 5564
rect 36547 5440 36556 5480
rect 36596 5440 41740 5480
rect 41780 5440 41789 5480
rect 55420 5440 64588 5480
rect 64628 5440 64637 5480
rect 72931 5440 72940 5480
rect 72980 5440 79756 5480
rect 79796 5440 79805 5480
rect 55420 5396 55460 5440
rect 52195 5356 52204 5396
rect 52244 5356 55460 5396
rect 3679 5335 4065 5354
rect 3679 5312 3745 5335
rect 3831 5312 3913 5335
rect 3999 5312 4065 5335
rect 3679 5272 3688 5312
rect 3728 5272 3745 5312
rect 3831 5272 3852 5312
rect 3892 5272 3913 5312
rect 3999 5272 4016 5312
rect 4056 5272 4065 5312
rect 3679 5249 3745 5272
rect 3831 5249 3913 5272
rect 3999 5249 4065 5272
rect 3679 5230 4065 5249
rect 18799 5335 19185 5354
rect 18799 5312 18865 5335
rect 18951 5312 19033 5335
rect 19119 5312 19185 5335
rect 18799 5272 18808 5312
rect 18848 5272 18865 5312
rect 18951 5272 18972 5312
rect 19012 5272 19033 5312
rect 19119 5272 19136 5312
rect 19176 5272 19185 5312
rect 18799 5249 18865 5272
rect 18951 5249 19033 5272
rect 19119 5249 19185 5272
rect 18799 5230 19185 5249
rect 33919 5335 34305 5354
rect 33919 5312 33985 5335
rect 34071 5312 34153 5335
rect 34239 5312 34305 5335
rect 33919 5272 33928 5312
rect 33968 5272 33985 5312
rect 34071 5272 34092 5312
rect 34132 5272 34153 5312
rect 34239 5272 34256 5312
rect 34296 5272 34305 5312
rect 33919 5249 33985 5272
rect 34071 5249 34153 5272
rect 34239 5249 34305 5272
rect 33919 5230 34305 5249
rect 49039 5335 49425 5354
rect 49039 5312 49105 5335
rect 49191 5312 49273 5335
rect 49359 5312 49425 5335
rect 49039 5272 49048 5312
rect 49088 5272 49105 5312
rect 49191 5272 49212 5312
rect 49252 5272 49273 5312
rect 49359 5272 49376 5312
rect 49416 5272 49425 5312
rect 49039 5249 49105 5272
rect 49191 5249 49273 5272
rect 49359 5249 49425 5272
rect 49039 5230 49425 5249
rect 64159 5335 64545 5354
rect 64159 5312 64225 5335
rect 64311 5312 64393 5335
rect 64479 5312 64545 5335
rect 64159 5272 64168 5312
rect 64208 5272 64225 5312
rect 64311 5272 64332 5312
rect 64372 5272 64393 5312
rect 64479 5272 64496 5312
rect 64536 5272 64545 5312
rect 64159 5249 64225 5272
rect 64311 5249 64393 5272
rect 64479 5249 64545 5272
rect 64159 5230 64545 5249
rect 79279 5335 79665 5354
rect 79279 5312 79345 5335
rect 79431 5312 79513 5335
rect 79599 5312 79665 5335
rect 79279 5272 79288 5312
rect 79328 5272 79345 5312
rect 79431 5272 79452 5312
rect 79492 5272 79513 5312
rect 79599 5272 79616 5312
rect 79656 5272 79665 5312
rect 79279 5249 79345 5272
rect 79431 5249 79513 5272
rect 79599 5249 79665 5272
rect 79279 5230 79665 5249
rect 94399 5335 94785 5354
rect 94399 5312 94465 5335
rect 94551 5312 94633 5335
rect 94719 5312 94785 5335
rect 94399 5272 94408 5312
rect 94448 5272 94465 5312
rect 94551 5272 94572 5312
rect 94612 5272 94633 5312
rect 94719 5272 94736 5312
rect 94776 5272 94785 5312
rect 94399 5249 94465 5272
rect 94551 5249 94633 5272
rect 94719 5249 94785 5272
rect 94399 5230 94785 5249
rect 21379 5020 21388 5060
rect 21428 5020 24652 5060
rect 24692 5020 24701 5060
rect 75139 5020 75148 5060
rect 75188 5020 76684 5060
rect 76724 5020 76733 5060
rect 82531 5020 82540 5060
rect 82580 5020 85612 5060
rect 85652 5020 85661 5060
rect 2083 4936 2092 4976
rect 2132 4936 34252 4976
rect 34292 4936 34301 4976
rect 76003 4936 76012 4976
rect 76052 4936 76780 4976
rect 76820 4936 76829 4976
rect 80611 4936 80620 4976
rect 80660 4936 97708 4976
rect 97748 4936 97757 4976
rect 97892 4936 98092 4976
rect 98132 4936 98141 4976
rect 97892 4892 97932 4936
rect 17539 4852 17548 4892
rect 17588 4852 24364 4892
rect 24404 4852 27628 4892
rect 27668 4852 27677 4892
rect 34819 4852 34828 4892
rect 34868 4852 39724 4892
rect 39764 4852 39773 4892
rect 44227 4852 44236 4892
rect 44276 4852 63244 4892
rect 63284 4852 63293 4892
rect 81859 4852 81868 4892
rect 81908 4852 97932 4892
rect 21283 4768 21292 4808
rect 21332 4768 25516 4808
rect 25556 4768 25565 4808
rect 72067 4768 72076 4808
rect 72116 4768 88492 4808
rect 88532 4768 88541 4808
rect 18499 4684 18508 4724
rect 18548 4684 25036 4724
rect 25076 4684 25085 4724
rect 32707 4684 32716 4724
rect 32756 4684 35788 4724
rect 35828 4684 35837 4724
rect 72835 4684 72844 4724
rect 72884 4684 88972 4724
rect 89012 4684 89021 4724
rect 67555 4600 67564 4640
rect 67604 4600 69964 4640
rect 70004 4600 71884 4640
rect 71924 4600 73516 4640
rect 73556 4600 73565 4640
rect 4919 4579 5305 4598
rect 4919 4556 4985 4579
rect 5071 4556 5153 4579
rect 5239 4556 5305 4579
rect 4919 4516 4928 4556
rect 4968 4516 4985 4556
rect 5071 4516 5092 4556
rect 5132 4516 5153 4556
rect 5239 4516 5256 4556
rect 5296 4516 5305 4556
rect 2090 4495 2214 4514
rect 2090 4409 2109 4495
rect 2195 4472 2214 4495
rect 4919 4493 4985 4516
rect 5071 4493 5153 4516
rect 5239 4493 5305 4516
rect 4919 4474 5305 4493
rect 20039 4579 20425 4598
rect 20039 4556 20105 4579
rect 20191 4556 20273 4579
rect 20359 4556 20425 4579
rect 20039 4516 20048 4556
rect 20088 4516 20105 4556
rect 20191 4516 20212 4556
rect 20252 4516 20273 4556
rect 20359 4516 20376 4556
rect 20416 4516 20425 4556
rect 20039 4493 20105 4516
rect 20191 4493 20273 4516
rect 20359 4493 20425 4516
rect 20039 4474 20425 4493
rect 35159 4579 35545 4598
rect 35159 4556 35225 4579
rect 35311 4556 35393 4579
rect 35479 4556 35545 4579
rect 35159 4516 35168 4556
rect 35208 4516 35225 4556
rect 35311 4516 35332 4556
rect 35372 4516 35393 4556
rect 35479 4516 35496 4556
rect 35536 4516 35545 4556
rect 35159 4493 35225 4516
rect 35311 4493 35393 4516
rect 35479 4493 35545 4516
rect 35159 4474 35545 4493
rect 50279 4579 50665 4598
rect 50279 4556 50345 4579
rect 50431 4556 50513 4579
rect 50599 4556 50665 4579
rect 50279 4516 50288 4556
rect 50328 4516 50345 4556
rect 50431 4516 50452 4556
rect 50492 4516 50513 4556
rect 50599 4516 50616 4556
rect 50656 4516 50665 4556
rect 50279 4493 50345 4516
rect 50431 4493 50513 4516
rect 50599 4493 50665 4516
rect 50279 4474 50665 4493
rect 65399 4579 65785 4598
rect 65399 4556 65465 4579
rect 65551 4556 65633 4579
rect 65719 4556 65785 4579
rect 65399 4516 65408 4556
rect 65448 4516 65465 4556
rect 65551 4516 65572 4556
rect 65612 4516 65633 4556
rect 65719 4516 65736 4556
rect 65776 4516 65785 4556
rect 65399 4493 65465 4516
rect 65551 4493 65633 4516
rect 65719 4493 65785 4516
rect 65399 4474 65785 4493
rect 80519 4579 80905 4598
rect 80519 4556 80585 4579
rect 80671 4556 80753 4579
rect 80839 4556 80905 4579
rect 80519 4516 80528 4556
rect 80568 4516 80585 4556
rect 80671 4516 80692 4556
rect 80732 4516 80753 4556
rect 80839 4516 80856 4556
rect 80896 4516 80905 4556
rect 80519 4493 80585 4516
rect 80671 4493 80753 4516
rect 80839 4493 80905 4516
rect 80519 4474 80905 4493
rect 95639 4579 96025 4598
rect 95639 4556 95705 4579
rect 95791 4556 95873 4579
rect 95959 4556 96025 4579
rect 95639 4516 95648 4556
rect 95688 4516 95705 4556
rect 95791 4516 95812 4556
rect 95852 4516 95873 4556
rect 95959 4516 95976 4556
rect 96016 4516 96025 4556
rect 95639 4493 95705 4516
rect 95791 4493 95873 4516
rect 95959 4493 96025 4516
rect 95639 4474 96025 4493
rect 2195 4432 2476 4472
rect 2516 4432 2525 4472
rect 2195 4409 2214 4432
rect 2090 4390 2214 4409
rect 33098 4411 33222 4430
rect 33098 4325 33117 4411
rect 33203 4388 33222 4411
rect 33203 4348 35020 4388
rect 35060 4348 35069 4388
rect 50371 4348 50380 4388
rect 50420 4348 61804 4388
rect 61844 4348 61853 4388
rect 33203 4325 33222 4348
rect 33098 4306 33222 4325
rect 17347 4264 17356 4304
rect 17396 4264 22732 4304
rect 22772 4264 22781 4304
rect 65443 4264 65452 4304
rect 65492 4264 67948 4304
rect 67988 4264 70540 4304
rect 70580 4264 70589 4304
rect 72547 4264 72556 4304
rect 72596 4264 87724 4304
rect 87764 4264 87773 4304
rect 19555 4180 19564 4220
rect 19604 4180 19948 4220
rect 19988 4180 20180 4220
rect 20227 4180 20236 4220
rect 20276 4180 21292 4220
rect 21332 4180 21341 4220
rect 27212 4180 28588 4220
rect 28628 4180 28637 4220
rect 49123 4180 49132 4220
rect 49172 4180 57964 4220
rect 58004 4180 58013 4220
rect 64771 4180 64780 4220
rect 64820 4180 67084 4220
rect 67124 4180 75148 4220
rect 75188 4180 75197 4220
rect 20140 4136 20180 4180
rect 27212 4136 27252 4180
rect 20140 4096 23788 4136
rect 23828 4096 27252 4136
rect 27619 4096 27628 4136
rect 27668 4096 29932 4136
rect 29972 4096 34060 4136
rect 34100 4096 34540 4136
rect 34580 4096 34924 4136
rect 34964 4096 34973 4136
rect 36643 4096 36652 4136
rect 36692 4096 42988 4136
rect 43028 4096 43037 4136
rect 73699 4096 73708 4136
rect 73748 4096 86284 4136
rect 86324 4096 86333 4136
rect 28994 3991 29118 4010
rect 28994 3905 29013 3991
rect 29099 3968 29118 3991
rect 29108 3928 29118 3968
rect 49699 3928 49708 3968
rect 49748 3928 58252 3968
rect 58292 3928 58301 3968
rect 29099 3905 29118 3928
rect 28994 3886 29118 3905
rect 3679 3823 4065 3842
rect 3679 3800 3745 3823
rect 3831 3800 3913 3823
rect 3999 3800 4065 3823
rect 3679 3760 3688 3800
rect 3728 3760 3745 3800
rect 3831 3760 3852 3800
rect 3892 3760 3913 3800
rect 3999 3760 4016 3800
rect 4056 3760 4065 3800
rect 3679 3737 3745 3760
rect 3831 3737 3913 3760
rect 3999 3737 4065 3760
rect 3679 3718 4065 3737
rect 18799 3823 19185 3842
rect 18799 3800 18865 3823
rect 18951 3800 19033 3823
rect 19119 3800 19185 3823
rect 18799 3760 18808 3800
rect 18848 3760 18865 3800
rect 18951 3760 18972 3800
rect 19012 3760 19033 3800
rect 19119 3760 19136 3800
rect 19176 3760 19185 3800
rect 18799 3737 18865 3760
rect 18951 3737 19033 3760
rect 19119 3737 19185 3760
rect 18799 3718 19185 3737
rect 33919 3823 34305 3842
rect 33919 3800 33985 3823
rect 34071 3800 34153 3823
rect 34239 3800 34305 3823
rect 49039 3823 49425 3842
rect 49039 3800 49105 3823
rect 49191 3800 49273 3823
rect 49359 3800 49425 3823
rect 33919 3760 33928 3800
rect 33968 3760 33985 3800
rect 34071 3760 34092 3800
rect 34132 3760 34153 3800
rect 34239 3760 34256 3800
rect 34296 3760 34305 3800
rect 38659 3760 38668 3800
rect 38708 3760 40300 3800
rect 40340 3760 40349 3800
rect 49039 3760 49048 3800
rect 49088 3760 49105 3800
rect 49191 3760 49212 3800
rect 49252 3760 49273 3800
rect 49359 3760 49376 3800
rect 49416 3760 49425 3800
rect 33919 3737 33985 3760
rect 34071 3737 34153 3760
rect 34239 3737 34305 3760
rect 33919 3718 34305 3737
rect 49039 3737 49105 3760
rect 49191 3737 49273 3760
rect 49359 3737 49425 3760
rect 49039 3718 49425 3737
rect 64159 3823 64545 3842
rect 64159 3800 64225 3823
rect 64311 3800 64393 3823
rect 64479 3800 64545 3823
rect 64159 3760 64168 3800
rect 64208 3760 64225 3800
rect 64311 3760 64332 3800
rect 64372 3760 64393 3800
rect 64479 3760 64496 3800
rect 64536 3760 64545 3800
rect 64159 3737 64225 3760
rect 64311 3737 64393 3760
rect 64479 3737 64545 3760
rect 64159 3718 64545 3737
rect 79279 3823 79665 3842
rect 79279 3800 79345 3823
rect 79431 3800 79513 3823
rect 79599 3800 79665 3823
rect 79279 3760 79288 3800
rect 79328 3760 79345 3800
rect 79431 3760 79452 3800
rect 79492 3760 79513 3800
rect 79599 3760 79616 3800
rect 79656 3760 79665 3800
rect 79279 3737 79345 3760
rect 79431 3737 79513 3760
rect 79599 3737 79665 3760
rect 79279 3718 79665 3737
rect 94399 3823 94785 3842
rect 94399 3800 94465 3823
rect 94551 3800 94633 3823
rect 94719 3800 94785 3823
rect 94399 3760 94408 3800
rect 94448 3760 94465 3800
rect 94551 3760 94572 3800
rect 94612 3760 94633 3800
rect 94719 3760 94736 3800
rect 94776 3760 94785 3800
rect 94399 3737 94465 3760
rect 94551 3737 94633 3760
rect 94719 3737 94785 3760
rect 94399 3718 94785 3737
rect 20131 3676 20140 3716
rect 20180 3676 33484 3716
rect 33524 3676 33533 3716
rect 6979 3592 6988 3632
rect 7028 3592 22348 3632
rect 22388 3592 22397 3632
rect 67075 3592 67084 3632
rect 67124 3592 95884 3632
rect 95924 3592 95933 3632
rect 2132 3508 19756 3548
rect 19796 3508 19805 3548
rect 32995 3508 33004 3548
rect 33044 3508 42300 3548
rect 49507 3508 49516 3548
rect 49556 3508 55460 3548
rect 60451 3508 60460 3548
rect 60500 3508 64280 3548
rect 64771 3508 64780 3548
rect 64820 3508 92916 3548
rect 1634 3487 1758 3506
rect 1634 3464 1653 3487
rect 1603 3424 1612 3464
rect 1652 3424 1653 3464
rect 1634 3401 1653 3424
rect 1739 3401 1758 3487
rect 2132 3464 2172 3508
rect 42260 3464 42300 3508
rect 55420 3464 55460 3508
rect 64240 3464 64280 3508
rect 92876 3464 92916 3508
rect 1987 3424 1996 3464
rect 2036 3424 2172 3464
rect 2371 3424 2380 3464
rect 2420 3424 2540 3464
rect 18499 3424 18508 3464
rect 18548 3424 25420 3464
rect 25460 3424 25469 3464
rect 37699 3424 37708 3464
rect 37748 3424 41600 3464
rect 42260 3424 43372 3464
rect 43412 3424 43421 3464
rect 43628 3424 47980 3464
rect 48020 3424 48029 3464
rect 55420 3424 60748 3464
rect 60788 3424 60797 3464
rect 64240 3424 92460 3464
rect 92876 3424 95500 3464
rect 95540 3424 95549 3464
rect 95612 3424 96652 3464
rect 96692 3424 96701 3464
rect 1634 3382 1758 3401
rect 2500 3380 2540 3424
rect 41560 3380 41600 3424
rect 43628 3380 43668 3424
rect 92420 3380 92460 3424
rect 95612 3380 95652 3424
rect 2500 3340 16396 3380
rect 16436 3340 16445 3380
rect 41560 3340 43668 3380
rect 80611 3340 80620 3380
rect 80660 3340 91948 3380
rect 91988 3340 91997 3380
rect 92420 3340 95652 3380
rect 1219 3256 1228 3296
rect 1268 3256 19948 3296
rect 19988 3256 19997 3296
rect 49219 3256 49228 3296
rect 49268 3256 58060 3296
rect 58100 3256 58109 3296
rect 60259 3256 60268 3296
rect 60308 3256 94732 3296
rect 94772 3256 94781 3296
rect 59491 3172 59500 3212
rect 59540 3172 90740 3212
rect 92035 3172 92044 3212
rect 92084 3172 97420 3212
rect 97460 3172 97469 3212
rect 90700 3128 90740 3172
rect 90700 3088 95116 3128
rect 95156 3088 95165 3128
rect 4919 3067 5305 3086
rect 4919 3044 4985 3067
rect 5071 3044 5153 3067
rect 5239 3044 5305 3067
rect 4919 3004 4928 3044
rect 4968 3004 4985 3044
rect 5071 3004 5092 3044
rect 5132 3004 5153 3044
rect 5239 3004 5256 3044
rect 5296 3004 5305 3044
rect 4919 2981 4985 3004
rect 5071 2981 5153 3004
rect 5239 2981 5305 3004
rect 4919 2962 5305 2981
rect 20039 3067 20425 3086
rect 20039 3044 20105 3067
rect 20191 3044 20273 3067
rect 20359 3044 20425 3067
rect 20039 3004 20048 3044
rect 20088 3004 20105 3044
rect 20191 3004 20212 3044
rect 20252 3004 20273 3044
rect 20359 3004 20376 3044
rect 20416 3004 20425 3044
rect 20039 2981 20105 3004
rect 20191 2981 20273 3004
rect 20359 2981 20425 3004
rect 20039 2962 20425 2981
rect 35159 3067 35545 3086
rect 35159 3044 35225 3067
rect 35311 3044 35393 3067
rect 35479 3044 35545 3067
rect 35159 3004 35168 3044
rect 35208 3004 35225 3044
rect 35311 3004 35332 3044
rect 35372 3004 35393 3044
rect 35479 3004 35496 3044
rect 35536 3004 35545 3044
rect 35159 2981 35225 3004
rect 35311 2981 35393 3004
rect 35479 2981 35545 3004
rect 35159 2962 35545 2981
rect 50279 3067 50665 3086
rect 50279 3044 50345 3067
rect 50431 3044 50513 3067
rect 50599 3044 50665 3067
rect 50279 3004 50288 3044
rect 50328 3004 50345 3044
rect 50431 3004 50452 3044
rect 50492 3004 50513 3044
rect 50599 3004 50616 3044
rect 50656 3004 50665 3044
rect 50279 2981 50345 3004
rect 50431 2981 50513 3004
rect 50599 2981 50665 3004
rect 50279 2962 50665 2981
rect 65399 3067 65785 3086
rect 65399 3044 65465 3067
rect 65551 3044 65633 3067
rect 65719 3044 65785 3067
rect 65399 3004 65408 3044
rect 65448 3004 65465 3044
rect 65551 3004 65572 3044
rect 65612 3004 65633 3044
rect 65719 3004 65736 3044
rect 65776 3004 65785 3044
rect 65399 2981 65465 3004
rect 65551 2981 65633 3004
rect 65719 2981 65785 3004
rect 65399 2962 65785 2981
rect 80519 3067 80905 3086
rect 80519 3044 80585 3067
rect 80671 3044 80753 3067
rect 80839 3044 80905 3067
rect 80519 3004 80528 3044
rect 80568 3004 80585 3044
rect 80671 3004 80692 3044
rect 80732 3004 80753 3044
rect 80839 3004 80856 3044
rect 80896 3004 80905 3044
rect 80519 2981 80585 3004
rect 80671 2981 80753 3004
rect 80839 2981 80905 3004
rect 80519 2962 80905 2981
rect 95639 3067 96025 3086
rect 95639 3044 95705 3067
rect 95791 3044 95873 3067
rect 95959 3044 96025 3067
rect 95639 3004 95648 3044
rect 95688 3004 95705 3044
rect 95791 3004 95812 3044
rect 95852 3004 95873 3044
rect 95959 3004 95976 3044
rect 96016 3004 96025 3044
rect 95639 2981 95705 3004
rect 95791 2981 95873 3004
rect 95959 2981 96025 3004
rect 95639 2962 96025 2981
<< via5 >>
rect 3745 11360 3831 11383
rect 3913 11360 3999 11383
rect 3745 11320 3770 11360
rect 3770 11320 3810 11360
rect 3810 11320 3831 11360
rect 3913 11320 3934 11360
rect 3934 11320 3974 11360
rect 3974 11320 3999 11360
rect 3745 11297 3831 11320
rect 3913 11297 3999 11320
rect 18865 11360 18951 11383
rect 19033 11360 19119 11383
rect 18865 11320 18890 11360
rect 18890 11320 18930 11360
rect 18930 11320 18951 11360
rect 19033 11320 19054 11360
rect 19054 11320 19094 11360
rect 19094 11320 19119 11360
rect 18865 11297 18951 11320
rect 19033 11297 19119 11320
rect 33985 11360 34071 11383
rect 34153 11360 34239 11383
rect 33985 11320 34010 11360
rect 34010 11320 34050 11360
rect 34050 11320 34071 11360
rect 34153 11320 34174 11360
rect 34174 11320 34214 11360
rect 34214 11320 34239 11360
rect 33985 11297 34071 11320
rect 34153 11297 34239 11320
rect 49105 11360 49191 11383
rect 49273 11360 49359 11383
rect 49105 11320 49130 11360
rect 49130 11320 49170 11360
rect 49170 11320 49191 11360
rect 49273 11320 49294 11360
rect 49294 11320 49334 11360
rect 49334 11320 49359 11360
rect 49105 11297 49191 11320
rect 49273 11297 49359 11320
rect 64225 11360 64311 11383
rect 64393 11360 64479 11383
rect 64225 11320 64250 11360
rect 64250 11320 64290 11360
rect 64290 11320 64311 11360
rect 64393 11320 64414 11360
rect 64414 11320 64454 11360
rect 64454 11320 64479 11360
rect 64225 11297 64311 11320
rect 64393 11297 64479 11320
rect 79345 11360 79431 11383
rect 79513 11360 79599 11383
rect 79345 11320 79370 11360
rect 79370 11320 79410 11360
rect 79410 11320 79431 11360
rect 79513 11320 79534 11360
rect 79534 11320 79574 11360
rect 79574 11320 79599 11360
rect 79345 11297 79431 11320
rect 79513 11297 79599 11320
rect 94465 11360 94551 11383
rect 94633 11360 94719 11383
rect 94465 11320 94490 11360
rect 94490 11320 94530 11360
rect 94530 11320 94551 11360
rect 94633 11320 94654 11360
rect 94654 11320 94694 11360
rect 94694 11320 94719 11360
rect 94465 11297 94551 11320
rect 94633 11297 94719 11320
rect 4985 10604 5071 10627
rect 5153 10604 5239 10627
rect 4985 10564 5010 10604
rect 5010 10564 5050 10604
rect 5050 10564 5071 10604
rect 5153 10564 5174 10604
rect 5174 10564 5214 10604
rect 5214 10564 5239 10604
rect 4985 10541 5071 10564
rect 5153 10541 5239 10564
rect 20105 10604 20191 10627
rect 20273 10604 20359 10627
rect 20105 10564 20130 10604
rect 20130 10564 20170 10604
rect 20170 10564 20191 10604
rect 20273 10564 20294 10604
rect 20294 10564 20334 10604
rect 20334 10564 20359 10604
rect 20105 10541 20191 10564
rect 20273 10541 20359 10564
rect 35225 10604 35311 10627
rect 35393 10604 35479 10627
rect 35225 10564 35250 10604
rect 35250 10564 35290 10604
rect 35290 10564 35311 10604
rect 35393 10564 35414 10604
rect 35414 10564 35454 10604
rect 35454 10564 35479 10604
rect 35225 10541 35311 10564
rect 35393 10541 35479 10564
rect 50345 10604 50431 10627
rect 50513 10604 50599 10627
rect 50345 10564 50370 10604
rect 50370 10564 50410 10604
rect 50410 10564 50431 10604
rect 50513 10564 50534 10604
rect 50534 10564 50574 10604
rect 50574 10564 50599 10604
rect 50345 10541 50431 10564
rect 50513 10541 50599 10564
rect 65465 10604 65551 10627
rect 65633 10604 65719 10627
rect 65465 10564 65490 10604
rect 65490 10564 65530 10604
rect 65530 10564 65551 10604
rect 65633 10564 65654 10604
rect 65654 10564 65694 10604
rect 65694 10564 65719 10604
rect 65465 10541 65551 10564
rect 65633 10541 65719 10564
rect 80585 10604 80671 10627
rect 80753 10604 80839 10627
rect 80585 10564 80610 10604
rect 80610 10564 80650 10604
rect 80650 10564 80671 10604
rect 80753 10564 80774 10604
rect 80774 10564 80814 10604
rect 80814 10564 80839 10604
rect 80585 10541 80671 10564
rect 80753 10541 80839 10564
rect 95705 10604 95791 10627
rect 95873 10604 95959 10627
rect 95705 10564 95730 10604
rect 95730 10564 95770 10604
rect 95770 10564 95791 10604
rect 95873 10564 95894 10604
rect 95894 10564 95934 10604
rect 95934 10564 95959 10604
rect 95705 10541 95791 10564
rect 95873 10541 95959 10564
rect 3745 9848 3831 9871
rect 3913 9848 3999 9871
rect 3745 9808 3770 9848
rect 3770 9808 3810 9848
rect 3810 9808 3831 9848
rect 3913 9808 3934 9848
rect 3934 9808 3974 9848
rect 3974 9808 3999 9848
rect 3745 9785 3831 9808
rect 3913 9785 3999 9808
rect 18865 9848 18951 9871
rect 19033 9848 19119 9871
rect 18865 9808 18890 9848
rect 18890 9808 18930 9848
rect 18930 9808 18951 9848
rect 19033 9808 19054 9848
rect 19054 9808 19094 9848
rect 19094 9808 19119 9848
rect 18865 9785 18951 9808
rect 19033 9785 19119 9808
rect 33985 9848 34071 9871
rect 34153 9848 34239 9871
rect 33985 9808 34010 9848
rect 34010 9808 34050 9848
rect 34050 9808 34071 9848
rect 34153 9808 34174 9848
rect 34174 9808 34214 9848
rect 34214 9808 34239 9848
rect 33985 9785 34071 9808
rect 34153 9785 34239 9808
rect 49105 9848 49191 9871
rect 49273 9848 49359 9871
rect 49105 9808 49130 9848
rect 49130 9808 49170 9848
rect 49170 9808 49191 9848
rect 49273 9808 49294 9848
rect 49294 9808 49334 9848
rect 49334 9808 49359 9848
rect 49105 9785 49191 9808
rect 49273 9785 49359 9808
rect 64225 9848 64311 9871
rect 64393 9848 64479 9871
rect 64225 9808 64250 9848
rect 64250 9808 64290 9848
rect 64290 9808 64311 9848
rect 64393 9808 64414 9848
rect 64414 9808 64454 9848
rect 64454 9808 64479 9848
rect 64225 9785 64311 9808
rect 64393 9785 64479 9808
rect 79345 9848 79431 9871
rect 79513 9848 79599 9871
rect 79345 9808 79370 9848
rect 79370 9808 79410 9848
rect 79410 9808 79431 9848
rect 79513 9808 79534 9848
rect 79534 9808 79574 9848
rect 79574 9808 79599 9848
rect 79345 9785 79431 9808
rect 79513 9785 79599 9808
rect 94465 9848 94551 9871
rect 94633 9848 94719 9871
rect 94465 9808 94490 9848
rect 94490 9808 94530 9848
rect 94530 9808 94551 9848
rect 94633 9808 94654 9848
rect 94654 9808 94694 9848
rect 94694 9808 94719 9848
rect 94465 9785 94551 9808
rect 94633 9785 94719 9808
rect 4985 9092 5071 9115
rect 5153 9092 5239 9115
rect 4985 9052 5010 9092
rect 5010 9052 5050 9092
rect 5050 9052 5071 9092
rect 5153 9052 5174 9092
rect 5174 9052 5214 9092
rect 5214 9052 5239 9092
rect 4985 9029 5071 9052
rect 5153 9029 5239 9052
rect 20105 9092 20191 9115
rect 20273 9092 20359 9115
rect 20105 9052 20130 9092
rect 20130 9052 20170 9092
rect 20170 9052 20191 9092
rect 20273 9052 20294 9092
rect 20294 9052 20334 9092
rect 20334 9052 20359 9092
rect 20105 9029 20191 9052
rect 20273 9029 20359 9052
rect 35225 9092 35311 9115
rect 35393 9092 35479 9115
rect 35225 9052 35250 9092
rect 35250 9052 35290 9092
rect 35290 9052 35311 9092
rect 35393 9052 35414 9092
rect 35414 9052 35454 9092
rect 35454 9052 35479 9092
rect 35225 9029 35311 9052
rect 35393 9029 35479 9052
rect 50345 9092 50431 9115
rect 50513 9092 50599 9115
rect 50345 9052 50370 9092
rect 50370 9052 50410 9092
rect 50410 9052 50431 9092
rect 50513 9052 50534 9092
rect 50534 9052 50574 9092
rect 50574 9052 50599 9092
rect 50345 9029 50431 9052
rect 50513 9029 50599 9052
rect 65465 9092 65551 9115
rect 65633 9092 65719 9115
rect 65465 9052 65490 9092
rect 65490 9052 65530 9092
rect 65530 9052 65551 9092
rect 65633 9052 65654 9092
rect 65654 9052 65694 9092
rect 65694 9052 65719 9092
rect 65465 9029 65551 9052
rect 65633 9029 65719 9052
rect 80585 9092 80671 9115
rect 80753 9092 80839 9115
rect 80585 9052 80610 9092
rect 80610 9052 80650 9092
rect 80650 9052 80671 9092
rect 80753 9052 80774 9092
rect 80774 9052 80814 9092
rect 80814 9052 80839 9092
rect 80585 9029 80671 9052
rect 80753 9029 80839 9052
rect 95705 9092 95791 9115
rect 95873 9092 95959 9115
rect 95705 9052 95730 9092
rect 95730 9052 95770 9092
rect 95770 9052 95791 9092
rect 95873 9052 95894 9092
rect 95894 9052 95934 9092
rect 95934 9052 95959 9092
rect 95705 9029 95791 9052
rect 95873 9029 95959 9052
rect 3745 8336 3831 8359
rect 3913 8336 3999 8359
rect 3745 8296 3770 8336
rect 3770 8296 3810 8336
rect 3810 8296 3831 8336
rect 3913 8296 3934 8336
rect 3934 8296 3974 8336
rect 3974 8296 3999 8336
rect 3745 8273 3831 8296
rect 3913 8273 3999 8296
rect 18865 8336 18951 8359
rect 19033 8336 19119 8359
rect 18865 8296 18890 8336
rect 18890 8296 18930 8336
rect 18930 8296 18951 8336
rect 19033 8296 19054 8336
rect 19054 8296 19094 8336
rect 19094 8296 19119 8336
rect 18865 8273 18951 8296
rect 19033 8273 19119 8296
rect 33985 8336 34071 8359
rect 34153 8336 34239 8359
rect 33985 8296 34010 8336
rect 34010 8296 34050 8336
rect 34050 8296 34071 8336
rect 34153 8296 34174 8336
rect 34174 8296 34214 8336
rect 34214 8296 34239 8336
rect 33985 8273 34071 8296
rect 34153 8273 34239 8296
rect 49105 8336 49191 8359
rect 49273 8336 49359 8359
rect 49105 8296 49130 8336
rect 49130 8296 49170 8336
rect 49170 8296 49191 8336
rect 49273 8296 49294 8336
rect 49294 8296 49334 8336
rect 49334 8296 49359 8336
rect 49105 8273 49191 8296
rect 49273 8273 49359 8296
rect 64225 8336 64311 8359
rect 64393 8336 64479 8359
rect 64225 8296 64250 8336
rect 64250 8296 64290 8336
rect 64290 8296 64311 8336
rect 64393 8296 64414 8336
rect 64414 8296 64454 8336
rect 64454 8296 64479 8336
rect 64225 8273 64311 8296
rect 64393 8273 64479 8296
rect 79345 8336 79431 8359
rect 79513 8336 79599 8359
rect 79345 8296 79370 8336
rect 79370 8296 79410 8336
rect 79410 8296 79431 8336
rect 79513 8296 79534 8336
rect 79534 8296 79574 8336
rect 79574 8296 79599 8336
rect 79345 8273 79431 8296
rect 79513 8273 79599 8296
rect 94465 8336 94551 8359
rect 94633 8336 94719 8359
rect 94465 8296 94490 8336
rect 94490 8296 94530 8336
rect 94530 8296 94551 8336
rect 94633 8296 94654 8336
rect 94654 8296 94694 8336
rect 94694 8296 94719 8336
rect 94465 8273 94551 8296
rect 94633 8273 94719 8296
rect 4985 7580 5071 7603
rect 5153 7580 5239 7603
rect 4985 7540 5010 7580
rect 5010 7540 5050 7580
rect 5050 7540 5071 7580
rect 5153 7540 5174 7580
rect 5174 7540 5214 7580
rect 5214 7540 5239 7580
rect 4985 7517 5071 7540
rect 5153 7517 5239 7540
rect 20105 7580 20191 7603
rect 20273 7580 20359 7603
rect 20105 7540 20130 7580
rect 20130 7540 20170 7580
rect 20170 7540 20191 7580
rect 20273 7540 20294 7580
rect 20294 7540 20334 7580
rect 20334 7540 20359 7580
rect 20105 7517 20191 7540
rect 20273 7517 20359 7540
rect 35225 7580 35311 7603
rect 35393 7580 35479 7603
rect 35225 7540 35250 7580
rect 35250 7540 35290 7580
rect 35290 7540 35311 7580
rect 35393 7540 35414 7580
rect 35414 7540 35454 7580
rect 35454 7540 35479 7580
rect 35225 7517 35311 7540
rect 35393 7517 35479 7540
rect 50345 7580 50431 7603
rect 50513 7580 50599 7603
rect 50345 7540 50370 7580
rect 50370 7540 50410 7580
rect 50410 7540 50431 7580
rect 50513 7540 50534 7580
rect 50534 7540 50574 7580
rect 50574 7540 50599 7580
rect 50345 7517 50431 7540
rect 50513 7517 50599 7540
rect 65465 7580 65551 7603
rect 65633 7580 65719 7603
rect 80585 7580 80671 7603
rect 80753 7580 80839 7603
rect 95705 7580 95791 7603
rect 95873 7580 95959 7603
rect 65465 7540 65490 7580
rect 65490 7540 65530 7580
rect 65530 7540 65551 7580
rect 65633 7540 65654 7580
rect 65654 7540 65694 7580
rect 65694 7540 65719 7580
rect 80585 7540 80610 7580
rect 80610 7540 80650 7580
rect 80650 7540 80671 7580
rect 80753 7540 80774 7580
rect 80774 7540 80814 7580
rect 80814 7540 80839 7580
rect 95705 7540 95730 7580
rect 95730 7540 95770 7580
rect 95770 7540 95791 7580
rect 95873 7540 95894 7580
rect 95894 7540 95934 7580
rect 95934 7540 95959 7580
rect 65465 7517 65551 7540
rect 65633 7517 65719 7540
rect 80585 7517 80671 7540
rect 80753 7517 80839 7540
rect 95705 7517 95791 7540
rect 95873 7517 95959 7540
rect 3745 6824 3831 6847
rect 3913 6824 3999 6847
rect 3745 6784 3770 6824
rect 3770 6784 3810 6824
rect 3810 6784 3831 6824
rect 3913 6784 3934 6824
rect 3934 6784 3974 6824
rect 3974 6784 3999 6824
rect 3745 6761 3831 6784
rect 3913 6761 3999 6784
rect 18865 6824 18951 6847
rect 19033 6824 19119 6847
rect 18865 6784 18890 6824
rect 18890 6784 18930 6824
rect 18930 6784 18951 6824
rect 19033 6784 19054 6824
rect 19054 6784 19094 6824
rect 19094 6784 19119 6824
rect 18865 6761 18951 6784
rect 19033 6761 19119 6784
rect 33985 6824 34071 6847
rect 34153 6824 34239 6847
rect 33985 6784 34010 6824
rect 34010 6784 34050 6824
rect 34050 6784 34071 6824
rect 34153 6784 34174 6824
rect 34174 6784 34214 6824
rect 34214 6784 34239 6824
rect 33985 6761 34071 6784
rect 34153 6761 34239 6784
rect 49105 6824 49191 6847
rect 49273 6824 49359 6847
rect 49105 6784 49130 6824
rect 49130 6784 49170 6824
rect 49170 6784 49191 6824
rect 49273 6784 49294 6824
rect 49294 6784 49334 6824
rect 49334 6784 49359 6824
rect 49105 6761 49191 6784
rect 49273 6761 49359 6784
rect 64225 6824 64311 6847
rect 64393 6824 64479 6847
rect 64225 6784 64250 6824
rect 64250 6784 64290 6824
rect 64290 6784 64311 6824
rect 64393 6784 64414 6824
rect 64414 6784 64454 6824
rect 64454 6784 64479 6824
rect 64225 6761 64311 6784
rect 64393 6761 64479 6784
rect 79345 6824 79431 6847
rect 79513 6824 79599 6847
rect 79345 6784 79370 6824
rect 79370 6784 79410 6824
rect 79410 6784 79431 6824
rect 79513 6784 79534 6824
rect 79534 6784 79574 6824
rect 79574 6784 79599 6824
rect 79345 6761 79431 6784
rect 79513 6761 79599 6784
rect 94465 6824 94551 6847
rect 94633 6824 94719 6847
rect 94465 6784 94490 6824
rect 94490 6784 94530 6824
rect 94530 6784 94551 6824
rect 94633 6784 94654 6824
rect 94654 6784 94694 6824
rect 94694 6784 94719 6824
rect 94465 6761 94551 6784
rect 94633 6761 94719 6784
rect 4985 6068 5071 6091
rect 5153 6068 5239 6091
rect 4985 6028 5010 6068
rect 5010 6028 5050 6068
rect 5050 6028 5071 6068
rect 5153 6028 5174 6068
rect 5174 6028 5214 6068
rect 5214 6028 5239 6068
rect 4985 6005 5071 6028
rect 5153 6005 5239 6028
rect 20105 6068 20191 6091
rect 20273 6068 20359 6091
rect 20105 6028 20130 6068
rect 20130 6028 20170 6068
rect 20170 6028 20191 6068
rect 20273 6028 20294 6068
rect 20294 6028 20334 6068
rect 20334 6028 20359 6068
rect 20105 6005 20191 6028
rect 20273 6005 20359 6028
rect 35225 6068 35311 6091
rect 35393 6068 35479 6091
rect 35225 6028 35250 6068
rect 35250 6028 35290 6068
rect 35290 6028 35311 6068
rect 35393 6028 35414 6068
rect 35414 6028 35454 6068
rect 35454 6028 35479 6068
rect 35225 6005 35311 6028
rect 35393 6005 35479 6028
rect 50345 6068 50431 6091
rect 50513 6068 50599 6091
rect 50345 6028 50370 6068
rect 50370 6028 50410 6068
rect 50410 6028 50431 6068
rect 50513 6028 50534 6068
rect 50534 6028 50574 6068
rect 50574 6028 50599 6068
rect 50345 6005 50431 6028
rect 50513 6005 50599 6028
rect 65465 6068 65551 6091
rect 65633 6068 65719 6091
rect 65465 6028 65490 6068
rect 65490 6028 65530 6068
rect 65530 6028 65551 6068
rect 65633 6028 65654 6068
rect 65654 6028 65694 6068
rect 65694 6028 65719 6068
rect 65465 6005 65551 6028
rect 65633 6005 65719 6028
rect 80585 6068 80671 6091
rect 80753 6068 80839 6091
rect 80585 6028 80610 6068
rect 80610 6028 80650 6068
rect 80650 6028 80671 6068
rect 80753 6028 80774 6068
rect 80774 6028 80814 6068
rect 80814 6028 80839 6068
rect 80585 6005 80671 6028
rect 80753 6005 80839 6028
rect 95705 6068 95791 6091
rect 95873 6068 95959 6091
rect 95705 6028 95730 6068
rect 95730 6028 95770 6068
rect 95770 6028 95791 6068
rect 95873 6028 95894 6068
rect 95894 6028 95934 6068
rect 95934 6028 95959 6068
rect 95705 6005 95791 6028
rect 95873 6005 95959 6028
rect 3745 5312 3831 5335
rect 3913 5312 3999 5335
rect 3745 5272 3770 5312
rect 3770 5272 3810 5312
rect 3810 5272 3831 5312
rect 3913 5272 3934 5312
rect 3934 5272 3974 5312
rect 3974 5272 3999 5312
rect 3745 5249 3831 5272
rect 3913 5249 3999 5272
rect 18865 5312 18951 5335
rect 19033 5312 19119 5335
rect 18865 5272 18890 5312
rect 18890 5272 18930 5312
rect 18930 5272 18951 5312
rect 19033 5272 19054 5312
rect 19054 5272 19094 5312
rect 19094 5272 19119 5312
rect 18865 5249 18951 5272
rect 19033 5249 19119 5272
rect 33985 5312 34071 5335
rect 34153 5312 34239 5335
rect 33985 5272 34010 5312
rect 34010 5272 34050 5312
rect 34050 5272 34071 5312
rect 34153 5272 34174 5312
rect 34174 5272 34214 5312
rect 34214 5272 34239 5312
rect 33985 5249 34071 5272
rect 34153 5249 34239 5272
rect 49105 5312 49191 5335
rect 49273 5312 49359 5335
rect 49105 5272 49130 5312
rect 49130 5272 49170 5312
rect 49170 5272 49191 5312
rect 49273 5272 49294 5312
rect 49294 5272 49334 5312
rect 49334 5272 49359 5312
rect 49105 5249 49191 5272
rect 49273 5249 49359 5272
rect 64225 5312 64311 5335
rect 64393 5312 64479 5335
rect 64225 5272 64250 5312
rect 64250 5272 64290 5312
rect 64290 5272 64311 5312
rect 64393 5272 64414 5312
rect 64414 5272 64454 5312
rect 64454 5272 64479 5312
rect 64225 5249 64311 5272
rect 64393 5249 64479 5272
rect 79345 5312 79431 5335
rect 79513 5312 79599 5335
rect 79345 5272 79370 5312
rect 79370 5272 79410 5312
rect 79410 5272 79431 5312
rect 79513 5272 79534 5312
rect 79534 5272 79574 5312
rect 79574 5272 79599 5312
rect 79345 5249 79431 5272
rect 79513 5249 79599 5272
rect 94465 5312 94551 5335
rect 94633 5312 94719 5335
rect 94465 5272 94490 5312
rect 94490 5272 94530 5312
rect 94530 5272 94551 5312
rect 94633 5272 94654 5312
rect 94654 5272 94694 5312
rect 94694 5272 94719 5312
rect 94465 5249 94551 5272
rect 94633 5249 94719 5272
rect 4985 4556 5071 4579
rect 5153 4556 5239 4579
rect 4985 4516 5010 4556
rect 5010 4516 5050 4556
rect 5050 4516 5071 4556
rect 5153 4516 5174 4556
rect 5174 4516 5214 4556
rect 5214 4516 5239 4556
rect 2109 4409 2195 4495
rect 4985 4493 5071 4516
rect 5153 4493 5239 4516
rect 20105 4556 20191 4579
rect 20273 4556 20359 4579
rect 20105 4516 20130 4556
rect 20130 4516 20170 4556
rect 20170 4516 20191 4556
rect 20273 4516 20294 4556
rect 20294 4516 20334 4556
rect 20334 4516 20359 4556
rect 20105 4493 20191 4516
rect 20273 4493 20359 4516
rect 35225 4556 35311 4579
rect 35393 4556 35479 4579
rect 35225 4516 35250 4556
rect 35250 4516 35290 4556
rect 35290 4516 35311 4556
rect 35393 4516 35414 4556
rect 35414 4516 35454 4556
rect 35454 4516 35479 4556
rect 35225 4493 35311 4516
rect 35393 4493 35479 4516
rect 50345 4556 50431 4579
rect 50513 4556 50599 4579
rect 50345 4516 50370 4556
rect 50370 4516 50410 4556
rect 50410 4516 50431 4556
rect 50513 4516 50534 4556
rect 50534 4516 50574 4556
rect 50574 4516 50599 4556
rect 50345 4493 50431 4516
rect 50513 4493 50599 4516
rect 65465 4556 65551 4579
rect 65633 4556 65719 4579
rect 65465 4516 65490 4556
rect 65490 4516 65530 4556
rect 65530 4516 65551 4556
rect 65633 4516 65654 4556
rect 65654 4516 65694 4556
rect 65694 4516 65719 4556
rect 65465 4493 65551 4516
rect 65633 4493 65719 4516
rect 80585 4556 80671 4579
rect 80753 4556 80839 4579
rect 80585 4516 80610 4556
rect 80610 4516 80650 4556
rect 80650 4516 80671 4556
rect 80753 4516 80774 4556
rect 80774 4516 80814 4556
rect 80814 4516 80839 4556
rect 80585 4493 80671 4516
rect 80753 4493 80839 4516
rect 95705 4556 95791 4579
rect 95873 4556 95959 4579
rect 95705 4516 95730 4556
rect 95730 4516 95770 4556
rect 95770 4516 95791 4556
rect 95873 4516 95894 4556
rect 95894 4516 95934 4556
rect 95934 4516 95959 4556
rect 95705 4493 95791 4516
rect 95873 4493 95959 4516
rect 33117 4325 33203 4411
rect 29013 3968 29099 3991
rect 29013 3928 29068 3968
rect 29068 3928 29099 3968
rect 29013 3905 29099 3928
rect 3745 3800 3831 3823
rect 3913 3800 3999 3823
rect 3745 3760 3770 3800
rect 3770 3760 3810 3800
rect 3810 3760 3831 3800
rect 3913 3760 3934 3800
rect 3934 3760 3974 3800
rect 3974 3760 3999 3800
rect 3745 3737 3831 3760
rect 3913 3737 3999 3760
rect 18865 3800 18951 3823
rect 19033 3800 19119 3823
rect 18865 3760 18890 3800
rect 18890 3760 18930 3800
rect 18930 3760 18951 3800
rect 19033 3760 19054 3800
rect 19054 3760 19094 3800
rect 19094 3760 19119 3800
rect 18865 3737 18951 3760
rect 19033 3737 19119 3760
rect 33985 3800 34071 3823
rect 34153 3800 34239 3823
rect 49105 3800 49191 3823
rect 49273 3800 49359 3823
rect 33985 3760 34010 3800
rect 34010 3760 34050 3800
rect 34050 3760 34071 3800
rect 34153 3760 34174 3800
rect 34174 3760 34214 3800
rect 34214 3760 34239 3800
rect 49105 3760 49130 3800
rect 49130 3760 49170 3800
rect 49170 3760 49191 3800
rect 49273 3760 49294 3800
rect 49294 3760 49334 3800
rect 49334 3760 49359 3800
rect 33985 3737 34071 3760
rect 34153 3737 34239 3760
rect 49105 3737 49191 3760
rect 49273 3737 49359 3760
rect 64225 3800 64311 3823
rect 64393 3800 64479 3823
rect 64225 3760 64250 3800
rect 64250 3760 64290 3800
rect 64290 3760 64311 3800
rect 64393 3760 64414 3800
rect 64414 3760 64454 3800
rect 64454 3760 64479 3800
rect 64225 3737 64311 3760
rect 64393 3737 64479 3760
rect 79345 3800 79431 3823
rect 79513 3800 79599 3823
rect 79345 3760 79370 3800
rect 79370 3760 79410 3800
rect 79410 3760 79431 3800
rect 79513 3760 79534 3800
rect 79534 3760 79574 3800
rect 79574 3760 79599 3800
rect 79345 3737 79431 3760
rect 79513 3737 79599 3760
rect 94465 3800 94551 3823
rect 94633 3800 94719 3823
rect 94465 3760 94490 3800
rect 94490 3760 94530 3800
rect 94530 3760 94551 3800
rect 94633 3760 94654 3800
rect 94654 3760 94694 3800
rect 94694 3760 94719 3800
rect 94465 3737 94551 3760
rect 94633 3737 94719 3760
rect 1653 3401 1739 3487
rect 4985 3044 5071 3067
rect 5153 3044 5239 3067
rect 4985 3004 5010 3044
rect 5010 3004 5050 3044
rect 5050 3004 5071 3044
rect 5153 3004 5174 3044
rect 5174 3004 5214 3044
rect 5214 3004 5239 3044
rect 4985 2981 5071 3004
rect 5153 2981 5239 3004
rect 20105 3044 20191 3067
rect 20273 3044 20359 3067
rect 20105 3004 20130 3044
rect 20130 3004 20170 3044
rect 20170 3004 20191 3044
rect 20273 3004 20294 3044
rect 20294 3004 20334 3044
rect 20334 3004 20359 3044
rect 20105 2981 20191 3004
rect 20273 2981 20359 3004
rect 35225 3044 35311 3067
rect 35393 3044 35479 3067
rect 35225 3004 35250 3044
rect 35250 3004 35290 3044
rect 35290 3004 35311 3044
rect 35393 3004 35414 3044
rect 35414 3004 35454 3044
rect 35454 3004 35479 3044
rect 35225 2981 35311 3004
rect 35393 2981 35479 3004
rect 50345 3044 50431 3067
rect 50513 3044 50599 3067
rect 50345 3004 50370 3044
rect 50370 3004 50410 3044
rect 50410 3004 50431 3044
rect 50513 3004 50534 3044
rect 50534 3004 50574 3044
rect 50574 3004 50599 3044
rect 50345 2981 50431 3004
rect 50513 2981 50599 3004
rect 65465 3044 65551 3067
rect 65633 3044 65719 3067
rect 65465 3004 65490 3044
rect 65490 3004 65530 3044
rect 65530 3004 65551 3044
rect 65633 3004 65654 3044
rect 65654 3004 65694 3044
rect 65694 3004 65719 3044
rect 65465 2981 65551 3004
rect 65633 2981 65719 3004
rect 80585 3044 80671 3067
rect 80753 3044 80839 3067
rect 80585 3004 80610 3044
rect 80610 3004 80650 3044
rect 80650 3004 80671 3044
rect 80753 3004 80774 3044
rect 80774 3004 80814 3044
rect 80814 3004 80839 3044
rect 80585 2981 80671 3004
rect 80753 2981 80839 3004
rect 95705 3044 95791 3067
rect 95873 3044 95959 3067
rect 95705 3004 95730 3044
rect 95730 3004 95770 3044
rect 95770 3004 95791 3044
rect 95873 3004 95894 3044
rect 95894 3004 95934 3044
rect 95934 3004 95959 3044
rect 95705 2981 95791 3004
rect 95873 2981 95959 3004
<< metal6 >>
rect 3652 11383 4092 11466
rect 3652 11297 3745 11383
rect 3831 11297 3913 11383
rect 3999 11297 4092 11383
rect 3652 9871 4092 11297
rect 3652 9785 3745 9871
rect 3831 9785 3913 9871
rect 3999 9785 4092 9871
rect 3652 8359 4092 9785
rect 3652 8273 3745 8359
rect 3831 8273 3913 8359
rect 3999 8273 4092 8359
rect 3652 6847 4092 8273
rect 3652 6761 3745 6847
rect 3831 6761 3913 6847
rect 3999 6761 4092 6847
rect 3652 5934 4092 6761
rect 3652 5554 3682 5934
rect 4062 5554 4092 5934
rect 3652 5335 4092 5554
rect 3652 5249 3745 5335
rect 3831 5249 3913 5335
rect 3999 5249 4092 5335
rect 1988 4590 2316 4616
rect 3652 3823 4092 5249
rect 3652 3737 3745 3823
rect 3831 3737 3913 3823
rect 3999 3737 4092 3823
rect 1532 3401 1653 3410
rect 1739 3401 1860 3410
rect 1532 3280 1860 3401
rect 3652 2980 4092 3737
rect 4892 10627 5332 11384
rect 4892 10541 4985 10627
rect 5071 10541 5153 10627
rect 5239 10541 5332 10627
rect 4892 9115 5332 10541
rect 4892 9029 4985 9115
rect 5071 9029 5153 9115
rect 5239 9029 5332 9115
rect 4892 7603 5332 9029
rect 4892 7517 4985 7603
rect 5071 7517 5153 7603
rect 5239 7517 5332 7603
rect 4892 7174 5332 7517
rect 4892 6794 4922 7174
rect 5302 6794 5332 7174
rect 4892 6091 5332 6794
rect 4892 6005 4985 6091
rect 5071 6005 5153 6091
rect 5239 6005 5332 6091
rect 4892 4579 5332 6005
rect 4892 4493 4985 4579
rect 5071 4493 5153 4579
rect 5239 4493 5332 4579
rect 4892 3067 5332 4493
rect 4892 2981 4985 3067
rect 5071 2981 5153 3067
rect 5239 2981 5332 3067
rect 4892 2898 5332 2981
rect 18772 11383 19212 11466
rect 18772 11297 18865 11383
rect 18951 11297 19033 11383
rect 19119 11297 19212 11383
rect 18772 9871 19212 11297
rect 18772 9785 18865 9871
rect 18951 9785 19033 9871
rect 19119 9785 19212 9871
rect 18772 8359 19212 9785
rect 18772 8273 18865 8359
rect 18951 8273 19033 8359
rect 19119 8273 19212 8359
rect 18772 6847 19212 8273
rect 18772 6761 18865 6847
rect 18951 6761 19033 6847
rect 19119 6761 19212 6847
rect 18772 5934 19212 6761
rect 18772 5554 18802 5934
rect 19182 5554 19212 5934
rect 18772 5335 19212 5554
rect 18772 5249 18865 5335
rect 18951 5249 19033 5335
rect 19119 5249 19212 5335
rect 18772 3823 19212 5249
rect 18772 3737 18865 3823
rect 18951 3737 19033 3823
rect 19119 3737 19212 3823
rect 18772 2980 19212 3737
rect 20012 10627 20452 11384
rect 20012 10541 20105 10627
rect 20191 10541 20273 10627
rect 20359 10541 20452 10627
rect 20012 9115 20452 10541
rect 20012 9029 20105 9115
rect 20191 9029 20273 9115
rect 20359 9029 20452 9115
rect 20012 7603 20452 9029
rect 20012 7517 20105 7603
rect 20191 7517 20273 7603
rect 20359 7517 20452 7603
rect 20012 7174 20452 7517
rect 20012 6794 20042 7174
rect 20422 6794 20452 7174
rect 20012 6091 20452 6794
rect 20012 6005 20105 6091
rect 20191 6005 20273 6091
rect 20359 6005 20452 6091
rect 20012 4579 20452 6005
rect 33892 11383 34332 11466
rect 33892 11297 33985 11383
rect 34071 11297 34153 11383
rect 34239 11297 34332 11383
rect 33892 9871 34332 11297
rect 33892 9785 33985 9871
rect 34071 9785 34153 9871
rect 34239 9785 34332 9871
rect 33892 8359 34332 9785
rect 33892 8273 33985 8359
rect 34071 8273 34153 8359
rect 34239 8273 34332 8359
rect 33892 6847 34332 8273
rect 33892 6761 33985 6847
rect 34071 6761 34153 6847
rect 34239 6761 34332 6847
rect 33892 5934 34332 6761
rect 33892 5554 33922 5934
rect 34302 5554 34332 5934
rect 33892 5335 34332 5554
rect 33892 5249 33985 5335
rect 34071 5249 34153 5335
rect 34239 5249 34332 5335
rect 20012 4493 20105 4579
rect 20191 4493 20273 4579
rect 20359 4493 20452 4579
rect 20012 3067 20452 4493
rect 32996 4204 33324 4210
rect 28892 3991 29220 4112
rect 28892 3905 29013 3991
rect 29099 3905 29220 3991
rect 28892 3790 29220 3905
rect 33892 3823 34332 5249
rect 33892 3737 33985 3823
rect 34071 3737 34153 3823
rect 34239 3737 34332 3823
rect 20012 2981 20105 3067
rect 20191 2981 20273 3067
rect 20359 2981 20452 3067
rect 20012 2898 20452 2981
rect 33892 2980 34332 3737
rect 35132 10627 35572 11384
rect 35132 10541 35225 10627
rect 35311 10541 35393 10627
rect 35479 10541 35572 10627
rect 35132 9115 35572 10541
rect 35132 9029 35225 9115
rect 35311 9029 35393 9115
rect 35479 9029 35572 9115
rect 35132 7603 35572 9029
rect 35132 7517 35225 7603
rect 35311 7517 35393 7603
rect 35479 7517 35572 7603
rect 35132 7174 35572 7517
rect 35132 6794 35162 7174
rect 35542 6794 35572 7174
rect 35132 6091 35572 6794
rect 35132 6005 35225 6091
rect 35311 6005 35393 6091
rect 35479 6005 35572 6091
rect 35132 4579 35572 6005
rect 35132 4493 35225 4579
rect 35311 4493 35393 4579
rect 35479 4493 35572 4579
rect 35132 3067 35572 4493
rect 35132 2981 35225 3067
rect 35311 2981 35393 3067
rect 35479 2981 35572 3067
rect 35132 2898 35572 2981
rect 49012 11383 49452 11466
rect 49012 11297 49105 11383
rect 49191 11297 49273 11383
rect 49359 11297 49452 11383
rect 49012 9871 49452 11297
rect 49012 9785 49105 9871
rect 49191 9785 49273 9871
rect 49359 9785 49452 9871
rect 49012 8359 49452 9785
rect 49012 8273 49105 8359
rect 49191 8273 49273 8359
rect 49359 8273 49452 8359
rect 49012 6847 49452 8273
rect 49012 6761 49105 6847
rect 49191 6761 49273 6847
rect 49359 6761 49452 6847
rect 49012 5934 49452 6761
rect 49012 5554 49042 5934
rect 49422 5554 49452 5934
rect 49012 5335 49452 5554
rect 49012 5249 49105 5335
rect 49191 5249 49273 5335
rect 49359 5249 49452 5335
rect 49012 3823 49452 5249
rect 49012 3737 49105 3823
rect 49191 3737 49273 3823
rect 49359 3737 49452 3823
rect 49012 2980 49452 3737
rect 50252 10627 50692 11384
rect 50252 10541 50345 10627
rect 50431 10541 50513 10627
rect 50599 10541 50692 10627
rect 50252 9115 50692 10541
rect 50252 9029 50345 9115
rect 50431 9029 50513 9115
rect 50599 9029 50692 9115
rect 50252 7603 50692 9029
rect 50252 7517 50345 7603
rect 50431 7517 50513 7603
rect 50599 7517 50692 7603
rect 50252 7174 50692 7517
rect 50252 6794 50282 7174
rect 50662 6794 50692 7174
rect 50252 6091 50692 6794
rect 50252 6005 50345 6091
rect 50431 6005 50513 6091
rect 50599 6005 50692 6091
rect 50252 4579 50692 6005
rect 50252 4493 50345 4579
rect 50431 4493 50513 4579
rect 50599 4493 50692 4579
rect 50252 3067 50692 4493
rect 50252 2981 50345 3067
rect 50431 2981 50513 3067
rect 50599 2981 50692 3067
rect 50252 2898 50692 2981
rect 64132 11383 64572 11466
rect 64132 11297 64225 11383
rect 64311 11297 64393 11383
rect 64479 11297 64572 11383
rect 64132 9871 64572 11297
rect 64132 9785 64225 9871
rect 64311 9785 64393 9871
rect 64479 9785 64572 9871
rect 64132 8359 64572 9785
rect 64132 8273 64225 8359
rect 64311 8273 64393 8359
rect 64479 8273 64572 8359
rect 64132 6847 64572 8273
rect 64132 6761 64225 6847
rect 64311 6761 64393 6847
rect 64479 6761 64572 6847
rect 64132 5934 64572 6761
rect 64132 5554 64162 5934
rect 64542 5554 64572 5934
rect 64132 5335 64572 5554
rect 64132 5249 64225 5335
rect 64311 5249 64393 5335
rect 64479 5249 64572 5335
rect 64132 3823 64572 5249
rect 64132 3737 64225 3823
rect 64311 3737 64393 3823
rect 64479 3737 64572 3823
rect 64132 2980 64572 3737
rect 65372 10627 65812 11384
rect 65372 10541 65465 10627
rect 65551 10541 65633 10627
rect 65719 10541 65812 10627
rect 65372 9115 65812 10541
rect 65372 9029 65465 9115
rect 65551 9029 65633 9115
rect 65719 9029 65812 9115
rect 65372 7603 65812 9029
rect 65372 7517 65465 7603
rect 65551 7517 65633 7603
rect 65719 7517 65812 7603
rect 65372 7174 65812 7517
rect 65372 6794 65402 7174
rect 65782 6794 65812 7174
rect 65372 6091 65812 6794
rect 65372 6005 65465 6091
rect 65551 6005 65633 6091
rect 65719 6005 65812 6091
rect 65372 4579 65812 6005
rect 65372 4493 65465 4579
rect 65551 4493 65633 4579
rect 65719 4493 65812 4579
rect 65372 3067 65812 4493
rect 65372 2981 65465 3067
rect 65551 2981 65633 3067
rect 65719 2981 65812 3067
rect 65372 2898 65812 2981
rect 79252 11383 79692 11466
rect 79252 11297 79345 11383
rect 79431 11297 79513 11383
rect 79599 11297 79692 11383
rect 79252 9871 79692 11297
rect 79252 9785 79345 9871
rect 79431 9785 79513 9871
rect 79599 9785 79692 9871
rect 79252 8359 79692 9785
rect 79252 8273 79345 8359
rect 79431 8273 79513 8359
rect 79599 8273 79692 8359
rect 79252 6847 79692 8273
rect 79252 6761 79345 6847
rect 79431 6761 79513 6847
rect 79599 6761 79692 6847
rect 79252 5934 79692 6761
rect 79252 5554 79282 5934
rect 79662 5554 79692 5934
rect 79252 5335 79692 5554
rect 79252 5249 79345 5335
rect 79431 5249 79513 5335
rect 79599 5249 79692 5335
rect 79252 3823 79692 5249
rect 79252 3737 79345 3823
rect 79431 3737 79513 3823
rect 79599 3737 79692 3823
rect 79252 2980 79692 3737
rect 80492 10627 80932 11384
rect 80492 10541 80585 10627
rect 80671 10541 80753 10627
rect 80839 10541 80932 10627
rect 80492 9115 80932 10541
rect 80492 9029 80585 9115
rect 80671 9029 80753 9115
rect 80839 9029 80932 9115
rect 80492 7603 80932 9029
rect 80492 7517 80585 7603
rect 80671 7517 80753 7603
rect 80839 7517 80932 7603
rect 80492 7174 80932 7517
rect 80492 6794 80522 7174
rect 80902 6794 80932 7174
rect 80492 6091 80932 6794
rect 80492 6005 80585 6091
rect 80671 6005 80753 6091
rect 80839 6005 80932 6091
rect 80492 4579 80932 6005
rect 80492 4493 80585 4579
rect 80671 4493 80753 4579
rect 80839 4493 80932 4579
rect 80492 3067 80932 4493
rect 80492 2981 80585 3067
rect 80671 2981 80753 3067
rect 80839 2981 80932 3067
rect 80492 2898 80932 2981
rect 94372 11383 94812 11466
rect 94372 11297 94465 11383
rect 94551 11297 94633 11383
rect 94719 11297 94812 11383
rect 94372 9871 94812 11297
rect 94372 9785 94465 9871
rect 94551 9785 94633 9871
rect 94719 9785 94812 9871
rect 94372 8359 94812 9785
rect 94372 8273 94465 8359
rect 94551 8273 94633 8359
rect 94719 8273 94812 8359
rect 94372 6847 94812 8273
rect 94372 6761 94465 6847
rect 94551 6761 94633 6847
rect 94719 6761 94812 6847
rect 94372 5934 94812 6761
rect 94372 5554 94402 5934
rect 94782 5554 94812 5934
rect 94372 5335 94812 5554
rect 94372 5249 94465 5335
rect 94551 5249 94633 5335
rect 94719 5249 94812 5335
rect 94372 3823 94812 5249
rect 94372 3737 94465 3823
rect 94551 3737 94633 3823
rect 94719 3737 94812 3823
rect 94372 2980 94812 3737
rect 95612 10627 96052 11384
rect 95612 10541 95705 10627
rect 95791 10541 95873 10627
rect 95959 10541 96052 10627
rect 95612 9115 96052 10541
rect 95612 9029 95705 9115
rect 95791 9029 95873 9115
rect 95959 9029 96052 9115
rect 95612 7603 96052 9029
rect 95612 7517 95705 7603
rect 95791 7517 95873 7603
rect 95959 7517 96052 7603
rect 95612 7174 96052 7517
rect 95612 6794 95642 7174
rect 96022 6794 96052 7174
rect 95612 6091 96052 6794
rect 95612 6005 95705 6091
rect 95791 6005 95873 6091
rect 95959 6005 96052 6091
rect 95612 4579 96052 6005
rect 95612 4493 95705 4579
rect 95791 4493 95873 4579
rect 95959 4493 96052 4579
rect 95612 3067 96052 4493
rect 95612 2981 95705 3067
rect 95791 2981 95873 3067
rect 95959 2981 96052 3067
rect 95612 2898 96052 2981
<< via6 >>
rect 3682 5554 4062 5934
rect 1962 4495 2342 4590
rect 1962 4409 2109 4495
rect 2109 4409 2195 4495
rect 2195 4409 2342 4495
rect 1962 4210 2342 4409
rect 1506 3487 1886 3790
rect 1506 3410 1653 3487
rect 1653 3410 1739 3487
rect 1739 3410 1886 3487
rect 4922 6794 5302 7174
rect 18802 5554 19182 5934
rect 20042 6794 20422 7174
rect 33922 5554 34302 5934
rect 32970 4411 33350 4590
rect 32970 4325 33117 4411
rect 33117 4325 33203 4411
rect 33203 4325 33350 4411
rect 32970 4210 33350 4325
rect 28866 3410 29246 3790
rect 35162 6794 35542 7174
rect 49042 5554 49422 5934
rect 50282 6794 50662 7174
rect 64162 5554 64542 5934
rect 65402 6794 65782 7174
rect 79282 5554 79662 5934
rect 80522 6794 80902 7174
rect 94402 5554 94782 5934
rect 95642 6794 96022 7174
<< metal7 >>
rect 1108 7174 98828 7204
rect 1108 6794 4922 7174
rect 5302 6794 20042 7174
rect 20422 6794 35162 7174
rect 35542 6794 50282 7174
rect 50662 6794 65402 7174
rect 65782 6794 80522 7174
rect 80902 6794 95642 7174
rect 96022 6794 98828 7174
rect 1108 6764 98828 6794
rect 1108 5934 98828 5964
rect 1108 5554 3682 5934
rect 4062 5554 18802 5934
rect 19182 5554 33922 5934
rect 34302 5554 49042 5934
rect 49422 5554 64162 5934
rect 64542 5554 79282 5934
rect 79662 5554 94402 5934
rect 94782 5554 98828 5934
rect 1108 5524 98828 5554
rect 1952 4590 33360 4600
rect 1952 4210 1962 4590
rect 2342 4210 32970 4590
rect 33350 4210 33360 4590
rect 1952 4200 33360 4210
rect 1496 3790 29256 3800
rect 1496 3410 1506 3790
rect 1886 3410 28866 3790
rect 29246 3410 29256 3790
rect 1496 3400 29256 3410
use sg13g2_inv_1  _095_
timestamp 1676382929
transform 1 0 37152 0 -1 6048
box -48 -56 336 834
use sg13g2_nor2_1  _096_
timestamp 1676627187
transform 1 0 51168 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _097_
timestamp 1676627187
transform -1 0 49824 0 -1 7560
box -48 -56 432 834
use sg13g2_nor4_2  _098_
timestamp 1685199459
transform 1 0 49920 0 -1 7560
box -48 -56 1200 834
use sg13g2_nor2b_2  _099_
timestamp 1685188981
transform -1 0 60864 0 1 6048
box -54 -56 720 834
use sg13g2_and4_1  _100_
timestamp 1676985977
transform 1 0 61632 0 1 6048
box -48 -56 816 834
use sg13g2_nand4_1  _101_
timestamp 1685201930
transform 1 0 60192 0 -1 7560
box -48 -56 624 834
use sg13g2_and2_1  _102_
timestamp 1676901763
transform -1 0 62880 0 1 6048
box -48 -56 528 834
use sg13g2_nand2_1  _103_
timestamp 1676557249
transform -1 0 63264 0 1 6048
box -48 -56 432 834
use sg13g2_and2_1  _104_
timestamp 1676901763
transform -1 0 50592 0 1 6048
box -48 -56 528 834
use sg13g2_and2_1  _105_
timestamp 1676901763
transform 1 0 49824 0 -1 9072
box -48 -56 528 834
use sg13g2_nand2_2  _106_
timestamp 1685180049
transform 1 0 51360 0 -1 4536
box -48 -56 624 834
use sg13g2_nor2b_2  _107_
timestamp 1685188981
transform -1 0 77376 0 1 6048
box -54 -56 720 834
use sg13g2_and3_1  _108_
timestamp 1676971669
transform -1 0 61632 0 -1 6048
box -48 -56 720 834
use sg13g2_nand3_1  _109_
timestamp 1683988354
transform -1 0 60192 0 -1 7560
box -48 -56 528 834
use sg13g2_nor2_1  _110_
timestamp 1676627187
transform -1 0 55392 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2b_1  _111_
timestamp 1676567195
transform 1 0 60864 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2b_2  _112_
timestamp 1685188981
transform 1 0 49728 0 1 7560
box -54 -56 720 834
use sg13g2_nand2_1  _113_
timestamp 1676557249
transform 1 0 49440 0 1 4536
box -48 -56 432 834
use sg13g2_nor2_1  _114_
timestamp 1676627187
transform 1 0 48960 0 -1 4536
box -48 -56 432 834
use sg13g2_or2_1  _115_
timestamp 1684236171
transform 1 0 49344 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2b_2  _116_
timestamp 1685188981
transform -1 0 49728 0 1 7560
box -54 -56 720 834
use sg13g2_nand2_1  _117_
timestamp 1676557249
transform -1 0 50208 0 1 4536
box -48 -56 432 834
use sg13g2_nor2_1  _118_
timestamp 1676627187
transform 1 0 49056 0 1 3024
box -48 -56 432 834
use sg13g2_or2_1  _119_
timestamp 1684236171
transform 1 0 49440 0 1 3024
box -48 -56 528 834
use sg13g2_nand2_1  _120_
timestamp 1676557249
transform 1 0 51936 0 -1 4536
box -48 -56 432 834
use sg13g2_nor2_1  _121_
timestamp 1676627187
transform -1 0 53664 0 -1 4536
box -48 -56 432 834
use sg13g2_or2_1  _122_
timestamp 1684236171
transform 1 0 52800 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2b_1  _123_
timestamp 1685181386
transform -1 0 51648 0 -1 7560
box -54 -56 528 834
use sg13g2_nand2_1  _124_
timestamp 1676557249
transform -1 0 54624 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _125_
timestamp 1676627187
transform 1 0 53664 0 -1 6048
box -48 -56 432 834
use sg13g2_or2_1  _126_
timestamp 1684236171
transform 1 0 54240 0 1 6048
box -48 -56 528 834
use sg13g2_nand2_1  _127_
timestamp 1676557249
transform 1 0 55872 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _128_
timestamp 1676627187
transform 1 0 56736 0 1 7560
box -48 -56 432 834
use sg13g2_or2_1  _129_
timestamp 1684236171
transform 1 0 57024 0 -1 9072
box -48 -56 528 834
use sg13g2_nand2_1  _130_
timestamp 1676557249
transform -1 0 55104 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _131_
timestamp 1676627187
transform 1 0 54720 0 1 7560
box -48 -56 432 834
use sg13g2_or2_1  _132_
timestamp 1684236171
transform 1 0 55104 0 -1 9072
box -48 -56 528 834
use sg13g2_nand2_1  _133_
timestamp 1676557249
transform 1 0 55968 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _134_
timestamp 1676627187
transform 1 0 57600 0 1 7560
box -48 -56 432 834
use sg13g2_or2_1  _135_
timestamp 1684236171
transform 1 0 58176 0 -1 7560
box -48 -56 528 834
use sg13g2_nor2b_1  _136_
timestamp 1685181386
transform 1 0 51552 0 1 6048
box -54 -56 528 834
use sg13g2_nand2_1  _137_
timestamp 1676557249
transform 1 0 55968 0 1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _138_
timestamp 1676627187
transform 1 0 56448 0 1 6048
box -48 -56 432 834
use sg13g2_or2_1  _139_
timestamp 1684236171
transform 1 0 56832 0 1 6048
box -48 -56 528 834
use sg13g2_nand2_1  _140_
timestamp 1676557249
transform 1 0 55584 0 -1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _141_
timestamp 1676627187
transform 1 0 56640 0 -1 6048
box -48 -56 432 834
use sg13g2_or2_1  _142_
timestamp 1684236171
transform 1 0 57504 0 -1 6048
box -48 -56 528 834
use sg13g2_nand2_1  _143_
timestamp 1676557249
transform 1 0 55872 0 1 4536
box -48 -56 432 834
use sg13g2_nor2_1  _144_
timestamp 1676627187
transform 1 0 57408 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _145_
timestamp 1684236171
transform 1 0 56352 0 -1 4536
box -48 -56 528 834
use sg13g2_nand2_1  _146_
timestamp 1676557249
transform 1 0 56256 0 1 4536
box -48 -56 432 834
use sg13g2_nor2_1  _147_
timestamp 1676627187
transform 1 0 56256 0 -1 6048
box -48 -56 432 834
use sg13g2_or2_1  _148_
timestamp 1684236171
transform 1 0 56832 0 -1 4536
box -48 -56 528 834
use sg13g2_nand2_1  _149_
timestamp 1676557249
transform 1 0 55680 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _150_
timestamp 1676627187
transform 1 0 60192 0 -1 10584
box -48 -56 432 834
use sg13g2_or2_1  _151_
timestamp 1684236171
transform 1 0 60672 0 1 9072
box -48 -56 528 834
use sg13g2_nand2_1  _152_
timestamp 1676557249
transform 1 0 56448 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _153_
timestamp 1676627187
transform -1 0 59712 0 1 9072
box -48 -56 432 834
use sg13g2_or2_1  _154_
timestamp 1684236171
transform 1 0 59712 0 1 9072
box -48 -56 528 834
use sg13g2_nand2_1  _155_
timestamp 1676557249
transform 1 0 56064 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _156_
timestamp 1676627187
transform 1 0 59808 0 -1 10584
box -48 -56 432 834
use sg13g2_or2_1  _157_
timestamp 1684236171
transform 1 0 60192 0 1 9072
box -48 -56 528 834
use sg13g2_and2_1  _158_
timestamp 1676901763
transform 1 0 61152 0 1 4536
box -48 -56 528 834
use sg13g2_nand2_1  _159_
timestamp 1676557249
transform 1 0 61632 0 1 4536
box -48 -56 432 834
use sg13g2_nor2b_2  _160_
timestamp 1685188981
transform -1 0 71616 0 1 6048
box -54 -56 720 834
use sg13g2_and2_1  _161_
timestamp 1676901763
transform -1 0 72960 0 1 7560
box -48 -56 528 834
use sg13g2_nand2_1  _162_
timestamp 1676557249
transform 1 0 67104 0 1 6048
box -48 -56 432 834
use sg13g2_and3_2  _163_
timestamp 1683976310
transform -1 0 45504 0 -1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _164_
timestamp 1683988354
transform -1 0 44928 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _165_
timestamp 1676627187
transform -1 0 67872 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _166_
timestamp 1676557249
transform 1 0 69696 0 1 7560
box -48 -56 432 834
use sg13g2_and3_2  _167_
timestamp 1683976310
transform -1 0 44640 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _168_
timestamp 1683988354
transform 1 0 45024 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _169_
timestamp 1676627187
transform -1 0 68448 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _170_
timestamp 1676557249
transform -1 0 70464 0 1 7560
box -48 -56 432 834
use sg13g2_and3_2  _171_
timestamp 1683976310
transform 1 0 44640 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _172_
timestamp 1683988354
transform -1 0 46272 0 1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _173_
timestamp 1676627187
transform -1 0 67488 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _174_
timestamp 1676557249
transform -1 0 70272 0 -1 9072
box -48 -56 432 834
use sg13g2_and3_2  _175_
timestamp 1683976310
transform -1 0 44928 0 -1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _176_
timestamp 1683988354
transform -1 0 44448 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _177_
timestamp 1676627187
transform -1 0 68064 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _178_
timestamp 1676557249
transform -1 0 70848 0 -1 7560
box -48 -56 432 834
use sg13g2_and3_2  _179_
timestamp 1683976310
transform -1 0 47520 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _180_
timestamp 1683988354
transform 1 0 47424 0 1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _181_
timestamp 1676627187
transform -1 0 68256 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _182_
timestamp 1676557249
transform -1 0 70848 0 1 7560
box -48 -56 432 834
use sg13g2_and3_2  _183_
timestamp 1683976310
transform -1 0 46848 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _184_
timestamp 1683988354
transform -1 0 46464 0 1 3024
box -48 -56 528 834
use sg13g2_nor2_1  _185_
timestamp 1676627187
transform -1 0 68832 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _186_
timestamp 1676557249
transform -1 0 70752 0 -1 9072
box -48 -56 432 834
use sg13g2_and3_2  _187_
timestamp 1683976310
transform -1 0 46176 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _188_
timestamp 1683988354
transform 1 0 46464 0 1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _189_
timestamp 1676627187
transform -1 0 68640 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _190_
timestamp 1676557249
transform -1 0 71232 0 1 7560
box -48 -56 432 834
use sg13g2_and3_2  _191_
timestamp 1683976310
transform -1 0 46944 0 -1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _192_
timestamp 1683988354
transform 1 0 46944 0 1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _193_
timestamp 1676627187
transform 1 0 68832 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _194_
timestamp 1676557249
transform -1 0 71136 0 -1 9072
box -48 -56 432 834
use sg13g2_and3_2  _195_
timestamp 1683976310
transform 1 0 49056 0 -1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _196_
timestamp 1683988354
transform -1 0 49440 0 -1 7560
box -48 -56 528 834
use sg13g2_nor2_1  _197_
timestamp 1676627187
transform -1 0 68640 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _198_
timestamp 1676557249
transform -1 0 72288 0 1 9072
box -48 -56 432 834
use sg13g2_and3_2  _199_
timestamp 1683976310
transform 1 0 49248 0 1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _200_
timestamp 1683988354
transform -1 0 52608 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _201_
timestamp 1676627187
transform -1 0 68832 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _202_
timestamp 1676557249
transform -1 0 73440 0 1 9072
box -48 -56 432 834
use sg13g2_and3_2  _203_
timestamp 1683976310
transform -1 0 49248 0 1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _204_
timestamp 1683988354
transform -1 0 52992 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _205_
timestamp 1676627187
transform -1 0 69408 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _206_
timestamp 1676557249
transform -1 0 73248 0 -1 10584
box -48 -56 432 834
use sg13g2_and3_2  _207_
timestamp 1683976310
transform -1 0 48768 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _208_
timestamp 1683988354
transform -1 0 48288 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _209_
timestamp 1676627187
transform -1 0 68352 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _210_
timestamp 1676557249
transform -1 0 71904 0 1 9072
box -48 -56 432 834
use sg13g2_and3_2  _211_
timestamp 1683976310
transform -1 0 51744 0 1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _212_
timestamp 1683988354
transform 1 0 51072 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _213_
timestamp 1676627187
transform 1 0 69408 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _214_
timestamp 1676557249
transform 1 0 71232 0 -1 10584
box -48 -56 432 834
use sg13g2_and3_2  _215_
timestamp 1683976310
transform 1 0 52320 0 -1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _216_
timestamp 1683988354
transform -1 0 52512 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _217_
timestamp 1676627187
transform 1 0 67968 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _218_
timestamp 1676557249
transform -1 0 74592 0 -1 10584
box -48 -56 432 834
use sg13g2_and3_2  _219_
timestamp 1683976310
transform 1 0 51744 0 1 9072
box -48 -56 720 834
use sg13g2_nand3_1  _220_
timestamp 1683988354
transform 1 0 51648 0 -1 7560
box -48 -56 528 834
use sg13g2_nor2_1  _221_
timestamp 1676627187
transform -1 0 69312 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _222_
timestamp 1676557249
transform -1 0 74016 0 1 9072
box -48 -56 432 834
use sg13g2_and2_1  _223_
timestamp 1676901763
transform 1 0 61728 0 -1 7560
box -48 -56 528 834
use sg13g2_nand2_2  _224_
timestamp 1685180049
transform -1 0 62208 0 -1 6048
box -48 -56 624 834
use sg13g2_nor2_1  _225_
timestamp 1676627187
transform 1 0 68640 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _226_
timestamp 1676557249
transform -1 0 73536 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_2  _227_
timestamp 1683979924
transform 1 0 71616 0 1 6048
box -48 -56 624 834
use sg13g2_and2_1  _228_
timestamp 1676901763
transform 1 0 74688 0 1 7560
box -48 -56 528 834
use sg13g2_nand2_1  _229_
timestamp 1676557249
transform 1 0 72576 0 1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _230_
timestamp 1676627187
transform 1 0 69888 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _231_
timestamp 1676557249
transform -1 0 75552 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _232_
timestamp 1676627187
transform -1 0 70752 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _233_
timestamp 1676557249
transform 1 0 75648 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _234_
timestamp 1676627187
transform 1 0 69984 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _235_
timestamp 1676557249
transform -1 0 75648 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _236_
timestamp 1676627187
transform 1 0 69504 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _237_
timestamp 1676557249
transform -1 0 74304 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _238_
timestamp 1676627187
transform -1 0 71136 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _239_
timestamp 1676557249
transform -1 0 74688 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _240_
timestamp 1676627187
transform 1 0 70272 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _241_
timestamp 1676557249
transform -1 0 74880 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _242_
timestamp 1676627187
transform -1 0 71520 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _243_
timestamp 1676557249
transform -1 0 75264 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _244_
timestamp 1676627187
transform 1 0 69504 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _245_
timestamp 1676557249
transform -1 0 75168 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _246_
timestamp 1676627187
transform -1 0 75072 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _247_
timestamp 1676557249
transform 1 0 77664 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _248_
timestamp 1676627187
transform 1 0 74112 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _249_
timestamp 1676557249
transform -1 0 77664 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _250_
timestamp 1676627187
transform -1 0 74688 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _251_
timestamp 1676557249
transform -1 0 76800 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _252_
timestamp 1676627187
transform 1 0 74208 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _253_
timestamp 1676557249
transform -1 0 77280 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _254_
timestamp 1676627187
transform 1 0 73920 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _255_
timestamp 1676557249
transform -1 0 77952 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _256_
timestamp 1676627187
transform -1 0 75456 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _257_
timestamp 1676557249
transform -1 0 77568 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _258_
timestamp 1676627187
transform 1 0 73728 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _259_
timestamp 1676557249
transform 1 0 76800 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _260_
timestamp 1676627187
transform 1 0 73344 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _261_
timestamp 1676557249
transform 1 0 76608 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_2  _262_
timestamp 1683979924
transform 1 0 60864 0 1 6048
box -48 -56 624 834
use sg13g2_and3_2  _263_
timestamp 1683976310
transform 1 0 76992 0 -1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _264_
timestamp 1683988354
transform -1 0 77856 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _265_
timestamp 1676627187
transform 1 0 73440 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _266_
timestamp 1676557249
transform -1 0 78336 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _267_
timestamp 1676627187
transform 1 0 72288 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _268_
timestamp 1676557249
transform -1 0 78240 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _269_
timestamp 1676627187
transform 1 0 71904 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _270_
timestamp 1676557249
transform -1 0 79008 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _271_
timestamp 1676627187
transform 1 0 72672 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _272_
timestamp 1676557249
transform -1 0 77856 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _273_
timestamp 1676627187
transform -1 0 79104 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _274_
timestamp 1676557249
transform -1 0 78624 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _275_
timestamp 1676627187
transform 1 0 75744 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _276_
timestamp 1676557249
transform 1 0 78240 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _277_
timestamp 1676627187
transform 1 0 75648 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _278_
timestamp 1676557249
transform 1 0 77856 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _279_
timestamp 1676627187
transform 1 0 72672 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _280_
timestamp 1676557249
transform 1 0 78720 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _281_
timestamp 1676627187
transform 1 0 79008 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _282_
timestamp 1676557249
transform -1 0 80928 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _283_
timestamp 1676627187
transform 1 0 79200 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _284_
timestamp 1676557249
transform -1 0 82176 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _285_
timestamp 1676627187
transform 1 0 78624 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _286_
timestamp 1676557249
transform -1 0 82848 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _287_
timestamp 1676627187
transform 1 0 78816 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _288_
timestamp 1676557249
transform 1 0 80928 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _289_
timestamp 1676627187
transform 1 0 79200 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _290_
timestamp 1676557249
transform -1 0 84288 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _291_
timestamp 1676627187
transform 1 0 79584 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _292_
timestamp 1676557249
transform -1 0 83904 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _293_
timestamp 1676627187
transform 1 0 78432 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _294_
timestamp 1676557249
transform -1 0 83520 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _295_
timestamp 1676627187
transform -1 0 80352 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _296_
timestamp 1676557249
transform 1 0 84000 0 -1 9072
box -48 -56 432 834
use sg13g2_and2_1  _297_
timestamp 1676901763
transform 1 0 78336 0 -1 7560
box -48 -56 528 834
use sg13g2_nand2_2  _298_
timestamp 1685180049
transform -1 0 78240 0 -1 6048
box -48 -56 624 834
use sg13g2_nor2_1  _299_
timestamp 1676627187
transform 1 0 71904 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _300_
timestamp 1676557249
transform 1 0 80640 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _301_
timestamp 1676627187
transform 1 0 71040 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _302_
timestamp 1676557249
transform 1 0 81024 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _303_
timestamp 1676627187
transform 1 0 71424 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _304_
timestamp 1676557249
transform 1 0 81120 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _305_
timestamp 1676627187
transform 1 0 71520 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _306_
timestamp 1676557249
transform 1 0 81792 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _307_
timestamp 1676627187
transform 1 0 77184 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _308_
timestamp 1676557249
transform 1 0 81888 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _309_
timestamp 1676627187
transform 1 0 73056 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _310_
timestamp 1676557249
transform 1 0 81504 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _311_
timestamp 1676627187
transform 1 0 76128 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _312_
timestamp 1676557249
transform 1 0 80736 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _313_
timestamp 1676627187
transform 1 0 74592 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _314_
timestamp 1676557249
transform 1 0 81408 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _315_
timestamp 1676627187
transform 1 0 83040 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _316_
timestamp 1676557249
transform -1 0 88128 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _317_
timestamp 1676627187
transform 1 0 84864 0 1 3024
box -48 -56 432 834
use sg13g2_nand2_1  _318_
timestamp 1676557249
transform -1 0 87552 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _319_
timestamp 1676627187
transform 1 0 83616 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _320_
timestamp 1676557249
transform -1 0 87456 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _321_
timestamp 1676627187
transform 1 0 80832 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _322_
timestamp 1676557249
transform -1 0 88320 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _323_
timestamp 1676627187
transform 1 0 82464 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _324_
timestamp 1676557249
transform -1 0 88512 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _325_
timestamp 1676627187
transform 1 0 83424 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _326_
timestamp 1676557249
transform -1 0 88896 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _327_
timestamp 1676627187
transform 1 0 85248 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _328_
timestamp 1676557249
transform -1 0 89664 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _329_
timestamp 1676627187
transform 1 0 80736 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _330_
timestamp 1676557249
transform -1 0 88320 0 -1 7560
box -48 -56 432 834
use sg13g2_and2_1  _331_
timestamp 1676901763
transform 1 0 84480 0 1 6048
box -48 -56 528 834
use sg13g2_nand2_2  _332_
timestamp 1685180049
transform -1 0 84768 0 -1 6048
box -48 -56 624 834
use sg13g2_nor2_1  _333_
timestamp 1676627187
transform 1 0 72288 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _334_
timestamp 1676557249
transform 1 0 84096 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _335_
timestamp 1676627187
transform 1 0 73056 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _336_
timestamp 1676557249
transform 1 0 83712 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _337_
timestamp 1676627187
transform 1 0 72672 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _338_
timestamp 1676557249
transform -1 0 82752 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _339_
timestamp 1676627187
transform 1 0 71904 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _340_
timestamp 1676557249
transform 1 0 83040 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _341_
timestamp 1676627187
transform 1 0 80640 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _342_
timestamp 1676557249
transform 1 0 83424 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _343_
timestamp 1676627187
transform 1 0 76512 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _344_
timestamp 1676557249
transform -1 0 83904 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _345_
timestamp 1676627187
transform 1 0 76896 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _346_
timestamp 1676557249
transform 1 0 83136 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _347_
timestamp 1676627187
transform 1 0 75744 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _348_
timestamp 1676557249
transform -1 0 88896 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _349_
timestamp 1676627187
transform 1 0 83232 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _350_
timestamp 1676557249
transform 1 0 89376 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _351_
timestamp 1676627187
transform 1 0 82656 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _352_
timestamp 1676557249
transform 1 0 89280 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _353_
timestamp 1676627187
transform 1 0 82848 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _354_
timestamp 1676557249
transform 1 0 89376 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _355_
timestamp 1676627187
transform 1 0 81216 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _356_
timestamp 1676557249
transform -1 0 87936 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _357_
timestamp 1676627187
transform 1 0 82080 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _358_
timestamp 1676557249
transform -1 0 88896 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _359_
timestamp 1676627187
transform 1 0 83808 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _360_
timestamp 1676557249
transform 1 0 88128 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _361_
timestamp 1676627187
transform 1 0 82560 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _362_
timestamp 1676557249
transform 1 0 88896 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _363_
timestamp 1676627187
transform 1 0 81504 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _364_
timestamp 1676557249
transform 1 0 86592 0 1 6048
box -48 -56 432 834
use sg13g2_and2_1  _365_
timestamp 1676901763
transform 1 0 78816 0 -1 7560
box -48 -56 528 834
use sg13g2_nand2_2  _366_
timestamp 1685180049
transform -1 0 75264 0 -1 6048
box -48 -56 624 834
use sg13g2_nor2_2  _367_
timestamp 1683979924
transform 1 0 59904 0 1 3024
box -48 -56 624 834
use sg13g2_nand2_1  _368_
timestamp 1676557249
transform -1 0 85440 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _369_
timestamp 1683979924
transform 1 0 59328 0 1 3024
box -48 -56 624 834
use sg13g2_nand2_1  _370_
timestamp 1676557249
transform -1 0 85056 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _371_
timestamp 1683979924
transform 1 0 64416 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _372_
timestamp 1676557249
transform -1 0 83136 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _373_
timestamp 1683979924
transform 1 0 66720 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _374_
timestamp 1676557249
transform 1 0 82944 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _375_
timestamp 1676627187
transform 1 0 81120 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _376_
timestamp 1676557249
transform -1 0 84672 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _377_
timestamp 1683979924
transform -1 0 60864 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _378_
timestamp 1676557249
transform 1 0 83328 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _379_
timestamp 1676627187
transform 1 0 76512 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _380_
timestamp 1676557249
transform -1 0 84288 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _381_
timestamp 1683979924
transform 1 0 59520 0 1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _382_
timestamp 1676557249
transform 1 0 88128 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _383_
timestamp 1676627187
transform 1 0 82656 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _384_
timestamp 1676557249
transform 1 0 88992 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _385_
timestamp 1676627187
transform 1 0 83136 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _386_
timestamp 1676557249
transform 1 0 88896 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _387_
timestamp 1676627187
transform 1 0 82080 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _388_
timestamp 1676557249
transform 1 0 89664 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _389_
timestamp 1676627187
transform 1 0 80352 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _390_
timestamp 1676557249
transform -1 0 87168 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _391_
timestamp 1676627187
transform 1 0 81600 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _392_
timestamp 1676557249
transform 1 0 87648 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _393_
timestamp 1676627187
transform 1 0 83232 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _394_
timestamp 1676557249
transform 1 0 87744 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _395_
timestamp 1676627187
transform -1 0 84000 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _396_
timestamp 1676557249
transform 1 0 88896 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_2  _397_
timestamp 1683979924
transform 1 0 74112 0 -1 6048
box -48 -56 624 834
use sg13g2_nand2_1  _398_
timestamp 1676557249
transform 1 0 85536 0 -1 7560
box -48 -56 432 834
use sg13g2_and3_2  _399_
timestamp 1683976310
transform -1 0 23328 0 -1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _400_
timestamp 1683988354
transform -1 0 23424 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _401_
timestamp 1676627187
transform -1 0 22176 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _402_
timestamp 1676557249
transform -1 0 9984 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _403_
timestamp 1676627187
transform -1 0 21792 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _404_
timestamp 1676557249
transform -1 0 11328 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _405_
timestamp 1676627187
transform -1 0 22176 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _406_
timestamp 1676557249
transform -1 0 10752 0 1 6048
box -48 -56 432 834
use sg13g2_nor2_1  _407_
timestamp 1676627187
transform -1 0 22560 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _408_
timestamp 1676557249
transform -1 0 10944 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _409_
timestamp 1676627187
transform -1 0 21024 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _410_
timestamp 1676557249
transform -1 0 11904 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _411_
timestamp 1676627187
transform -1 0 17664 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _412_
timestamp 1676557249
transform -1 0 12672 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _413_
timestamp 1676627187
transform -1 0 18912 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _414_
timestamp 1676557249
transform -1 0 12192 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _415_
timestamp 1676627187
transform -1 0 17472 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _416_
timestamp 1676557249
transform -1 0 12864 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _417_
timestamp 1676627187
transform -1 0 16416 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _418_
timestamp 1676557249
transform 1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _419_
timestamp 1676627187
transform -1 0 16032 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _420_
timestamp 1676557249
transform 1 0 15264 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _421_
timestamp 1676627187
transform -1 0 17184 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _422_
timestamp 1676557249
transform 1 0 14880 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _423_
timestamp 1676627187
transform -1 0 20832 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _424_
timestamp 1676557249
transform 1 0 15552 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _425_
timestamp 1676627187
transform -1 0 19296 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _426_
timestamp 1676557249
transform -1 0 12480 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _427_
timestamp 1676627187
transform -1 0 16128 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _428_
timestamp 1676557249
transform 1 0 11520 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _429_
timestamp 1676627187
transform -1 0 15648 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _430_
timestamp 1676557249
transform -1 0 11520 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _431_
timestamp 1676627187
transform -1 0 20064 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _432_
timestamp 1676557249
transform 1 0 14880 0 1 9072
box -48 -56 432 834
use sg13g2_and3_2  _433_
timestamp 1683976310
transform -1 0 22944 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _434_
timestamp 1683988354
transform -1 0 23040 0 1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _435_
timestamp 1676627187
transform -1 0 22560 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _436_
timestamp 1676557249
transform 1 0 9600 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _437_
timestamp 1676627187
transform -1 0 22944 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _438_
timestamp 1676557249
transform 1 0 8832 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _439_
timestamp 1676627187
transform -1 0 21408 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _440_
timestamp 1676557249
transform 1 0 9216 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _441_
timestamp 1676627187
transform -1 0 23712 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _442_
timestamp 1676557249
transform 1 0 9984 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _443_
timestamp 1676627187
transform -1 0 21408 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _444_
timestamp 1676557249
transform 1 0 11904 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _445_
timestamp 1676627187
transform -1 0 19296 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _446_
timestamp 1676557249
transform 1 0 12672 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _447_
timestamp 1676627187
transform -1 0 20256 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _448_
timestamp 1676557249
transform 1 0 13440 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _449_
timestamp 1676627187
transform 1 0 17472 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _450_
timestamp 1676557249
transform 1 0 13056 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _451_
timestamp 1676627187
transform -1 0 18816 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _452_
timestamp 1676557249
transform 1 0 14496 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _453_
timestamp 1676627187
transform -1 0 18432 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _454_
timestamp 1676557249
transform 1 0 15264 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _455_
timestamp 1676627187
transform -1 0 18432 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _456_
timestamp 1676557249
transform -1 0 16032 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _457_
timestamp 1676627187
transform -1 0 19680 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _458_
timestamp 1676557249
transform 1 0 15648 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _459_
timestamp 1676627187
transform -1 0 18912 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _460_
timestamp 1676557249
transform 1 0 11520 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _461_
timestamp 1676627187
transform -1 0 19200 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _462_
timestamp 1676557249
transform 1 0 11712 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _463_
timestamp 1676627187
transform 1 0 17664 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _464_
timestamp 1676557249
transform 1 0 10752 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _465_
timestamp 1676627187
transform -1 0 19680 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _466_
timestamp 1676557249
transform 1 0 16032 0 1 9072
box -48 -56 432 834
use sg13g2_and3_1  _467_
timestamp 1676971669
transform -1 0 23616 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _468_
timestamp 1683988354
transform -1 0 24864 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _469_
timestamp 1676627187
transform -1 0 25248 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _470_
timestamp 1676557249
transform 1 0 18144 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _471_
timestamp 1676627187
transform -1 0 24864 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _472_
timestamp 1676557249
transform -1 0 18912 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _473_
timestamp 1676627187
transform -1 0 24480 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _474_
timestamp 1676557249
transform -1 0 18144 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _475_
timestamp 1676627187
transform -1 0 25248 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _476_
timestamp 1676557249
transform 1 0 18624 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _477_
timestamp 1676627187
transform -1 0 25632 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _478_
timestamp 1676557249
transform 1 0 19296 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _479_
timestamp 1676627187
transform -1 0 24864 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _480_
timestamp 1676557249
transform 1 0 18912 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _481_
timestamp 1676627187
transform 1 0 23712 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _482_
timestamp 1676557249
transform -1 0 20064 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _483_
timestamp 1676627187
transform -1 0 24480 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _484_
timestamp 1676557249
transform 1 0 18528 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _485_
timestamp 1676627187
transform -1 0 25248 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _486_
timestamp 1676557249
transform -1 0 20064 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _487_
timestamp 1676627187
transform -1 0 23904 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _488_
timestamp 1676557249
transform 1 0 20064 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _489_
timestamp 1676627187
transform 1 0 23136 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _490_
timestamp 1676557249
transform 1 0 19392 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _491_
timestamp 1676627187
transform -1 0 24096 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _492_
timestamp 1676557249
transform 1 0 19680 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _493_
timestamp 1676627187
transform -1 0 25632 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _494_
timestamp 1676557249
transform 1 0 19296 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _495_
timestamp 1676627187
transform -1 0 24288 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _496_
timestamp 1676557249
transform 1 0 19296 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _497_
timestamp 1676627187
transform -1 0 24480 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _498_
timestamp 1676557249
transform 1 0 18912 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _499_
timestamp 1676627187
transform -1 0 24672 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _500_
timestamp 1676557249
transform 1 0 18912 0 1 9072
box -48 -56 432 834
use sg13g2_nand3_1  _501_
timestamp 1683988354
transform 1 0 39360 0 1 7560
box -48 -56 528 834
use sg13g2_nor2_1  _502_
timestamp 1676627187
transform -1 0 34272 0 -1 9072
box -48 -56 432 834
use sg13g2_nand2b_1  _503_
timestamp 1676567195
transform -1 0 33408 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _504_
timestamp 1676627187
transform -1 0 28704 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _505_
timestamp 1676557249
transform -1 0 25632 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _506_
timestamp 1676627187
transform -1 0 28320 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _507_
timestamp 1676557249
transform -1 0 24864 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _508_
timestamp 1676627187
transform -1 0 27936 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _509_
timestamp 1676557249
transform 1 0 25632 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _510_
timestamp 1676627187
transform -1 0 29088 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _511_
timestamp 1676557249
transform 1 0 24960 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _512_
timestamp 1676627187
transform -1 0 28320 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _513_
timestamp 1676557249
transform 1 0 24480 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _514_
timestamp 1676627187
transform 1 0 27168 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _515_
timestamp 1676557249
transform 1 0 24864 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _516_
timestamp 1676627187
transform -1 0 28800 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _517_
timestamp 1676557249
transform 1 0 24864 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _518_
timestamp 1676627187
transform 1 0 27552 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _519_
timestamp 1676557249
transform -1 0 24480 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _520_
timestamp 1676627187
transform -1 0 27264 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _521_
timestamp 1676557249
transform 1 0 24480 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _522_
timestamp 1676627187
transform 1 0 26496 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _523_
timestamp 1676557249
transform 1 0 24864 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _524_
timestamp 1676627187
transform 1 0 26880 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _525_
timestamp 1676557249
transform 1 0 24480 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _526_
timestamp 1676627187
transform 1 0 27648 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _527_
timestamp 1676557249
transform 1 0 24480 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _528_
timestamp 1676627187
transform 1 0 26112 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _529_
timestamp 1676557249
transform -1 0 24096 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _530_
timestamp 1676627187
transform 1 0 26880 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _531_
timestamp 1676557249
transform 1 0 24096 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _532_
timestamp 1676627187
transform 1 0 27264 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _533_
timestamp 1676557249
transform 1 0 24096 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _534_
timestamp 1676627187
transform 1 0 26496 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _535_
timestamp 1676557249
transform 1 0 24096 0 1 10584
box -48 -56 432 834
use sg13g2_and3_1  _536_
timestamp 1676971669
transform 1 0 29664 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _537_
timestamp 1683988354
transform -1 0 30144 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _538_
timestamp 1676627187
transform -1 0 30624 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _539_
timestamp 1676557249
transform 1 0 28320 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _540_
timestamp 1676627187
transform -1 0 31392 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _541_
timestamp 1676557249
transform 1 0 27936 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _542_
timestamp 1676627187
transform 1 0 30240 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _543_
timestamp 1676557249
transform 1 0 28704 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _544_
timestamp 1676627187
transform 1 0 30624 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _545_
timestamp 1676557249
transform 1 0 27552 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _546_
timestamp 1676627187
transform 1 0 31008 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _547_
timestamp 1676557249
transform 1 0 28128 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _548_
timestamp 1676627187
transform -1 0 31968 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _549_
timestamp 1676557249
transform 1 0 27744 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _550_
timestamp 1676627187
transform 1 0 30624 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _551_
timestamp 1676557249
transform 1 0 28512 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _552_
timestamp 1676627187
transform 1 0 29856 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _553_
timestamp 1676557249
transform -1 0 27744 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _554_
timestamp 1676627187
transform 1 0 32160 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _555_
timestamp 1676557249
transform 1 0 31104 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _556_
timestamp 1676627187
transform 1 0 31776 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _557_
timestamp 1676557249
transform 1 0 30912 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _558_
timestamp 1676627187
transform 1 0 32160 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _559_
timestamp 1676557249
transform 1 0 30528 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _560_
timestamp 1676627187
transform 1 0 31776 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _561_
timestamp 1676557249
transform 1 0 30912 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _562_
timestamp 1676627187
transform 1 0 32544 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _563_
timestamp 1676557249
transform 1 0 31296 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _564_
timestamp 1676627187
transform 1 0 32544 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _565_
timestamp 1676557249
transform 1 0 30720 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _566_
timestamp 1676627187
transform 1 0 31392 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _567_
timestamp 1676557249
transform 1 0 30144 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _568_
timestamp 1676627187
transform 1 0 31392 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _569_
timestamp 1676557249
transform 1 0 30528 0 1 9072
box -48 -56 432 834
use sg13g2_and3_1  _570_
timestamp 1676971669
transform 1 0 36480 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _571_
timestamp 1683988354
transform 1 0 35808 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _572_
timestamp 1676627187
transform -1 0 36864 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _573_
timestamp 1676557249
transform 1 0 34368 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _574_
timestamp 1676627187
transform 1 0 36384 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _575_
timestamp 1676557249
transform 1 0 35040 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _576_
timestamp 1676627187
transform 1 0 36000 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _577_
timestamp 1676557249
transform 1 0 34656 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _578_
timestamp 1676627187
transform 1 0 35616 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _579_
timestamp 1676557249
transform 1 0 34752 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _580_
timestamp 1676627187
transform 1 0 35232 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _581_
timestamp 1676557249
transform 1 0 34272 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _582_
timestamp 1676627187
transform 1 0 34848 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _583_
timestamp 1676557249
transform 1 0 35424 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _584_
timestamp 1676627187
transform 1 0 34464 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _585_
timestamp 1676557249
transform 1 0 34752 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _586_
timestamp 1676627187
transform 1 0 34848 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _587_
timestamp 1676557249
transform 1 0 34368 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _588_
timestamp 1676627187
transform 1 0 34368 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _589_
timestamp 1676557249
transform 1 0 36576 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _590_
timestamp 1676627187
transform 1 0 33984 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _591_
timestamp 1676557249
transform 1 0 36768 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _592_
timestamp 1676627187
transform 1 0 34752 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _593_
timestamp 1676557249
transform 1 0 36384 0 1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _594_
timestamp 1676627187
transform 1 0 34464 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _595_
timestamp 1676557249
transform 1 0 36672 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _596_
timestamp 1676627187
transform 1 0 34176 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _597_
timestamp 1676557249
transform 1 0 36288 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _598_
timestamp 1676627187
transform 1 0 34080 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _599_
timestamp 1676557249
transform 1 0 35904 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _600_
timestamp 1676627187
transform 1 0 33600 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _601_
timestamp 1676557249
transform -1 0 35904 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _602_
timestamp 1676627187
transform 1 0 33792 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _603_
timestamp 1676557249
transform 1 0 36192 0 1 9072
box -48 -56 432 834
use sg13g2_and3_1  _604_
timestamp 1676971669
transform 1 0 37152 0 1 7560
box -48 -56 720 834
use sg13g2_nand3_1  _605_
timestamp 1683988354
transform -1 0 38016 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _606_
timestamp 1676627187
transform 1 0 37920 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _607_
timestamp 1676557249
transform 1 0 31104 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _608_
timestamp 1676627187
transform 1 0 38208 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _609_
timestamp 1676557249
transform 1 0 32544 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _610_
timestamp 1676627187
transform 1 0 38592 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _611_
timestamp 1676557249
transform -1 0 31104 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _612_
timestamp 1676627187
transform 1 0 38688 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _613_
timestamp 1676557249
transform 1 0 33024 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _614_
timestamp 1676627187
transform 1 0 37536 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _615_
timestamp 1676557249
transform 1 0 32256 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _616_
timestamp 1676627187
transform -1 0 39936 0 1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _617_
timestamp 1676557249
transform 1 0 31488 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _618_
timestamp 1676627187
transform 1 0 39072 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _619_
timestamp 1676557249
transform 1 0 31872 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _620_
timestamp 1676627187
transform 1 0 38304 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _621_
timestamp 1676557249
transform 1 0 32640 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _622_
timestamp 1676627187
transform 1 0 37248 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _623_
timestamp 1676557249
transform 1 0 38688 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _624_
timestamp 1676627187
transform 1 0 38592 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _625_
timestamp 1676557249
transform -1 0 37728 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _626_
timestamp 1676627187
transform 1 0 36768 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _627_
timestamp 1676557249
transform 1 0 38304 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _628_
timestamp 1676627187
transform 1 0 39072 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _629_
timestamp 1676557249
transform 1 0 38880 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _630_
timestamp 1676627187
transform 1 0 37824 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _631_
timestamp 1676557249
transform 1 0 38496 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _632_
timestamp 1676627187
transform 1 0 37632 0 -1 7560
box -48 -56 432 834
use sg13g2_nand2_1  _633_
timestamp 1676557249
transform 1 0 38112 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _634_
timestamp 1676627187
transform 1 0 38016 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _635_
timestamp 1676557249
transform 1 0 37728 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _636_
timestamp 1676627187
transform 1 0 37440 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _637_
timestamp 1676557249
transform 1 0 37920 0 1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _638_
timestamp 1676627187
transform 1 0 55104 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _639_
timestamp 1684236171
transform -1 0 55008 0 1 3024
box -48 -56 528 834
use sg13g2_nor2_1  _640_
timestamp 1676627187
transform -1 0 50592 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _641_
timestamp 1684236171
transform 1 0 49824 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _642_
timestamp 1676627187
transform -1 0 50976 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _643_
timestamp 1684236171
transform 1 0 49920 0 1 3024
box -48 -56 528 834
use sg13g2_nor2_1  _644_
timestamp 1676627187
transform -1 0 52704 0 -1 4536
box -48 -56 432 834
use sg13g2_or2_1  _645_
timestamp 1684236171
transform -1 0 52896 0 1 3024
box -48 -56 528 834
use sg13g2_nor2_1  _646_
timestamp 1676627187
transform -1 0 54624 0 -1 6048
box -48 -56 432 834
use sg13g2_or2_1  _647_
timestamp 1684236171
transform -1 0 55200 0 1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _648_
timestamp 1676627187
transform -1 0 56736 0 1 7560
box -48 -56 432 834
use sg13g2_or2_1  _649_
timestamp 1684236171
transform -1 0 57024 0 -1 9072
box -48 -56 528 834
use sg13g2_nor2_1  _650_
timestamp 1676627187
transform 1 0 54240 0 -1 9072
box -48 -56 432 834
use sg13g2_or2_1  _651_
timestamp 1684236171
transform -1 0 55104 0 -1 9072
box -48 -56 528 834
use sg13g2_nor2_1  _652_
timestamp 1676627187
transform -1 0 58560 0 1 7560
box -48 -56 432 834
use sg13g2_or2_1  _653_
timestamp 1684236171
transform -1 0 59136 0 1 7560
box -48 -56 528 834
use sg13g2_nor2_1  _654_
timestamp 1676627187
transform -1 0 57696 0 1 6048
box -48 -56 432 834
use sg13g2_or2_1  _655_
timestamp 1684236171
transform -1 0 57504 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _656_
timestamp 1676627187
transform -1 0 57408 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _657_
timestamp 1684236171
transform -1 0 58464 0 -1 6048
box -48 -56 528 834
use sg13g2_nor2_1  _658_
timestamp 1676627187
transform -1 0 58560 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _659_
timestamp 1684236171
transform -1 0 57792 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2_1  _660_
timestamp 1676627187
transform -1 0 58176 0 1 4536
box -48 -56 432 834
use sg13g2_or2_1  _661_
timestamp 1684236171
transform -1 0 57504 0 1 3024
box -48 -56 528 834
use sg13g2_nor2_1  _662_
timestamp 1676627187
transform 1 0 58944 0 1 9072
box -48 -56 432 834
use sg13g2_or2_1  _663_
timestamp 1684236171
transform -1 0 58944 0 1 9072
box -48 -56 528 834
use sg13g2_nor2_1  _664_
timestamp 1676627187
transform 1 0 58848 0 -1 10584
box -48 -56 432 834
use sg13g2_or2_1  _665_
timestamp 1684236171
transform -1 0 58848 0 -1 10584
box -48 -56 528 834
use sg13g2_nor2_1  _666_
timestamp 1676627187
transform -1 0 57888 0 -1 10584
box -48 -56 432 834
use sg13g2_or2_1  _667_
timestamp 1684236171
transform -1 0 58368 0 -1 10584
box -48 -56 528 834
use sg13g2_nor2_2  _668_
timestamp 1683979924
transform 1 0 31488 0 -1 7560
box -48 -56 624 834
use sg13g2_or2_1  _669_
timestamp 1684236171
transform -1 0 32544 0 -1 7560
box -48 -56 528 834
use sg13g2_nor2_2  _670_
timestamp 1683979924
transform -1 0 35136 0 1 3024
box -48 -56 624 834
use sg13g2_nand2_1  _671_
timestamp 1676557249
transform -1 0 10368 0 -1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _672_
timestamp 1683979924
transform -1 0 36000 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _673_
timestamp 1676557249
transform -1 0 9984 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _674_
timestamp 1683979924
transform -1 0 34848 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _675_
timestamp 1676557249
transform -1 0 10368 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_2  _676_
timestamp 1683979924
transform -1 0 35424 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _677_
timestamp 1676557249
transform -1 0 10752 0 1 7560
box -48 -56 432 834
use sg13g2_nor2_1  _678_
timestamp 1676627187
transform -1 0 20256 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _679_
timestamp 1676557249
transform 1 0 11424 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_2  _680_
timestamp 1683979924
transform -1 0 29664 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _681_
timestamp 1676557249
transform 1 0 11808 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _682_
timestamp 1676627187
transform 1 0 19488 0 -1 4536
box -48 -56 432 834
use sg13g2_nand2_1  _683_
timestamp 1676557249
transform 1 0 11040 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_2  _684_
timestamp 1683979924
transform -1 0 34272 0 -1 4536
box -48 -56 624 834
use sg13g2_nand2_1  _685_
timestamp 1676557249
transform 1 0 12192 0 -1 9072
box -48 -56 432 834
use sg13g2_nor2_1  _686_
timestamp 1676627187
transform -1 0 16320 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_2  _687_
timestamp 1685180049
transform -1 0 25632 0 -1 10584
box -48 -56 624 834
use sg13g2_nor2_1  _688_
timestamp 1676627187
transform 1 0 15552 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_2  _689_
timestamp 1685180049
transform -1 0 21888 0 -1 10584
box -48 -56 624 834
use sg13g2_nor2_1  _690_
timestamp 1676627187
transform -1 0 17568 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _691_
timestamp 1676557249
transform -1 0 18912 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _692_
timestamp 1676627187
transform -1 0 20448 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _693_
timestamp 1676557249
transform -1 0 16416 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _694_
timestamp 1676627187
transform -1 0 19968 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _695_
timestamp 1676557249
transform -1 0 13056 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _696_
timestamp 1676627187
transform -1 0 16800 0 -1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _697_
timestamp 1676557249
transform -1 0 12288 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_1  _698_
timestamp 1676627187
transform -1 0 16704 0 1 6048
box -48 -56 432 834
use sg13g2_nand2_1  _699_
timestamp 1676557249
transform -1 0 12672 0 -1 10584
box -48 -56 432 834
use sg13g2_nor2_2  _700_
timestamp 1683979924
transform -1 0 31584 0 1 4536
box -48 -56 624 834
use sg13g2_nand2_2  _701_
timestamp 1685180049
transform 1 0 31872 0 -1 10584
box -48 -56 624 834
use sg13g2_buf_8  fanout1
timestamp 1676451365
transform -1 0 22944 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout2
timestamp 1676451365
transform -1 0 31488 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_2  fanout3
timestamp 1676381867
transform 1 0 11904 0 1 9072
box -48 -56 528 834
use sg13g2_buf_8  fanout4
timestamp 1676451365
transform -1 0 32640 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout5
timestamp 1676381867
transform 1 0 33408 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout6
timestamp 1676381867
transform -1 0 38688 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout7
timestamp 1676381867
transform -1 0 36480 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout8
timestamp 1676381867
transform 1 0 35232 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout9
timestamp 1676381867
transform 1 0 36864 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout10
timestamp 1676381867
transform -1 0 37536 0 1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout11
timestamp 1676381867
transform -1 0 30528 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout12
timestamp 1676381867
transform -1 0 31008 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout13
timestamp 1676381867
transform 1 0 29184 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout14
timestamp 1676381867
transform -1 0 30432 0 1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout15
timestamp 1676381867
transform 1 0 28800 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout16
timestamp 1676381867
transform 1 0 28320 0 1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout17
timestamp 1676381867
transform 1 0 25248 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout18
timestamp 1676381867
transform 1 0 25056 0 1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout19
timestamp 1676381867
transform -1 0 25152 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout20
timestamp 1676381867
transform 1 0 23904 0 1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout21
timestamp 1676381867
transform 1 0 20256 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout22
timestamp 1676381867
transform 1 0 20448 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_2  fanout23
timestamp 1676381867
transform -1 0 19296 0 -1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout24
timestamp 1676381867
transform 1 0 17856 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout25
timestamp 1676381867
transform 1 0 14016 0 1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout26
timestamp 1676451365
transform -1 0 16032 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout27
timestamp 1676381867
transform -1 0 18144 0 1 3024
box -48 -56 528 834
use sg13g2_buf_2  fanout28
timestamp 1676381867
transform 1 0 16800 0 -1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout29
timestamp 1676381867
transform 1 0 13248 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout30
timestamp 1676451365
transform -1 0 17376 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout31
timestamp 1676451365
transform 1 0 86496 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout32
timestamp 1676451365
transform 1 0 86208 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout33
timestamp 1676451365
transform 1 0 84000 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout34
timestamp 1676451365
transform 1 0 84288 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout35
timestamp 1676451365
transform -1 0 89760 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout36
timestamp 1676451365
transform 1 0 87264 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout37
timestamp 1676451365
transform -1 0 78720 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout38
timestamp 1676451365
transform 1 0 81120 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_2  fanout39
timestamp 1676381867
transform -1 0 81216 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout40
timestamp 1676381867
transform -1 0 87936 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout41
timestamp 1676381867
transform 1 0 76992 0 -1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout42
timestamp 1676381867
transform -1 0 78240 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout43
timestamp 1676381867
transform 1 0 78240 0 1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout44
timestamp 1676451365
transform 1 0 79104 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout45
timestamp 1676381867
transform 1 0 71136 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout46
timestamp 1676381867
transform -1 0 73632 0 1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout47
timestamp 1676381867
transform -1 0 75648 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout48
timestamp 1676381867
transform -1 0 76320 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_8  fanout49
timestamp 1676451365
transform -1 0 40320 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout50
timestamp 1676451365
transform 1 0 63840 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout51
timestamp 1676451365
transform -1 0 53280 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_2  fanout52
timestamp 1676381867
transform -1 0 74208 0 -1 10584
box -48 -56 528 834
use sg13g2_buf_8  fanout53
timestamp 1676451365
transform -1 0 43104 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout54
timestamp 1676451365
transform 1 0 65088 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout55
timestamp 1676451365
transform -1 0 53664 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout56
timestamp 1676381867
transform -1 0 73728 0 -1 10584
box -48 -56 528 834
use sg13g2_buf_8  fanout57
timestamp 1676451365
transform -1 0 49824 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout58
timestamp 1676381867
transform -1 0 69024 0 1 6048
box -48 -56 528 834
use sg13g2_buf_8  fanout59
timestamp 1676451365
transform -1 0 50496 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_2  fanout60
timestamp 1676381867
transform -1 0 69984 0 -1 10584
box -48 -56 528 834
use sg13g2_buf_8  fanout61
timestamp 1676451365
transform -1 0 41856 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout62
timestamp 1676381867
transform -1 0 65376 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout63
timestamp 1676451365
transform -1 0 41760 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout64
timestamp 1676381867
transform -1 0 70944 0 1 9072
box -48 -56 528 834
use sg13g2_buf_8  fanout65
timestamp 1676451365
transform -1 0 44640 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout66
timestamp 1676381867
transform -1 0 66816 0 1 6048
box -48 -56 528 834
use sg13g2_buf_8  fanout67
timestamp 1676451365
transform -1 0 43008 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  fanout68
timestamp 1676451365
transform 1 0 68256 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  fanout69
timestamp 1676451365
transform -1 0 42816 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout70
timestamp 1676451365
transform 1 0 64416 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout71
timestamp 1676451365
transform -1 0 41760 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  fanout72
timestamp 1676451365
transform 1 0 64992 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_8  fanout73
timestamp 1676451365
transform -1 0 40512 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout74
timestamp 1676381867
transform -1 0 67200 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout75
timestamp 1676451365
transform -1 0 40512 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_8  fanout76
timestamp 1676451365
transform 1 0 61920 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_8  fanout77
timestamp 1676451365
transform -1 0 36384 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout78
timestamp 1676451365
transform 1 0 62880 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout79
timestamp 1676451365
transform -1 0 41568 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout80
timestamp 1676451365
transform 1 0 62496 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout81
timestamp 1676451365
transform -1 0 43584 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_8  fanout82
timestamp 1676451365
transform 1 0 63840 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout83
timestamp 1676451365
transform -1 0 48672 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout84
timestamp 1676451365
transform 1 0 59040 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout85
timestamp 1676451365
transform -1 0 41088 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_2  fanout86
timestamp 1676381867
transform -1 0 64896 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout87
timestamp 1676451365
transform -1 0 42336 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_2  fanout88
timestamp 1676381867
transform -1 0 67584 0 1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout89
timestamp 1676451365
transform -1 0 43488 0 1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout90
timestamp 1676381867
transform -1 0 67392 0 -1 9072
box -48 -56 528 834
use sg13g2_buf_8  fanout91
timestamp 1676451365
transform -1 0 43584 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_2  fanout92
timestamp 1676381867
transform -1 0 68064 0 1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout93
timestamp 1676451365
transform -1 0 43680 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_2  fanout94
timestamp 1676381867
transform -1 0 69120 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout95
timestamp 1676381867
transform 1 0 71520 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout96
timestamp 1676381867
transform -1 0 72480 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout97
timestamp 1676381867
transform 1 0 53760 0 1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout98
timestamp 1676381867
transform 1 0 59328 0 1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout99
timestamp 1676381867
transform 1 0 59040 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform 1 0 59904 0 1 7560
box -48 -56 432 834
use sg13g2_buf_2  fanout101
timestamp 1676381867
transform -1 0 55008 0 -1 4536
box -48 -56 528 834
use sg13g2_buf_8  fanout102
timestamp 1676451365
transform -1 0 60384 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_2  fanout103
timestamp 1676381867
transform 1 0 58080 0 1 6048
box -48 -56 528 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform -1 0 59040 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform -1 0 61152 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_8  fanout106
timestamp 1676451365
transform 1 0 52128 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform 1 0 52992 0 1 6048
box -48 -56 432 834
use sg13g2_buf_2  fanout108
timestamp 1676381867
transform 1 0 46944 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform 1 0 54336 0 1 7560
box -48 -56 432 834
use sg13g2_buf_8  fanout110
timestamp 1676451365
transform -1 0 47328 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_1  fanout111
timestamp 1676381911
transform 1 0 48192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_8  fanout112
timestamp 1676451365
transform -1 0 48576 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_1  fanout113
timestamp 1676381911
transform 1 0 48672 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_8  fanout114
timestamp 1676451365
transform 1 0 50304 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_1  fanout115
timestamp 1676381911
transform 1 0 50496 0 1 7560
box -48 -56 432 834
use sg13g2_buf_2  fanout116
timestamp 1676381867
transform 1 0 45984 0 1 6048
box -48 -56 528 834
use sg13g2_buf_1  fanout117
timestamp 1676381911
transform -1 0 50208 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_8  fanout118
timestamp 1676451365
transform -1 0 49536 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout119
timestamp 1676381867
transform -1 0 52032 0 1 7560
box -48 -56 528 834
use sg13g2_buf_8  fanout120
timestamp 1676451365
transform -1 0 30240 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_1  fanout121
timestamp 1676381911
transform 1 0 36384 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_8  fanout122
timestamp 1676451365
transform -1 0 60192 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout123
timestamp 1676451365
transform -1 0 45888 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_2  fanout124
timestamp 1676381867
transform 1 0 45600 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_1  fanout125
timestamp 1676381911
transform -1 0 47328 0 1 6048
box -48 -56 432 834
use sg13g2_buf_2  fanout126
timestamp 1676381867
transform -1 0 48960 0 -1 7560
box -48 -56 528 834
use sg13g2_buf_2  fanout127
timestamp 1676381867
transform -1 0 51072 0 1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout128
timestamp 1676381867
transform -1 0 55968 0 1 6048
box -48 -56 528 834
use sg13g2_buf_1  fanout129
timestamp 1676381911
transform 1 0 53088 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_2  fanout130
timestamp 1676381867
transform -1 0 39456 0 1 4536
box -48 -56 528 834
use sg13g2_buf_2  fanout131
timestamp 1676381867
transform -1 0 38976 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_8  fanout132
timestamp 1676451365
transform -1 0 46848 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout133
timestamp 1676451365
transform 1 0 64608 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout134
timestamp 1676451365
transform -1 0 44832 0 -1 9072
box -48 -56 1296 834
use sg13g2_buf_8  fanout135
timestamp 1676451365
transform 1 0 65088 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  fanout136
timestamp 1676451365
transform -1 0 47424 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout137
timestamp 1676451365
transform 1 0 57792 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout138
timestamp 1676451365
transform -1 0 47712 0 1 3024
box -48 -56 1296 834
use sg13g2_buf_2  fanout139
timestamp 1676381867
transform -1 0 62976 0 1 3024
box -48 -56 528 834
use sg13g2_buf_8  fanout140
timestamp 1676451365
transform -1 0 46176 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout141
timestamp 1676451365
transform 1 0 63168 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout142
timestamp 1676451365
transform -1 0 43296 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_2  fanout143
timestamp 1676381867
transform -1 0 63648 0 1 4536
box -48 -56 528 834
use sg13g2_buf_8  fanout144
timestamp 1676451365
transform -1 0 44928 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_2  fanout145
timestamp 1676381867
transform -1 0 62496 0 1 4536
box -48 -56 528 834
use sg13g2_buf_8  fanout146
timestamp 1676451365
transform -1 0 45792 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout147
timestamp 1676451365
transform 1 0 52608 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout148
timestamp 1676451365
transform -1 0 44544 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  fanout149
timestamp 1676451365
transform 1 0 53856 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_2  fanout150
timestamp 1676381867
transform 1 0 67104 0 -1 6048
box -48 -56 528 834
use sg13g2_buf_2  fanout151
timestamp 1676381867
transform -1 0 67968 0 1 6048
box -48 -56 528 834
use sg13g2_buf_8  fanout152
timestamp 1676451365
transform -1 0 37536 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  fanout153
timestamp 1676451365
transform 1 0 80928 0 1 3024
box -48 -56 1296 834
use sg13g2_buf_8  fanout154
timestamp 1676451365
transform 1 0 74496 0 1 4536
box -48 -56 1296 834
use sg13g2_fill_2  FILLER_0_177
timestamp 1677580104
transform 1 0 18144 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_179
timestamp 1677579658
transform 1 0 18336 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_354
timestamp 1677579658
transform 1 0 35136 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_485
timestamp 1677580104
transform 1 0 47712 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_533
timestamp 1677579658
transform 1 0 52320 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_555
timestamp 1677579658
transform 1 0 54432 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_581
timestamp 1677579658
transform 1 0 56928 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_603
timestamp 1677580104
transform 1 0 59040 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_605
timestamp 1677579658
transform 1 0 59232 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_638
timestamp 1677579658
transform 1 0 62400 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_828
timestamp 1677580104
transform 1 0 80640 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_830
timestamp 1677579658
transform 1 0 80832 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_1016
timestamp 1677579658
transform 1 0 98688 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_2
timestamp 1677579658
transform 1 0 1344 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_189
timestamp 1677580104
transform 1 0 19296 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_297
timestamp 1677580104
transform 1 0 29664 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_495
timestamp 1677580104
transform 1 0 48672 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_497
timestamp 1677579658
transform 1 0 48864 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_512
timestamp 1677580104
transform 1 0 50304 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_514
timestamp 1677579658
transform 1 0 50496 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_537
timestamp 1677579658
transform 1 0 52704 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_555
timestamp 1677579658
transform 1 0 54432 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_573
timestamp 1677580104
transform 1 0 56160 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_643
timestamp 1677580104
transform 1 0 62880 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_645
timestamp 1677579658
transform 1 0 63072 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_681
timestamp 1677580104
transform 1 0 66528 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_789
timestamp 1677579658
transform 1 0 76896 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_832
timestamp 1677579658
transform 1 0 81024 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_862
timestamp 1677579658
transform 1 0 83904 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_1016
timestamp 1677579658
transform 1 0 98688 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_2
timestamp 1677579658
transform 1 0 1344 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_19
timestamp 1679581782
transform 1 0 2976 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_26
timestamp 1679581782
transform 1 0 3648 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_33
timestamp 1679581782
transform 1 0 4320 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_40
timestamp 1679581782
transform 1 0 4992 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_47
timestamp 1679581782
transform 1 0 5664 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_54
timestamp 1679581782
transform 1 0 6336 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_61
timestamp 1679581782
transform 1 0 7008 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_68
timestamp 1679581782
transform 1 0 7680 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_75
timestamp 1679581782
transform 1 0 8352 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_82
timestamp 1679581782
transform 1 0 9024 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_89
timestamp 1679581782
transform 1 0 9696 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_96
timestamp 1679581782
transform 1 0 10368 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_103
timestamp 1679581782
transform 1 0 11040 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_110
timestamp 1679581782
transform 1 0 11712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_117
timestamp 1679581782
transform 1 0 12384 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_124
timestamp 1679577901
transform 1 0 13056 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_156
timestamp 1677580104
transform 1 0 16128 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_179
timestamp 1677580104
transform 1 0 18336 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_193
timestamp 1677580104
transform 1 0 19680 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_228
timestamp 1677580104
transform 1 0 23040 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_230
timestamp 1677579658
transform 1 0 23232 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_321
timestamp 1677580104
transform 1 0 31968 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_372
timestamp 1677580104
transform 1 0 36864 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_399
timestamp 1677579658
transform 1 0 39456 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_404
timestamp 1677580104
transform 1 0 39936 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_470
timestamp 1677580104
transform 1 0 46272 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_519
timestamp 1679581782
transform 1 0 50976 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_526
timestamp 1679577901
transform 1 0 51648 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_530
timestamp 1677579658
transform 1 0 52032 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_535
timestamp 1677579658
transform 1 0 52512 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_606
timestamp 1677580104
transform 1 0 59328 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_622
timestamp 1677580104
transform 1 0 60864 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_624
timestamp 1677579658
transform 1 0 61056 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_643
timestamp 1677580104
transform 1 0 62880 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_645
timestamp 1677579658
transform 1 0 63072 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_659
timestamp 1677580104
transform 1 0 64416 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_686
timestamp 1677579658
transform 1 0 67008 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_711
timestamp 1677579658
transform 1 0 69408 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_736
timestamp 1677579658
transform 1 0 71808 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_757
timestamp 1677580104
transform 1 0 73824 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_759
timestamp 1677579658
transform 1 0 74016 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_797
timestamp 1677579658
transform 1 0 77664 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_811
timestamp 1677580104
transform 1 0 79008 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_853
timestamp 1677580104
transform 1 0 83040 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_863
timestamp 1677580104
transform 1 0 84000 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_865
timestamp 1677579658
transform 1 0 84192 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_911
timestamp 1679581782
transform 1 0 88608 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_918
timestamp 1679581782
transform 1 0 89280 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_925
timestamp 1679581782
transform 1 0 89952 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_932
timestamp 1679581782
transform 1 0 90624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_939
timestamp 1679581782
transform 1 0 91296 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_946
timestamp 1679581782
transform 1 0 91968 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_953
timestamp 1679581782
transform 1 0 92640 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_960
timestamp 1679581782
transform 1 0 93312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_967
timestamp 1679581782
transform 1 0 93984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_974
timestamp 1679581782
transform 1 0 94656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_981
timestamp 1679581782
transform 1 0 95328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_988
timestamp 1679581782
transform 1 0 96000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_995
timestamp 1679577901
transform 1 0 96672 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_1015
timestamp 1677580104
transform 1 0 98592 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_0
timestamp 1677580104
transform 1 0 1152 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_2
timestamp 1677579658
transform 1 0 1344 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 2208 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2880 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 3552 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 4224 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4896 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 5568 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 6240 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6912 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7584 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 8256 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9600 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 10272 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10944 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11616 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 12288 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12960 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13632 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 14304 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_144
timestamp 1677580104
transform 1 0 14976 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_146
timestamp 1677579658
transform 1 0 15168 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_171
timestamp 1677579658
transform 1 0 17568 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_180
timestamp 1677579658
transform 1 0 18432 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_205
timestamp 1677579658
transform 1 0 20832 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_232
timestamp 1677580104
transform 1 0 23424 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_234
timestamp 1677579658
transform 1 0 23616 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_243
timestamp 1677580104
transform 1 0 24480 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_250
timestamp 1679581782
transform 1 0 25152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_257
timestamp 1679581782
transform 1 0 25824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_272
timestamp 1679581782
transform 1 0 27264 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_279
timestamp 1677579658
transform 1 0 27936 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_331
timestamp 1679581782
transform 1 0 32928 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_338
timestamp 1677579658
transform 1 0 33600 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_360
timestamp 1677580104
transform 1 0 35712 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_362
timestamp 1677579658
transform 1 0 35904 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_386
timestamp 1677580104
transform 1 0 38208 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_388
timestamp 1677579658
transform 1 0 38400 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_394
timestamp 1677579658
transform 1 0 38976 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_407
timestamp 1679581782
transform 1 0 40224 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_414
timestamp 1677579658
transform 1 0 40896 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_419
timestamp 1677580104
transform 1 0 41376 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_456
timestamp 1677579658
transform 1 0 44928 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_462
timestamp 1677579658
transform 1 0 45504 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_476
timestamp 1677580104
transform 1 0 46848 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_511
timestamp 1679581782
transform 1 0 50208 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_518
timestamp 1679581782
transform 1 0 50880 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_525
timestamp 1679577901
transform 1 0 51552 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_529
timestamp 1677580104
transform 1 0 51936 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_536
timestamp 1679577901
transform 1 0 52608 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_540
timestamp 1677579658
transform 1 0 52992 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_545
timestamp 1677580104
transform 1 0 53472 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_551
timestamp 1677580104
transform 1 0 54048 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_565
timestamp 1677580104
transform 1 0 55392 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_571
timestamp 1677580104
transform 1 0 55968 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_573
timestamp 1677579658
transform 1 0 56160 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_621
timestamp 1677580104
transform 1 0 60768 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_656
timestamp 1677580104
transform 1 0 64128 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_658
timestamp 1677579658
transform 1 0 64320 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_672
timestamp 1679581782
transform 1 0 65664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_679
timestamp 1679577901
transform 1 0 66336 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_696
timestamp 1677580104
transform 1 0 67968 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_698
timestamp 1677579658
transform 1 0 68160 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_711
timestamp 1677579658
transform 1 0 69408 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_728
timestamp 1677579658
transform 1 0 71040 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_734
timestamp 1677580104
transform 1 0 71616 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_736
timestamp 1677579658
transform 1 0 71808 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_749
timestamp 1677580104
transform 1 0 73056 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_751
timestamp 1677579658
transform 1 0 73248 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_796
timestamp 1677579658
transform 1 0 77568 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_803
timestamp 1677580104
transform 1 0 78240 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_829
timestamp 1677579658
transform 1 0 80736 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_842
timestamp 1677579658
transform 1 0 81984 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_863
timestamp 1677580104
transform 1 0 84000 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_891
timestamp 1679581782
transform 1 0 86688 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_898
timestamp 1679581782
transform 1 0 87360 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_905
timestamp 1679581782
transform 1 0 88032 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_912
timestamp 1679581782
transform 1 0 88704 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_919
timestamp 1679581782
transform 1 0 89376 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_926
timestamp 1679581782
transform 1 0 90048 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_933
timestamp 1679581782
transform 1 0 90720 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_940
timestamp 1679581782
transform 1 0 91392 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_947
timestamp 1679581782
transform 1 0 92064 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_954
timestamp 1679581782
transform 1 0 92736 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_961
timestamp 1679581782
transform 1 0 93408 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_968
timestamp 1679581782
transform 1 0 94080 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_975
timestamp 1679581782
transform 1 0 94752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_982
timestamp 1679581782
transform 1 0 95424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_989
timestamp 1679581782
transform 1 0 96096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_996
timestamp 1679581782
transform 1 0 96768 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1015
timestamp 1677580104
transform 1 0 98592 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 1536 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 2208 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2880 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 3552 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 4224 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4896 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 5568 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 6240 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6912 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7584 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 8256 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8928 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9600 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_95
timestamp 1677579658
transform 1 0 10272 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_100
timestamp 1679581782
transform 1 0 10752 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_107
timestamp 1679581782
transform 1 0 11424 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_114
timestamp 1679581782
transform 1 0 12096 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_121
timestamp 1679581782
transform 1 0 12768 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_128
timestamp 1679581782
transform 1 0 13440 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_135
timestamp 1679581782
transform 1 0 14112 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_142
timestamp 1679581782
transform 1 0 14784 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_149
timestamp 1677579658
transform 1 0 15456 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_162
timestamp 1679581782
transform 1 0 16704 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_169
timestamp 1677580104
transform 1 0 17376 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_171
timestamp 1677579658
transform 1 0 17568 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_196
timestamp 1679577901
transform 1 0 19968 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_200
timestamp 1677579658
transform 1 0 20352 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_209
timestamp 1679581782
transform 1 0 21216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_216
timestamp 1679581782
transform 1 0 21888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_223
timestamp 1679577901
transform 1 0 22560 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_227
timestamp 1677580104
transform 1 0 22944 0 1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_255
timestamp 1679577901
transform 1 0 25632 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_259
timestamp 1677579658
transform 1 0 26016 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_280
timestamp 1677580104
transform 1 0 28032 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_282
timestamp 1677579658
transform 1 0 28224 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_288
timestamp 1679581782
transform 1 0 28800 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_295
timestamp 1677580104
transform 1 0 29472 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1679581782
transform 1 0 30144 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_309
timestamp 1679577901
transform 1 0 30816 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_313
timestamp 1677580104
transform 1 0 31200 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_336
timestamp 1677580104
transform 1 0 33408 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_354
timestamp 1677580104
transform 1 0 35136 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_356
timestamp 1677579658
transform 1 0 35328 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_388
timestamp 1677580104
transform 1 0 38400 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_394
timestamp 1677580104
transform 1 0 38976 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_396
timestamp 1677579658
transform 1 0 39168 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_410
timestamp 1677579658
transform 1 0 40512 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_437
timestamp 1677580104
transform 1 0 43104 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_439
timestamp 1677579658
transform 1 0 43296 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_466
timestamp 1677579658
transform 1 0 45888 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_472
timestamp 1677579658
transform 1 0 46464 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_485
timestamp 1677579658
transform 1 0 47712 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_504
timestamp 1679577901
transform 1 0 49536 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_508
timestamp 1677580104
transform 1 0 49920 0 1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_544
timestamp 1679577901
transform 1 0 53376 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_563
timestamp 1677580104
transform 1 0 55200 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_565
timestamp 1677579658
transform 1 0 55392 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_575
timestamp 1677579658
transform 1 0 56352 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_628
timestamp 1677580104
transform 1 0 61440 0 1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_647
timestamp 1679577901
transform 1 0 63264 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_651
timestamp 1677580104
transform 1 0 63648 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_684
timestamp 1677580104
transform 1 0 66816 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_686
timestamp 1677579658
transform 1 0 67008 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_700
timestamp 1677580104
transform 1 0 68352 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_715
timestamp 1679581782
transform 1 0 69792 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_722
timestamp 1679577901
transform 1 0 70464 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_726
timestamp 1677579658
transform 1 0 70848 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_740
timestamp 1679577901
transform 1 0 72192 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_748
timestamp 1677580104
transform 1 0 72960 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_755
timestamp 1677580104
transform 1 0 73632 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_757
timestamp 1677579658
transform 1 0 73824 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_778
timestamp 1679581782
transform 1 0 75840 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_785
timestamp 1677580104
transform 1 0 76512 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_799
timestamp 1679581782
transform 1 0 77856 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_806
timestamp 1677579658
transform 1 0 78528 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_827
timestamp 1679581782
transform 1 0 80544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_834
timestamp 1679577901
transform 1 0 81216 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_838
timestamp 1677579658
transform 1 0 81600 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_847
timestamp 1677580104
transform 1 0 82464 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_865
timestamp 1677580104
transform 1 0 84192 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_867
timestamp 1677579658
transform 1 0 84384 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_873
timestamp 1679581782
transform 1 0 84960 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_880
timestamp 1679581782
transform 1 0 85632 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_887
timestamp 1677580104
transform 1 0 86304 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_889
timestamp 1677579658
transform 1 0 86496 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_894
timestamp 1677580104
transform 1 0 86976 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_896
timestamp 1677579658
transform 1 0 87168 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_910
timestamp 1679581782
transform 1 0 88512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_917
timestamp 1679581782
transform 1 0 89184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_924
timestamp 1679581782
transform 1 0 89856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_931
timestamp 1679581782
transform 1 0 90528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_938
timestamp 1679581782
transform 1 0 91200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_945
timestamp 1679581782
transform 1 0 91872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_952
timestamp 1679581782
transform 1 0 92544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_959
timestamp 1679581782
transform 1 0 93216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_966
timestamp 1679581782
transform 1 0 93888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_973
timestamp 1679581782
transform 1 0 94560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_980
timestamp 1679581782
transform 1 0 95232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_987
timestamp 1679581782
transform 1 0 95904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_994
timestamp 1679581782
transform 1 0 96576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1001
timestamp 1679581782
transform 1 0 97248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_1008
timestamp 1679577901
transform 1 0 97920 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_1012
timestamp 1677579658
transform 1 0 98304 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 8544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_84
timestamp 1679577901
transform 1 0 9216 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_96
timestamp 1677580104
transform 1 0 10368 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_106
timestamp 1679577901
transform 1 0 11328 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_110
timestamp 1677579658
transform 1 0 11712 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_115
timestamp 1677580104
transform 1 0 12192 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_117
timestamp 1677579658
transform 1 0 12384 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_122
timestamp 1679577901
transform 1 0 12864 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_131
timestamp 1679581782
transform 1 0 13728 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_138
timestamp 1679581782
transform 1 0 14400 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_145
timestamp 1679581782
transform 1 0 15072 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_152
timestamp 1679581782
transform 1 0 15744 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_159
timestamp 1679581782
transform 1 0 16416 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_166
timestamp 1679581782
transform 1 0 17088 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_173
timestamp 1679581782
transform 1 0 17760 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_180
timestamp 1677580104
transform 1 0 18432 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 19008 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19680 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 20352 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 21024 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21696 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_221
timestamp 1677580104
transform 1 0 22368 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_223
timestamp 1677579658
transform 1 0 22560 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_231
timestamp 1679577901
transform 1 0 23328 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_235
timestamp 1677580104
transform 1 0 23712 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_245
timestamp 1677580104
transform 1 0 24672 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_247
timestamp 1677579658
transform 1 0 24864 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679581782
transform 1 0 25344 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_259
timestamp 1679581782
transform 1 0 26016 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_266
timestamp 1677580104
transform 1 0 26688 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_272
timestamp 1679581782
transform 1 0 27264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_279
timestamp 1679581782
transform 1 0 27936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_286
timestamp 1679577901
transform 1 0 28608 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_331
timestamp 1679581782
transform 1 0 32928 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_338
timestamp 1677580104
transform 1 0 33600 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_348
timestamp 1679581782
transform 1 0 34560 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_355
timestamp 1679581782
transform 1 0 35232 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_362
timestamp 1679577901
transform 1 0 35904 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_366
timestamp 1677579658
transform 1 0 36288 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_371
timestamp 1679577901
transform 1 0 36768 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_375
timestamp 1677579658
transform 1 0 37152 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_384
timestamp 1679581782
transform 1 0 38016 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_391
timestamp 1679577901
transform 1 0 38688 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_421
timestamp 1679581782
transform 1 0 41568 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_428
timestamp 1677580104
transform 1 0 42240 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_443
timestamp 1679577901
transform 1 0 43680 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_447
timestamp 1677580104
transform 1 0 44064 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_456
timestamp 1679581782
transform 1 0 44928 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_468
timestamp 1677580104
transform 1 0 46080 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_482
timestamp 1679581782
transform 1 0 47424 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_489
timestamp 1679577901
transform 1 0 48096 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_507
timestamp 1677579658
transform 1 0 49824 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_520
timestamp 1677579658
transform 1 0 51072 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_544
timestamp 1679581782
transform 1 0 53376 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_551
timestamp 1677580104
transform 1 0 54048 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 55296 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_579
timestamp 1677580104
transform 1 0 56736 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 57312 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_592
timestamp 1677580104
transform 1 0 57984 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_599
timestamp 1679577901
transform 1 0 58656 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_608
timestamp 1677580104
transform 1 0 59520 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_625
timestamp 1679577901
transform 1 0 61152 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_629
timestamp 1677580104
transform 1 0 61536 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_636
timestamp 1679581782
transform 1 0 62208 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_656
timestamp 1677580104
transform 1 0 64128 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_658
timestamp 1677579658
transform 1 0 64320 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 65376 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 66048 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_688
timestamp 1679581782
transform 1 0 67200 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_695
timestamp 1677579658
transform 1 0 67872 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_700
timestamp 1677579658
transform 1 0 68352 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_705
timestamp 1677579658
transform 1 0 68832 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_710
timestamp 1679581782
transform 1 0 69312 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_717
timestamp 1679577901
transform 1 0 69984 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_721
timestamp 1677579658
transform 1 0 70368 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_726
timestamp 1679581782
transform 1 0 70848 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_733
timestamp 1679581782
transform 1 0 71520 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_740
timestamp 1679581782
transform 1 0 72192 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_747
timestamp 1679581782
transform 1 0 72864 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_754
timestamp 1679581782
transform 1 0 73536 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_765
timestamp 1677580104
transform 1 0 74592 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_775
timestamp 1679581782
transform 1 0 75552 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_782
timestamp 1679581782
transform 1 0 76224 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_789
timestamp 1677579658
transform 1 0 76896 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_797
timestamp 1677580104
transform 1 0 77664 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_799
timestamp 1677579658
transform 1 0 77856 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_814
timestamp 1679581782
transform 1 0 79296 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_821
timestamp 1679581782
transform 1 0 79968 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_828
timestamp 1677579658
transform 1 0 80640 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_834
timestamp 1679581782
transform 1 0 81216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_841
timestamp 1679581782
transform 1 0 81888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_868
timestamp 1679581782
transform 1 0 84480 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_875
timestamp 1679577901
transform 1 0 85152 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_883
timestamp 1677580104
transform 1 0 85920 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_885
timestamp 1677579658
transform 1 0 86112 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_908
timestamp 1677580104
transform 1 0 88320 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_923
timestamp 1679581782
transform 1 0 89760 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_930
timestamp 1679581782
transform 1 0 90432 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_937
timestamp 1679581782
transform 1 0 91104 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_944
timestamp 1679581782
transform 1 0 91776 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_951
timestamp 1679581782
transform 1 0 92448 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_958
timestamp 1679581782
transform 1 0 93120 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_965
timestamp 1679581782
transform 1 0 93792 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_972
timestamp 1679581782
transform 1 0 94464 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_979
timestamp 1679581782
transform 1 0 95136 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_986
timestamp 1679581782
transform 1 0 95808 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_993
timestamp 1679581782
transform 1 0 96480 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1000
timestamp 1679581782
transform 1 0 97152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1007
timestamp 1679581782
transform 1 0 97824 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_1014
timestamp 1677580104
transform 1 0 98496 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_1016
timestamp 1677579658
transform 1 0 98688 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_77
timestamp 1677580104
transform 1 0 8544 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_79
timestamp 1677579658
transform 1 0 8736 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_100
timestamp 1679581782
transform 1 0 10752 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_107
timestamp 1677579658
transform 1 0 11424 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_132
timestamp 1677580104
transform 1 0 13824 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_139
timestamp 1679581782
transform 1 0 14496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_146
timestamp 1679581782
transform 1 0 15168 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_153
timestamp 1677580104
transform 1 0 15840 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_155
timestamp 1677579658
transform 1 0 16032 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_169
timestamp 1679577901
transform 1 0 17376 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_197
timestamp 1677580104
transform 1 0 20064 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_204
timestamp 1679581782
transform 1 0 20736 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_211
timestamp 1679581782
transform 1 0 21408 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_218
timestamp 1677580104
transform 1 0 22080 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_234
timestamp 1679581782
transform 1 0 23616 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_241
timestamp 1677580104
transform 1 0 24288 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 26016 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679581782
transform 1 0 26688 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_273
timestamp 1677580104
transform 1 0 27360 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_291
timestamp 1679577901
transform 1 0 29088 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_295
timestamp 1677580104
transform 1 0 29472 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_304
timestamp 1679577901
transform 1 0 30336 0 1 7560
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_341
timestamp 1679577901
transform 1 0 33888 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_345
timestamp 1677579658
transform 1 0 34272 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_367
timestamp 1677579658
transform 1 0 36384 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 38496 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_396
timestamp 1677580104
transform 1 0 39168 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_442
timestamp 1679577901
transform 1 0 43584 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_460
timestamp 1677580104
transform 1 0 45312 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_483
timestamp 1679577901
transform 1 0 47520 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_487
timestamp 1677580104
transform 1 0 47904 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_496
timestamp 1677580104
transform 1 0 48768 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_498
timestamp 1677579658
transform 1 0 48960 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_513
timestamp 1677579658
transform 1 0 50400 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_518
timestamp 1677580104
transform 1 0 50880 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_520
timestamp 1677579658
transform 1 0 51072 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_530
timestamp 1679581782
transform 1 0 52032 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_537
timestamp 1679581782
transform 1 0 52704 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_544
timestamp 1679581782
transform 1 0 53376 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_551
timestamp 1677580104
transform 1 0 54048 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_553
timestamp 1677579658
transform 1 0 54240 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_562
timestamp 1679581782
transform 1 0 55104 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_569
timestamp 1677580104
transform 1 0 55776 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_583
timestamp 1679577901
transform 1 0 57120 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_587
timestamp 1677579658
transform 1 0 57504 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_592
timestamp 1677580104
transform 1 0 57984 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_598
timestamp 1677579658
transform 1 0 58560 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_604
timestamp 1677580104
transform 1 0 59136 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_611
timestamp 1677579658
transform 1 0 59808 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_616
timestamp 1679581782
transform 1 0 60288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_623
timestamp 1679581782
transform 1 0 60960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_630
timestamp 1679581782
transform 1 0 61632 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_637
timestamp 1677580104
transform 1 0 62304 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_652
timestamp 1677579658
transform 1 0 63744 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_679
timestamp 1679581782
transform 1 0 66336 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_686
timestamp 1677579658
transform 1 0 67008 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_697
timestamp 1679577901
transform 1 0 68064 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_701
timestamp 1677580104
transform 1 0 68448 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_708
timestamp 1679577901
transform 1 0 69120 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_712
timestamp 1677580104
transform 1 0 69504 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_730
timestamp 1677580104
transform 1 0 71232 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_732
timestamp 1677579658
transform 1 0 71424 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_748
timestamp 1679581782
transform 1 0 72960 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_755
timestamp 1677580104
transform 1 0 73632 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_757
timestamp 1677579658
transform 1 0 73824 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_780
timestamp 1679581782
transform 1 0 76032 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_787
timestamp 1679581782
transform 1 0 76704 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_794
timestamp 1677579658
transform 1 0 77376 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_812
timestamp 1679581782
transform 1 0 79104 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_819
timestamp 1679581782
transform 1 0 79776 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_826
timestamp 1677580104
transform 1 0 80448 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_844
timestamp 1677580104
transform 1 0 82176 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_878
timestamp 1679581782
transform 1 0 85440 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_885
timestamp 1679577901
transform 1 0 86112 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_914
timestamp 1677579658
transform 1 0 88896 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_923
timestamp 1679581782
transform 1 0 89760 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_930
timestamp 1679581782
transform 1 0 90432 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_937
timestamp 1679581782
transform 1 0 91104 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_944
timestamp 1679581782
transform 1 0 91776 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_951
timestamp 1679581782
transform 1 0 92448 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_958
timestamp 1679581782
transform 1 0 93120 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_965
timestamp 1679581782
transform 1 0 93792 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_972
timestamp 1679581782
transform 1 0 94464 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_979
timestamp 1679581782
transform 1 0 95136 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_986
timestamp 1679581782
transform 1 0 95808 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_993
timestamp 1679581782
transform 1 0 96480 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1000
timestamp 1679581782
transform 1 0 97152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1007
timestamp 1679581782
transform 1 0 97824 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1014
timestamp 1677580104
transform 1 0 98496 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_1016
timestamp 1677579658
transform 1 0 98688 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7872 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 8544 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_84
timestamp 1679577901
transform 1 0 9216 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679581782
transform 1 0 10368 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12576 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 13248 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13920 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_140
timestamp 1677580104
transform 1 0 14592 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_155
timestamp 1679581782
transform 1 0 16032 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_162
timestamp 1679581782
transform 1 0 16704 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_169
timestamp 1679581782
transform 1 0 17376 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_176
timestamp 1679577901
transform 1 0 18048 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_180
timestamp 1677579658
transform 1 0 18432 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_185
timestamp 1679581782
transform 1 0 18912 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_192
timestamp 1679581782
transform 1 0 19584 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_199
timestamp 1677580104
transform 1 0 20256 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_206
timestamp 1679581782
transform 1 0 20928 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_213
timestamp 1679581782
transform 1 0 21600 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_220
timestamp 1679581782
transform 1 0 22272 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_227
timestamp 1679581782
transform 1 0 22944 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_234
timestamp 1679577901
transform 1 0 23616 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_238
timestamp 1677579658
transform 1 0 24000 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_256
timestamp 1679581782
transform 1 0 25728 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_263
timestamp 1679581782
transform 1 0 26400 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_270
timestamp 1677580104
transform 1 0 27072 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_272
timestamp 1677579658
transform 1 0 27264 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_289
timestamp 1677580104
transform 1 0 28896 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_291
timestamp 1677579658
transform 1 0 29088 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_297
timestamp 1679581782
transform 1 0 29664 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_304
timestamp 1679581782
transform 1 0 30336 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_311
timestamp 1679577901
transform 1 0 31008 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_328
timestamp 1679581782
transform 1 0 32640 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_335
timestamp 1679577901
transform 1 0 33312 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_339
timestamp 1677580104
transform 1 0 33696 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_361
timestamp 1679581782
transform 1 0 35808 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_368
timestamp 1679577901
transform 1 0 36480 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_377
timestamp 1679581782
transform 1 0 37344 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_384
timestamp 1677580104
transform 1 0 38016 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_391
timestamp 1679581782
transform 1 0 38688 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_398
timestamp 1679581782
transform 1 0 39360 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_405
timestamp 1679581782
transform 1 0 40032 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_412
timestamp 1679581782
transform 1 0 40704 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_419
timestamp 1679581782
transform 1 0 41376 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_426
timestamp 1677580104
transform 1 0 42048 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_428
timestamp 1677579658
transform 1 0 42240 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_462
timestamp 1679577901
transform 1 0 45504 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_466
timestamp 1677580104
transform 1 0 45888 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_494
timestamp 1677579658
transform 1 0 48576 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_506
timestamp 1677579658
transform 1 0 49728 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679581782
transform 1 0 51552 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_532
timestamp 1677579658
transform 1 0 52224 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_540
timestamp 1679581782
transform 1 0 52992 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_547
timestamp 1679577901
transform 1 0 53664 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_551
timestamp 1677580104
transform 1 0 54048 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_567
timestamp 1677580104
transform 1 0 55584 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_569
timestamp 1677579658
transform 1 0 55776 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_574
timestamp 1677580104
transform 1 0 56256 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_576
timestamp 1677579658
transform 1 0 56448 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_587
timestamp 1679581782
transform 1 0 57504 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_594
timestamp 1679577901
transform 1 0 58176 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_598
timestamp 1677579658
transform 1 0 58560 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_603
timestamp 1677579658
transform 1 0 59040 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_617
timestamp 1679581782
transform 1 0 60384 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_624
timestamp 1679581782
transform 1 0 61056 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_631
timestamp 1679581782
transform 1 0 61728 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_638
timestamp 1679581782
transform 1 0 62400 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_645
timestamp 1679581782
transform 1 0 63072 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_652
timestamp 1679581782
transform 1 0 63744 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_659
timestamp 1679581782
transform 1 0 64416 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_666
timestamp 1679581782
transform 1 0 65088 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_673
timestamp 1679581782
transform 1 0 65760 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_680
timestamp 1679577901
transform 1 0 66432 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_684
timestamp 1677579658
transform 1 0 66816 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_690
timestamp 1679581782
transform 1 0 67392 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_697
timestamp 1679581782
transform 1 0 68064 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_704
timestamp 1679581782
transform 1 0 68736 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_711
timestamp 1679577901
transform 1 0 69408 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_715
timestamp 1677579658
transform 1 0 69792 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_720
timestamp 1677579658
transform 1 0 70272 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_729
timestamp 1679581782
transform 1 0 71136 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_736
timestamp 1679581782
transform 1 0 71808 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_743
timestamp 1679581782
transform 1 0 72480 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_754
timestamp 1679581782
transform 1 0 73536 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_761
timestamp 1677580104
transform 1 0 74208 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_763
timestamp 1677579658
transform 1 0 74400 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_776
timestamp 1677580104
transform 1 0 75648 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_783
timestamp 1677580104
transform 1 0 76320 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_785
timestamp 1677579658
transform 1 0 76512 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_790
timestamp 1679581782
transform 1 0 76992 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_797
timestamp 1677580104
transform 1 0 77664 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_811
timestamp 1679581782
transform 1 0 79008 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_818
timestamp 1679581782
transform 1 0 79680 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_825
timestamp 1679577901
transform 1 0 80352 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_845
timestamp 1679581782
transform 1 0 82272 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_852
timestamp 1677579658
transform 1 0 82944 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_861
timestamp 1677580104
transform 1 0 83808 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_867
timestamp 1679581782
transform 1 0 84384 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_874
timestamp 1679581782
transform 1 0 85056 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_881
timestamp 1679581782
transform 1 0 85728 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_888
timestamp 1679577901
transform 1 0 86400 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_908
timestamp 1679577901
transform 1 0 88320 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_912
timestamp 1677580104
transform 1 0 88704 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_922
timestamp 1679581782
transform 1 0 89664 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_929
timestamp 1679581782
transform 1 0 90336 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_936
timestamp 1679581782
transform 1 0 91008 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_943
timestamp 1679581782
transform 1 0 91680 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_950
timestamp 1679581782
transform 1 0 92352 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_957
timestamp 1679581782
transform 1 0 93024 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_964
timestamp 1679581782
transform 1 0 93696 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_971
timestamp 1679581782
transform 1 0 94368 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_978
timestamp 1679581782
transform 1 0 95040 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_985
timestamp 1679581782
transform 1 0 95712 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_992
timestamp 1679581782
transform 1 0 96384 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_999
timestamp 1679581782
transform 1 0 97056 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1006
timestamp 1679581782
transform 1 0 97728 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_1013
timestamp 1679577901
transform 1 0 98400 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_105
timestamp 1677580104
transform 1 0 11232 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_107
timestamp 1677579658
transform 1 0 11424 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_117
timestamp 1679581782
transform 1 0 12384 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_124
timestamp 1679581782
transform 1 0 13056 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_131
timestamp 1679581782
transform 1 0 13728 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_138
timestamp 1677579658
transform 1 0 14400 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_159
timestamp 1679581782
transform 1 0 16416 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_166
timestamp 1679581782
transform 1 0 17088 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_173
timestamp 1679581782
transform 1 0 17760 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_180
timestamp 1679577901
transform 1 0 18432 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_184
timestamp 1677579658
transform 1 0 18816 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_197
timestamp 1679581782
transform 1 0 20064 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_204
timestamp 1679581782
transform 1 0 20736 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_211
timestamp 1679581782
transform 1 0 21408 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_218
timestamp 1679581782
transform 1 0 22080 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_225
timestamp 1679581782
transform 1 0 22752 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_232
timestamp 1679581782
transform 1 0 23424 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_247
timestamp 1677580104
transform 1 0 24864 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_254
timestamp 1679581782
transform 1 0 25536 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_261
timestamp 1679581782
transform 1 0 26208 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_268
timestamp 1679581782
transform 1 0 26880 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_275
timestamp 1679581782
transform 1 0 27552 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_282
timestamp 1679581782
transform 1 0 28224 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_289
timestamp 1679581782
transform 1 0 28896 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_296
timestamp 1679577901
transform 1 0 29568 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_305
timestamp 1677579658
transform 1 0 30432 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_314
timestamp 1679581782
transform 1 0 31296 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_321
timestamp 1679581782
transform 1 0 31968 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_328
timestamp 1679581782
transform 1 0 32640 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_335
timestamp 1679581782
transform 1 0 33312 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_342
timestamp 1679577901
transform 1 0 33984 0 1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 35136 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_361
timestamp 1679577901
transform 1 0 35808 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_373
timestamp 1677579658
transform 1 0 36960 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_379
timestamp 1679577901
transform 1 0 37536 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_395
timestamp 1677580104
transform 1 0 39072 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_423
timestamp 1679577901
transform 1 0 41760 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_427
timestamp 1677579658
transform 1 0 42144 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 43488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 44160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 44832 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 45504 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 46176 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 46848 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 47520 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_508
timestamp 1679581782
transform 1 0 49920 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_515
timestamp 1679577901
transform 1 0 50592 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_519
timestamp 1677579658
transform 1 0 50976 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_547
timestamp 1679581782
transform 1 0 53664 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_554
timestamp 1679577901
transform 1 0 54336 0 1 9072
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_562
timestamp 1679577901
transform 1 0 55104 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_566
timestamp 1677580104
transform 1 0 55488 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_580
timestamp 1679581782
transform 1 0 56832 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_587
timestamp 1679581782
transform 1 0 57504 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_594
timestamp 1677580104
transform 1 0 58176 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_596
timestamp 1677579658
transform 1 0 58368 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_625
timestamp 1679581782
transform 1 0 61152 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_632
timestamp 1677579658
transform 1 0 61824 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_646
timestamp 1679581782
transform 1 0 63168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_653
timestamp 1679581782
transform 1 0 63840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_660
timestamp 1679577901
transform 1 0 64512 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_664
timestamp 1677579658
transform 1 0 64896 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_678
timestamp 1679581782
transform 1 0 66240 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_685
timestamp 1679581782
transform 1 0 66912 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_692
timestamp 1679581782
transform 1 0 67584 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_699
timestamp 1679581782
transform 1 0 68256 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_706
timestamp 1679581782
transform 1 0 68928 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_713
timestamp 1679581782
transform 1 0 69600 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_720
timestamp 1677580104
transform 1 0 70272 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_727
timestamp 1679577901
transform 1 0 70944 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_731
timestamp 1677580104
transform 1 0 71328 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_741
timestamp 1679581782
transform 1 0 72288 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_748
timestamp 1677579658
transform 1 0 72960 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_753
timestamp 1677580104
transform 1 0 73440 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_759
timestamp 1679581782
transform 1 0 74016 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_766
timestamp 1679581782
transform 1 0 74688 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_773
timestamp 1679581782
transform 1 0 75360 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_780
timestamp 1679581782
transform 1 0 76032 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_787
timestamp 1677580104
transform 1 0 76704 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_801
timestamp 1677580104
transform 1 0 78048 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_807
timestamp 1679577901
transform 1 0 78624 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_811
timestamp 1677579658
transform 1 0 79008 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_825
timestamp 1677580104
transform 1 0 80352 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_835
timestamp 1679577901
transform 1 0 81312 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_839
timestamp 1677579658
transform 1 0 81696 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_844
timestamp 1679581782
transform 1 0 82176 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_851
timestamp 1679581782
transform 1 0 82848 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_858
timestamp 1679581782
transform 1 0 83520 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_865
timestamp 1679581782
transform 1 0 84192 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_872
timestamp 1679581782
transform 1 0 84864 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_879
timestamp 1679581782
transform 1 0 85536 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_886
timestamp 1679581782
transform 1 0 86208 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_893
timestamp 1677580104
transform 1 0 86880 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_899
timestamp 1677580104
transform 1 0 87456 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_905
timestamp 1677579658
transform 1 0 88032 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_926
timestamp 1679581782
transform 1 0 90048 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_933
timestamp 1679581782
transform 1 0 90720 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_940
timestamp 1679581782
transform 1 0 91392 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_947
timestamp 1679581782
transform 1 0 92064 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_954
timestamp 1679581782
transform 1 0 92736 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_961
timestamp 1679581782
transform 1 0 93408 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_968
timestamp 1679581782
transform 1 0 94080 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_975
timestamp 1679581782
transform 1 0 94752 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_982
timestamp 1679581782
transform 1 0 95424 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_989
timestamp 1679581782
transform 1 0 96096 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_996
timestamp 1679581782
transform 1 0 96768 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1003
timestamp 1679581782
transform 1 0 97440 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1010
timestamp 1679581782
transform 1 0 98112 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 7200 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7872 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 8544 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 9216 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9888 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_98
timestamp 1677580104
transform 1 0 10560 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_124
timestamp 1679581782
transform 1 0 13056 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_131
timestamp 1679581782
transform 1 0 13728 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_138
timestamp 1677579658
transform 1 0 14400 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_159
timestamp 1679581782
transform 1 0 16416 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_166
timestamp 1679581782
transform 1 0 17088 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_173
timestamp 1679581782
transform 1 0 17760 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_180
timestamp 1677579658
transform 1 0 18432 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_201
timestamp 1679581782
transform 1 0 20448 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_208
timestamp 1677580104
transform 1 0 21120 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_216
timestamp 1679581782
transform 1 0 21888 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_223
timestamp 1679581782
transform 1 0 22560 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_230
timestamp 1679577901
transform 1 0 23232 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_234
timestamp 1677579658
transform 1 0 23616 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_247
timestamp 1677580104
transform 1 0 24864 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_255
timestamp 1679581782
transform 1 0 25632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_262
timestamp 1679581782
transform 1 0 26304 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_269
timestamp 1679581782
transform 1 0 26976 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_276
timestamp 1679581782
transform 1 0 27648 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_283
timestamp 1679581782
transform 1 0 28320 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_290
timestamp 1679581782
transform 1 0 28992 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_297
timestamp 1679577901
transform 1 0 29664 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_301
timestamp 1677579658
transform 1 0 30048 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_318
timestamp 1677580104
transform 1 0 31680 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 32448 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_333
timestamp 1679581782
transform 1 0 33120 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_340
timestamp 1679581782
transform 1 0 33792 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_347
timestamp 1679581782
transform 1 0 34464 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_354
timestamp 1679577901
transform 1 0 35136 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_374
timestamp 1677580104
transform 1 0 37056 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_376
timestamp 1677579658
transform 1 0 37248 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_397
timestamp 1679581782
transform 1 0 39264 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_404
timestamp 1679577901
transform 1 0 39936 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_408
timestamp 1677580104
transform 1 0 40320 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_436
timestamp 1679581782
transform 1 0 43008 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_443
timestamp 1679581782
transform 1 0 43680 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_450
timestamp 1679581782
transform 1 0 44352 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_457
timestamp 1679581782
transform 1 0 45024 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_464
timestamp 1679581782
transform 1 0 45696 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_471
timestamp 1679581782
transform 1 0 46368 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_478
timestamp 1679581782
transform 1 0 47040 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_485
timestamp 1679581782
transform 1 0 47712 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_492
timestamp 1679581782
transform 1 0 48384 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_499
timestamp 1677580104
transform 1 0 49056 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_514
timestamp 1679581782
transform 1 0 50496 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_521
timestamp 1679581782
transform 1 0 51168 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_528
timestamp 1677580104
transform 1 0 51840 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_543
timestamp 1679581782
transform 1 0 53280 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_550
timestamp 1679581782
transform 1 0 53952 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_557
timestamp 1679581782
transform 1 0 54624 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_564
timestamp 1679581782
transform 1 0 55296 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_571
timestamp 1679581782
transform 1 0 55968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_578
timestamp 1679581782
transform 1 0 56640 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_585
timestamp 1677580104
transform 1 0 57312 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_605
timestamp 1679577901
transform 1 0 59232 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_609
timestamp 1677580104
transform 1 0 59616 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_619
timestamp 1679581782
transform 1 0 60576 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_626
timestamp 1679581782
transform 1 0 61248 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_633
timestamp 1679581782
transform 1 0 61920 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_640
timestamp 1679581782
transform 1 0 62592 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_647
timestamp 1679581782
transform 1 0 63264 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_654
timestamp 1679581782
transform 1 0 63936 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_661
timestamp 1679581782
transform 1 0 64608 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_668
timestamp 1679581782
transform 1 0 65280 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_675
timestamp 1679581782
transform 1 0 65952 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_682
timestamp 1679581782
transform 1 0 66624 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_689
timestamp 1679581782
transform 1 0 67296 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_696
timestamp 1677580104
transform 1 0 67968 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_698
timestamp 1677579658
transform 1 0 68160 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_717
timestamp 1679581782
transform 1 0 69984 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_724
timestamp 1679577901
transform 1 0 70656 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_728
timestamp 1677580104
transform 1 0 71040 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_734
timestamp 1679581782
transform 1 0 71616 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_741
timestamp 1679577901
transform 1 0 72288 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_745
timestamp 1677580104
transform 1 0 72672 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_765
timestamp 1679581782
transform 1 0 74592 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_772
timestamp 1679581782
transform 1 0 75264 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_779
timestamp 1679577901
transform 1 0 75936 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_783
timestamp 1677579658
transform 1 0 76320 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_800
timestamp 1679581782
transform 1 0 77952 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679581782
transform 1 0 78624 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679581782
transform 1 0 79296 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_821
timestamp 1679581782
transform 1 0 79968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_828
timestamp 1679581782
transform 1 0 80640 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_835
timestamp 1679581782
transform 1 0 81312 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_842
timestamp 1679577901
transform 1 0 81984 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_846
timestamp 1677579658
transform 1 0 82368 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_851
timestamp 1677580104
transform 1 0 82848 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_853
timestamp 1677579658
transform 1 0 83040 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_866
timestamp 1679581782
transform 1 0 84288 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_873
timestamp 1679581782
transform 1 0 84960 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_880
timestamp 1679581782
transform 1 0 85632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_887
timestamp 1679581782
transform 1 0 86304 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_894
timestamp 1679581782
transform 1 0 86976 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_901
timestamp 1677579658
transform 1 0 87648 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_918
timestamp 1677579658
transform 1 0 89280 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_923
timestamp 1679581782
transform 1 0 89760 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_930
timestamp 1679581782
transform 1 0 90432 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_937
timestamp 1679581782
transform 1 0 91104 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_944
timestamp 1679581782
transform 1 0 91776 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_951
timestamp 1679581782
transform 1 0 92448 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_958
timestamp 1679581782
transform 1 0 93120 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_965
timestamp 1679581782
transform 1 0 93792 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_972
timestamp 1679581782
transform 1 0 94464 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_979
timestamp 1679581782
transform 1 0 95136 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_986
timestamp 1679581782
transform 1 0 95808 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_993
timestamp 1679581782
transform 1 0 96480 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1000
timestamp 1679581782
transform 1 0 97152 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1007
timestamp 1679581782
transform 1 0 97824 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_1014
timestamp 1677580104
transform 1 0 98496 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_1016
timestamp 1677579658
transform 1 0 98688 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 6528 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 7200 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7872 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 8544 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 10560 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_105
timestamp 1679577901
transform 1 0 11232 0 1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_109
timestamp 1677579658
transform 1 0 11616 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_118
timestamp 1679581782
transform 1 0 12480 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_125
timestamp 1679581782
transform 1 0 13152 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_132
timestamp 1679581782
transform 1 0 13824 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_139
timestamp 1679581782
transform 1 0 14496 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_146
timestamp 1679577901
transform 1 0 15168 0 1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679581782
transform 1 0 15936 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_161
timestamp 1679577901
transform 1 0 16608 0 1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_165
timestamp 1677580104
transform 1 0 16992 0 1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_172
timestamp 1679581782
transform 1 0 17664 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_179
timestamp 1679581782
transform 1 0 18336 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_186
timestamp 1679577901
transform 1 0 19008 0 1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_194
timestamp 1679581782
transform 1 0 19776 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_201
timestamp 1679581782
transform 1 0 20448 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_208
timestamp 1679581782
transform 1 0 21120 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_215
timestamp 1679581782
transform 1 0 21792 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_222
timestamp 1679581782
transform 1 0 22464 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_229
timestamp 1679581782
transform 1 0 23136 0 1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_236
timestamp 1677580104
transform 1 0 23808 0 1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_238
timestamp 1677579658
transform 1 0 24000 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_251
timestamp 1679581782
transform 1 0 25248 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_258
timestamp 1679581782
transform 1 0 25920 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_265
timestamp 1679581782
transform 1 0 26592 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_272
timestamp 1679581782
transform 1 0 27264 0 1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_279
timestamp 1677580104
transform 1 0 27936 0 1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_286
timestamp 1679581782
transform 1 0 28608 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_293
timestamp 1679581782
transform 1 0 29280 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_300
timestamp 1679581782
transform 1 0 29952 0 1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_307
timestamp 1677579658
transform 1 0 30624 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_316
timestamp 1679581782
transform 1 0 31488 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_323
timestamp 1679581782
transform 1 0 32160 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_330
timestamp 1679581782
transform 1 0 32832 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_337
timestamp 1679581782
transform 1 0 33504 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_344
timestamp 1679581782
transform 1 0 34176 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_351
timestamp 1679581782
transform 1 0 34848 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_358
timestamp 1679581782
transform 1 0 35520 0 1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_365
timestamp 1677580104
transform 1 0 36192 0 1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_375
timestamp 1679581782
transform 1 0 37152 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_382
timestamp 1679581782
transform 1 0 37824 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_389
timestamp 1679577901
transform 1 0 38496 0 1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_393
timestamp 1677580104
transform 1 0 38880 0 1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_400
timestamp 1679581782
transform 1 0 39552 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_407
timestamp 1679581782
transform 1 0 40224 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_414
timestamp 1679581782
transform 1 0 40896 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_421
timestamp 1679581782
transform 1 0 41568 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_428
timestamp 1679581782
transform 1 0 42240 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_435
timestamp 1679581782
transform 1 0 42912 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_442
timestamp 1679581782
transform 1 0 43584 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_449
timestamp 1679581782
transform 1 0 44256 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_456
timestamp 1679581782
transform 1 0 44928 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_463
timestamp 1679581782
transform 1 0 45600 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_470
timestamp 1679581782
transform 1 0 46272 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_477
timestamp 1679581782
transform 1 0 46944 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_484
timestamp 1679581782
transform 1 0 47616 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_491
timestamp 1679581782
transform 1 0 48288 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_498
timestamp 1679581782
transform 1 0 48960 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_505
timestamp 1679577901
transform 1 0 49632 0 1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_513
timestamp 1679581782
transform 1 0 50400 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_520
timestamp 1679581782
transform 1 0 51072 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_527
timestamp 1679581782
transform 1 0 51744 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_534
timestamp 1679581782
transform 1 0 52416 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_541
timestamp 1679581782
transform 1 0 53088 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_548
timestamp 1679581782
transform 1 0 53760 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_555
timestamp 1679581782
transform 1 0 54432 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_562
timestamp 1679581782
transform 1 0 55104 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_569
timestamp 1679581782
transform 1 0 55776 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_576
timestamp 1679581782
transform 1 0 56448 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_583
timestamp 1679581782
transform 1 0 57120 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_590
timestamp 1679581782
transform 1 0 57792 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_597
timestamp 1679581782
transform 1 0 58464 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_604
timestamp 1679581782
transform 1 0 59136 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_611
timestamp 1679581782
transform 1 0 59808 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_618
timestamp 1679577901
transform 1 0 60480 0 1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_622
timestamp 1677579658
transform 1 0 60864 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_628
timestamp 1679581782
transform 1 0 61440 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_635
timestamp 1679581782
transform 1 0 62112 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_642
timestamp 1679581782
transform 1 0 62784 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_649
timestamp 1679581782
transform 1 0 63456 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_656
timestamp 1679581782
transform 1 0 64128 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_663
timestamp 1679581782
transform 1 0 64800 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_670
timestamp 1679581782
transform 1 0 65472 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_677
timestamp 1679581782
transform 1 0 66144 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_684
timestamp 1679581782
transform 1 0 66816 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_691
timestamp 1679581782
transform 1 0 67488 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_698
timestamp 1679581782
transform 1 0 68160 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_705
timestamp 1679581782
transform 1 0 68832 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_712
timestamp 1679581782
transform 1 0 69504 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_719
timestamp 1679581782
transform 1 0 70176 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_726
timestamp 1679581782
transform 1 0 70848 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_733
timestamp 1679577901
transform 1 0 71520 0 1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_742
timestamp 1679581782
transform 1 0 72384 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_749
timestamp 1679581782
transform 1 0 73056 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_756
timestamp 1679581782
transform 1 0 73728 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_763
timestamp 1679581782
transform 1 0 74400 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_770
timestamp 1679581782
transform 1 0 75072 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_777
timestamp 1679581782
transform 1 0 75744 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_784
timestamp 1679581782
transform 1 0 76416 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_791
timestamp 1679581782
transform 1 0 77088 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_798
timestamp 1679581782
transform 1 0 77760 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_805
timestamp 1679581782
transform 1 0 78432 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_812
timestamp 1679581782
transform 1 0 79104 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_819
timestamp 1679581782
transform 1 0 79776 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_826
timestamp 1679581782
transform 1 0 80448 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_833
timestamp 1679581782
transform 1 0 81120 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_840
timestamp 1679581782
transform 1 0 81792 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_847
timestamp 1679577901
transform 1 0 82464 0 1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_856
timestamp 1679581782
transform 1 0 83328 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_863
timestamp 1679581782
transform 1 0 84000 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_870
timestamp 1679581782
transform 1 0 84672 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_877
timestamp 1679581782
transform 1 0 85344 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_884
timestamp 1679581782
transform 1 0 86016 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_891
timestamp 1679581782
transform 1 0 86688 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_898
timestamp 1679581782
transform 1 0 87360 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_905
timestamp 1679581782
transform 1 0 88032 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_912
timestamp 1679581782
transform 1 0 88704 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_919
timestamp 1679581782
transform 1 0 89376 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_926
timestamp 1679581782
transform 1 0 90048 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_933
timestamp 1679581782
transform 1 0 90720 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_940
timestamp 1679581782
transform 1 0 91392 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_947
timestamp 1679581782
transform 1 0 92064 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_954
timestamp 1679581782
transform 1 0 92736 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_961
timestamp 1679581782
transform 1 0 93408 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_968
timestamp 1679581782
transform 1 0 94080 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_975
timestamp 1679581782
transform 1 0 94752 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_982
timestamp 1679581782
transform 1 0 95424 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_989
timestamp 1679581782
transform 1 0 96096 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_996
timestamp 1679581782
transform 1 0 96768 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1003
timestamp 1679581782
transform 1 0 97440 0 1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1010
timestamp 1679581782
transform 1 0 98112 0 1 10584
box -48 -56 720 834
use sg13g2_buf_2  input1
timestamp 1676381867
transform -1 0 17664 0 1 10584
box -48 -56 528 834
use sg13g2_buf_2  input2
timestamp 1676381867
transform -1 0 28608 0 1 10584
box -48 -56 528 834
use sg13g2_buf_2  input3
timestamp 1676381867
transform -1 0 39552 0 1 10584
box -48 -56 528 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 50016 0 1 10584
box -48 -56 432 834
use sg13g2_buf_2  input5
timestamp 1676381867
transform -1 0 61440 0 1 10584
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1676381867
transform -1 0 72384 0 1 10584
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1676381867
transform -1 0 83328 0 1 10584
box -48 -56 528 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 1536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 37152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 37536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 37920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 40128 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 39456 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 40512 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 39840 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 39456 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 41280 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 40608 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 4128 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 40224 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 42816 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 41376 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 40992 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 43584 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 42144 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 42528 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 42912 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 43296 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 43296 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 4512 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 43680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform -1 0 47712 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform 1 0 47040 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform 1 0 47424 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform 1 0 47808 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform 1 0 48192 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform 1 0 48288 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform 1 0 49056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform 1 0 48288 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 51360 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform 1 0 4896 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform 1 0 50400 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 51552 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 52320 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 53664 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 54048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 54048 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 55392 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 56160 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 56544 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 56928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform 1 0 5280 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform -1 0 55872 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 57888 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform -1 0 57024 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 59040 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform -1 0 58944 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 59328 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform -1 0 57312 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 58848 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform -1 0 59232 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 59616 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 5664 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 60480 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform -1 0 60000 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform -1 0 62400 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform -1 0 60384 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 60768 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 63360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 63744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 62880 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 62592 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 62976 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform 1 0 6048 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 64032 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 65664 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 63744 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 65376 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 66432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 66816 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 67200 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 67584 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 67968 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 68352 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform 1 0 6432 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 67008 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 69120 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 69504 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 67968 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 69600 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 70656 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 69408 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 71424 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 71808 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 70272 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform 1 0 6816 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 72576 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 72960 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 73344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 73728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 74496 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 74208 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 73824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 75648 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 75360 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform -1 0 75744 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 7200 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform -1 0 77184 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform -1 0 77568 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform -1 0 77952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform -1 0 76416 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform -1 0 75840 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform -1 0 79104 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform -1 0 77184 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform -1 0 79872 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform -1 0 79488 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform -1 0 79008 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 7584 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform -1 0 2208 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform -1 0 80640 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform -1 0 80640 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform -1 0 80352 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform -1 0 82560 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform -1 0 82944 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform -1 0 83328 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform -1 0 80544 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform -1 0 82272 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform -1 0 84096 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform -1 0 84480 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform 1 0 7968 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform -1 0 84864 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform -1 0 85632 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform -1 0 86400 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform -1 0 86784 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform -1 0 87168 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform -1 0 85920 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform -1 0 87552 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform -1 0 86304 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform -1 0 87936 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform -1 0 86688 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform 1 0 8352 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform -1 0 88320 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform -1 0 87072 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 88704 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform -1 0 87456 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform -1 0 89088 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform -1 0 88704 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform -1 0 88224 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform -1 0 89856 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform -1 0 89472 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 89856 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform 1 0 8736 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform -1 0 90240 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform -1 0 90624 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform -1 0 91008 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform -1 0 91392 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform -1 0 91776 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform -1 0 92160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform -1 0 92544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform -1 0 92928 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform -1 0 93312 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform -1 0 93696 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform 1 0 9120 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output164
timestamp 1676381911
transform -1 0 94080 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output165
timestamp 1676381911
transform -1 0 94464 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output166
timestamp 1676381911
transform -1 0 94848 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output167
timestamp 1676381911
transform -1 0 95232 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output168
timestamp 1676381911
transform -1 0 95616 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output169
timestamp 1676381911
transform -1 0 96000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output170
timestamp 1676381911
transform -1 0 96384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output171
timestamp 1676381911
transform -1 0 96768 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output172
timestamp 1676381911
transform -1 0 97152 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output173
timestamp 1676381911
transform -1 0 97536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output174
timestamp 1676381911
transform 1 0 9504 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output175
timestamp 1676381911
transform -1 0 97920 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output176
timestamp 1676381911
transform -1 0 98304 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output177
timestamp 1676381911
transform -1 0 98688 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output178
timestamp 1676381911
transform -1 0 98592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output179
timestamp 1676381911
transform 1 0 97824 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output180
timestamp 1676381911
transform 1 0 97056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output181
timestamp 1676381911
transform 1 0 9888 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output182
timestamp 1676381911
transform 1 0 10272 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output183
timestamp 1676381911
transform 1 0 10656 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output184
timestamp 1676381911
transform 1 0 11040 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output185
timestamp 1676381911
transform 1 0 11424 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output186
timestamp 1676381911
transform -1 0 1824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output187
timestamp 1676381911
transform 1 0 11808 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output188
timestamp 1676381911
transform 1 0 12192 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output189
timestamp 1676381911
transform 1 0 12576 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output190
timestamp 1676381911
transform -1 0 13824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output191
timestamp 1676381911
transform 1 0 12288 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output192
timestamp 1676381911
transform 1 0 13344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output193
timestamp 1676381911
transform 1 0 14208 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output194
timestamp 1676381911
transform 1 0 13056 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output195
timestamp 1676381911
transform 1 0 14112 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output196
timestamp 1676381911
transform 1 0 14976 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output197
timestamp 1676381911
transform 1 0 1440 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output198
timestamp 1676381911
transform 1 0 13824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output199
timestamp 1676381911
transform 1 0 14880 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output200
timestamp 1676381911
transform 1 0 15264 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output201
timestamp 1676381911
transform 1 0 16320 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output202
timestamp 1676381911
transform 1 0 14976 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output203
timestamp 1676381911
transform 1 0 16032 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output204
timestamp 1676381911
transform 1 0 17664 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output205
timestamp 1676381911
transform 1 0 15744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output206
timestamp 1676381911
transform -1 0 19584 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output207
timestamp 1676381911
transform 1 0 16896 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output208
timestamp 1676381911
transform 1 0 1824 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output209
timestamp 1676381911
transform 1 0 17280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output210
timestamp 1676381911
transform -1 0 20832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output211
timestamp 1676381911
transform -1 0 21216 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output212
timestamp 1676381911
transform 1 0 20928 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output213
timestamp 1676381911
transform 1 0 18816 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output214
timestamp 1676381911
transform 1 0 19200 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output215
timestamp 1676381911
transform 1 0 19584 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output216
timestamp 1676381911
transform 1 0 21408 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output217
timestamp 1676381911
transform 1 0 20352 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output218
timestamp 1676381911
transform 1 0 21120 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output219
timestamp 1676381911
transform 1 0 2208 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output220
timestamp 1676381911
transform 1 0 21888 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output221
timestamp 1676381911
transform 1 0 23712 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output222
timestamp 1676381911
transform 1 0 23328 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output223
timestamp 1676381911
transform 1 0 23040 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output224
timestamp 1676381911
transform 1 0 23808 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output225
timestamp 1676381911
transform 1 0 24192 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output226
timestamp 1676381911
transform 1 0 26016 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output227
timestamp 1676381911
transform 1 0 25632 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output228
timestamp 1676381911
transform 1 0 24960 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output229
timestamp 1676381911
transform 1 0 26784 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output230
timestamp 1676381911
transform 1 0 2592 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output231
timestamp 1676381911
transform 1 0 26400 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output232
timestamp 1676381911
transform 1 0 25728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output233
timestamp 1676381911
transform 1 0 26784 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output234
timestamp 1676381911
transform 1 0 26496 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output235
timestamp 1676381911
transform -1 0 29664 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output236
timestamp 1676381911
transform -1 0 30048 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output237
timestamp 1676381911
transform 1 0 29088 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output238
timestamp 1676381911
transform 1 0 28704 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output239
timestamp 1676381911
transform 1 0 28032 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output240
timestamp 1676381911
transform 1 0 28416 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output241
timestamp 1676381911
transform 1 0 2976 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output242
timestamp 1676381911
transform 1 0 29184 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output243
timestamp 1676381911
transform 1 0 29952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output244
timestamp 1676381911
transform 1 0 31392 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output245
timestamp 1676381911
transform 1 0 30720 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output246
timestamp 1676381911
transform 1 0 32544 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output247
timestamp 1676381911
transform 1 0 32160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output248
timestamp 1676381911
transform 1 0 33696 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output249
timestamp 1676381911
transform 1 0 32544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output250
timestamp 1676381911
transform 1 0 31872 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output251
timestamp 1676381911
transform 1 0 33696 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output252
timestamp 1676381911
transform 1 0 3360 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output253
timestamp 1676381911
transform -1 0 35808 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output254
timestamp 1676381911
transform 1 0 34080 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output255
timestamp 1676381911
transform 1 0 33024 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output256
timestamp 1676381911
transform 1 0 33792 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output257
timestamp 1676381911
transform 1 0 35232 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output258
timestamp 1676381911
transform 1 0 37056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output259
timestamp 1676381911
transform 1 0 36384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output260
timestamp 1676381911
transform 1 0 36000 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output261
timestamp 1676381911
transform 1 0 37824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output262
timestamp 1676381911
transform 1 0 37152 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output263
timestamp 1676381911
transform 1 0 3744 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output264
timestamp 1676381911
transform -1 0 2976 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output265
timestamp 1676381911
transform -1 0 39840 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output266
timestamp 1676381911
transform -1 0 40224 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output267
timestamp 1676381911
transform 1 0 38304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output268
timestamp 1676381911
transform 1 0 38688 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output269
timestamp 1676381911
transform -1 0 41376 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output270
timestamp 1676381911
transform 1 0 39072 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output271
timestamp 1676381911
transform 1 0 40896 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output272
timestamp 1676381911
transform 1 0 40224 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output273
timestamp 1676381911
transform 1 0 39840 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output274
timestamp 1676381911
transform 1 0 41664 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output275
timestamp 1676381911
transform 1 0 3456 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output276
timestamp 1676381911
transform 1 0 40992 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output277
timestamp 1676381911
transform 1 0 40608 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output278
timestamp 1676381911
transform 1 0 43200 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output279
timestamp 1676381911
transform 1 0 41760 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output280
timestamp 1676381911
transform 1 0 41376 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output281
timestamp 1676381911
transform 1 0 41760 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output282
timestamp 1676381911
transform 1 0 42144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output283
timestamp 1676381911
transform 1 0 42528 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output284
timestamp 1676381911
transform 1 0 42912 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output285
timestamp 1676381911
transform 1 0 46560 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output286
timestamp 1676381911
transform 1 0 3840 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output287
timestamp 1676381911
transform 1 0 44064 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output288
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output289
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output290
timestamp 1676381911
transform 1 0 45216 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output291
timestamp 1676381911
transform 1 0 45600 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output292
timestamp 1676381911
transform 1 0 47904 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output293
timestamp 1676381911
transform 1 0 48672 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output294
timestamp 1676381911
transform 1 0 47904 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output295
timestamp 1676381911
transform 1 0 48672 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output296
timestamp 1676381911
transform -1 0 50976 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output297
timestamp 1676381911
transform 1 0 4224 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output298
timestamp 1676381911
transform 1 0 50784 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output299
timestamp 1676381911
transform -1 0 51936 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output300
timestamp 1676381911
transform -1 0 53280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output301
timestamp 1676381911
transform -1 0 52512 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output302
timestamp 1676381911
transform -1 0 54432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output303
timestamp 1676381911
transform -1 0 54432 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output304
timestamp 1676381911
transform -1 0 55776 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output305
timestamp 1676381911
transform -1 0 55776 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output306
timestamp 1676381911
transform -1 0 56160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output307
timestamp 1676381911
transform -1 0 55008 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output308
timestamp 1676381911
transform 1 0 4608 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output309
timestamp 1676381911
transform -1 0 55392 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output310
timestamp 1676381911
transform -1 0 58272 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output311
timestamp 1676381911
transform -1 0 58656 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output312
timestamp 1676381911
transform -1 0 56352 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output313
timestamp 1676381911
transform -1 0 56736 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output314
timestamp 1676381911
transform -1 0 60864 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output315
timestamp 1676381911
transform -1 0 58080 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output316
timestamp 1676381911
transform -1 0 61248 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output317
timestamp 1676381911
transform -1 0 61632 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output318
timestamp 1676381911
transform -1 0 58944 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output319
timestamp 1676381911
transform 1 0 4992 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output320
timestamp 1676381911
transform -1 0 62016 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output321
timestamp 1676381911
transform -1 0 60864 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output322
timestamp 1676381911
transform -1 0 61728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output323
timestamp 1676381911
transform -1 0 62112 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output324
timestamp 1676381911
transform -1 0 62496 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output325
timestamp 1676381911
transform -1 0 62880 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output326
timestamp 1676381911
transform -1 0 64128 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output327
timestamp 1676381911
transform -1 0 64512 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output328
timestamp 1676381911
transform -1 0 64896 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output329
timestamp 1676381911
transform -1 0 65280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output330
timestamp 1676381911
transform 1 0 5376 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output331
timestamp 1676381911
transform -1 0 63360 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output332
timestamp 1676381911
transform -1 0 64416 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output333
timestamp 1676381911
transform -1 0 66048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output334
timestamp 1676381911
transform -1 0 64128 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output335
timestamp 1676381911
transform -1 0 65760 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output336
timestamp 1676381911
transform -1 0 66144 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output337
timestamp 1676381911
transform -1 0 66528 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output338
timestamp 1676381911
transform -1 0 66240 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output339
timestamp 1676381911
transform -1 0 66624 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output340
timestamp 1676381911
transform -1 0 67680 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output341
timestamp 1676381911
transform 1 0 5760 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output342
timestamp 1676381911
transform -1 0 68736 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output343
timestamp 1676381911
transform -1 0 67104 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output344
timestamp 1676381911
transform -1 0 69888 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output345
timestamp 1676381911
transform -1 0 70272 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output346
timestamp 1676381911
transform -1 0 69024 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output347
timestamp 1676381911
transform -1 0 69984 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output348
timestamp 1676381911
transform -1 0 71040 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output349
timestamp 1676381911
transform -1 0 69408 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output350
timestamp 1676381911
transform -1 0 72192 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output351
timestamp 1676381911
transform -1 0 71040 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output352
timestamp 1676381911
transform 1 0 6144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output353
timestamp 1676381911
transform -1 0 70656 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output354
timestamp 1676381911
transform -1 0 71040 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output355
timestamp 1676381911
transform -1 0 72672 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output356
timestamp 1676381911
transform -1 0 74112 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output357
timestamp 1676381911
transform -1 0 74880 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output358
timestamp 1676381911
transform -1 0 75264 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output359
timestamp 1676381911
transform -1 0 74592 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output360
timestamp 1676381911
transform -1 0 76032 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output361
timestamp 1676381911
transform -1 0 76416 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output362
timestamp 1676381911
transform -1 0 76800 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output363
timestamp 1676381911
transform 1 0 6528 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output364
timestamp 1676381911
transform -1 0 76512 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output365
timestamp 1676381911
transform -1 0 75648 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output366
timestamp 1676381911
transform -1 0 78336 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output367
timestamp 1676381911
transform -1 0 78720 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output368
timestamp 1676381911
transform -1 0 76800 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output369
timestamp 1676381911
transform -1 0 77664 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output370
timestamp 1676381911
transform -1 0 79488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output371
timestamp 1676381911
transform -1 0 78624 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output372
timestamp 1676381911
transform -1 0 80256 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output373
timestamp 1676381911
transform -1 0 79872 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output374
timestamp 1676381911
transform 1 0 6912 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output375
timestamp 1676381911
transform -1 0 1824 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output376
timestamp 1676381911
transform -1 0 80256 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output377
timestamp 1676381911
transform -1 0 79968 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output378
timestamp 1676381911
transform -1 0 80736 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output379
timestamp 1676381911
transform -1 0 79776 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output380
timestamp 1676381911
transform -1 0 80160 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output381
timestamp 1676381911
transform -1 0 82752 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output382
timestamp 1676381911
transform -1 0 83712 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output383
timestamp 1676381911
transform -1 0 83136 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output384
timestamp 1676381911
transform -1 0 82656 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output385
timestamp 1676381911
transform -1 0 83904 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output386
timestamp 1676381911
transform 1 0 7296 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output387
timestamp 1676381911
transform -1 0 82080 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output388
timestamp 1676381911
transform -1 0 86016 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output389
timestamp 1676381911
transform -1 0 86016 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output390
timestamp 1676381911
transform -1 0 86400 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output391
timestamp 1676381911
transform -1 0 85152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output392
timestamp 1676381911
transform -1 0 86784 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output393
timestamp 1676381911
transform -1 0 85536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output394
timestamp 1676381911
transform -1 0 87168 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output395
timestamp 1676381911
transform -1 0 85920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output396
timestamp 1676381911
transform -1 0 87552 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output397
timestamp 1676381911
transform 1 0 7680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output398
timestamp 1676381911
transform -1 0 86304 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output399
timestamp 1676381911
transform -1 0 87936 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output400
timestamp 1676381911
transform -1 0 86688 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output401
timestamp 1676381911
transform -1 0 88320 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output402
timestamp 1676381911
transform -1 0 87840 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output403
timestamp 1676381911
transform -1 0 89472 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output404
timestamp 1676381911
transform -1 0 89088 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output405
timestamp 1676381911
transform -1 0 88608 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output406
timestamp 1676381911
transform -1 0 90240 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output407
timestamp 1676381911
transform -1 0 90624 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output408
timestamp 1676381911
transform 1 0 8064 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output409
timestamp 1676381911
transform -1 0 91008 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output410
timestamp 1676381911
transform -1 0 91392 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output411
timestamp 1676381911
transform -1 0 91776 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output412
timestamp 1676381911
transform -1 0 92160 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output413
timestamp 1676381911
transform -1 0 92544 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output414
timestamp 1676381911
transform -1 0 92928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output415
timestamp 1676381911
transform -1 0 93312 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output416
timestamp 1676381911
transform -1 0 93696 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output417
timestamp 1676381911
transform -1 0 94080 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output418
timestamp 1676381911
transform -1 0 94464 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output419
timestamp 1676381911
transform 1 0 8448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output420
timestamp 1676381911
transform -1 0 94848 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output421
timestamp 1676381911
transform -1 0 95232 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output422
timestamp 1676381911
transform -1 0 95616 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output423
timestamp 1676381911
transform -1 0 96000 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output424
timestamp 1676381911
transform -1 0 96384 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output425
timestamp 1676381911
transform -1 0 96768 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output426
timestamp 1676381911
transform -1 0 97152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output427
timestamp 1676381911
transform -1 0 97536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output428
timestamp 1676381911
transform -1 0 97920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output429
timestamp 1676381911
transform -1 0 98304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output430
timestamp 1676381911
transform 1 0 8832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output431
timestamp 1676381911
transform -1 0 98688 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output432
timestamp 1676381911
transform -1 0 97824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output433
timestamp 1676381911
transform -1 0 98208 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output434
timestamp 1676381911
transform -1 0 98592 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output435
timestamp 1676381911
transform 1 0 98400 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output436
timestamp 1676381911
transform 1 0 97440 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output437
timestamp 1676381911
transform 1 0 9216 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output438
timestamp 1676381911
transform 1 0 9600 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output439
timestamp 1676381911
transform 1 0 9984 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output440
timestamp 1676381911
transform 1 0 10368 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output441
timestamp 1676381911
transform 1 0 10752 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output442
timestamp 1676381911
transform -1 0 2208 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output443
timestamp 1676381911
transform 1 0 11136 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output444
timestamp 1676381911
transform 1 0 11520 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output445
timestamp 1676381911
transform 1 0 11904 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output446
timestamp 1676381911
transform 1 0 12960 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output447
timestamp 1676381911
transform 1 0 13824 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output448
timestamp 1676381911
transform 1 0 12672 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output449
timestamp 1676381911
transform 1 0 13728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output450
timestamp 1676381911
transform 1 0 14592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output451
timestamp 1676381911
transform 1 0 13440 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output452
timestamp 1676381911
transform 1 0 14496 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output453
timestamp 1676381911
transform -1 0 2592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output454
timestamp 1676381911
transform 1 0 15360 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output455
timestamp 1676381911
transform 1 0 14208 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output456
timestamp 1676381911
transform 1 0 14592 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output457
timestamp 1676381911
transform 1 0 15648 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output458
timestamp 1676381911
transform 1 0 16704 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output459
timestamp 1676381911
transform 1 0 15360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output460
timestamp 1676381911
transform 1 0 16416 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output461
timestamp 1676381911
transform 1 0 16128 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output462
timestamp 1676381911
transform 1 0 16512 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output463
timestamp 1676381911
transform 1 0 17664 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output464
timestamp 1676381911
transform 1 0 1152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output465
timestamp 1676381911
transform 1 0 18048 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output466
timestamp 1676381911
transform 1 0 18432 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output467
timestamp 1676381911
transform 1 0 18432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output468
timestamp 1676381911
transform 1 0 20256 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output469
timestamp 1676381911
transform 1 0 21312 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output470
timestamp 1676381911
transform 1 0 20256 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output471
timestamp 1676381911
transform 1 0 20640 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output472
timestamp 1676381911
transform 1 0 19968 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output473
timestamp 1676381911
transform 1 0 20736 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output474
timestamp 1676381911
transform 1 0 21504 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output475
timestamp 1676381911
transform 1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output476
timestamp 1676381911
transform 1 0 22944 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output477
timestamp 1676381911
transform 1 0 22272 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output478
timestamp 1676381911
transform 1 0 22656 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output479
timestamp 1676381911
transform 1 0 23424 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output480
timestamp 1676381911
transform -1 0 26016 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output481
timestamp 1676381911
transform 1 0 25248 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output482
timestamp 1676381911
transform 1 0 24576 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output483
timestamp 1676381911
transform 1 0 26400 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output484
timestamp 1676381911
transform 1 0 26016 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output485
timestamp 1676381911
transform 1 0 25344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output486
timestamp 1676381911
transform 1 0 1920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output487
timestamp 1676381911
transform 1 0 27168 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output488
timestamp 1676381911
transform 1 0 28032 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output489
timestamp 1676381911
transform 1 0 26112 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output490
timestamp 1676381911
transform 1 0 26880 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output491
timestamp 1676381911
transform 1 0 27264 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output492
timestamp 1676381911
transform 1 0 28320 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output493
timestamp 1676381911
transform 1 0 27648 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output494
timestamp 1676381911
transform 1 0 29472 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output495
timestamp 1676381911
transform 1 0 29856 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output496
timestamp 1676381911
transform 1 0 28800 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output497
timestamp 1676381911
transform 1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output498
timestamp 1676381911
transform 1 0 29568 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output499
timestamp 1676381911
transform 1 0 30336 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output500
timestamp 1676381911
transform 1 0 32160 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output501
timestamp 1676381911
transform 1 0 31776 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output502
timestamp 1676381911
transform 1 0 31104 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output503
timestamp 1676381911
transform 1 0 32928 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output504
timestamp 1676381911
transform 1 0 31488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output505
timestamp 1676381911
transform 1 0 33312 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output506
timestamp 1676381911
transform 1 0 32928 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output507
timestamp 1676381911
transform 1 0 32256 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output508
timestamp 1676381911
transform 1 0 2688 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output509
timestamp 1676381911
transform 1 0 33312 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output510
timestamp 1676381911
transform 1 0 32640 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output511
timestamp 1676381911
transform 1 0 33408 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output512
timestamp 1676381911
transform 1 0 34176 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output513
timestamp 1676381911
transform 1 0 36000 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output514
timestamp 1676381911
transform 1 0 35616 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output515
timestamp 1676381911
transform 1 0 37440 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output516
timestamp 1676381911
transform 1 0 36768 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output517
timestamp 1676381911
transform 1 0 36384 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output518
timestamp 1676381911
transform 1 0 36768 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output519
timestamp 1676381911
transform 1 0 3072 0 1 3024
box -48 -56 432 834
<< labels >>
flabel metal6 s 4892 2898 5332 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 20012 2898 20452 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 35132 2898 35572 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 50252 2898 50692 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 65372 2898 65812 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 80492 2898 80932 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95612 2898 96052 11384 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 1108 6764 98828 7204 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3652 2980 4092 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18772 2980 19212 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33892 2980 34332 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 49012 2980 49452 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 64132 2980 64572 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 79252 2980 79692 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 94372 2980 94812 11466 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 1108 5524 98828 5964 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6200 14920 6280 15000 0 FreeSans 320 0 0 0 ena_i
port 2 nsew signal input
flabel metal2 s 17144 14920 17224 15000 0 FreeSans 320 0 0 0 input_ni[0]
port 3 nsew signal input
flabel metal2 s 28088 14920 28168 15000 0 FreeSans 320 0 0 0 input_ni[1]
port 4 nsew signal input
flabel metal2 s 39032 14920 39112 15000 0 FreeSans 320 0 0 0 input_ni[2]
port 5 nsew signal input
flabel metal2 s 49976 14920 50056 15000 0 FreeSans 320 0 0 0 input_ni[3]
port 6 nsew signal input
flabel metal2 s 60920 14920 61000 15000 0 FreeSans 320 0 0 0 input_ni[4]
port 7 nsew signal input
flabel metal2 s 71864 14920 71944 15000 0 FreeSans 320 0 0 0 input_ni[5]
port 8 nsew signal input
flabel metal2 s 82808 14920 82888 15000 0 FreeSans 320 0 0 0 input_ni[6]
port 9 nsew signal input
flabel metal2 s 93752 14920 93832 15000 0 FreeSans 320 0 0 0 input_ni[7]
port 10 nsew signal input
flabel metal2 s 824 0 904 80 0 FreeSans 320 0 0 0 output_no[0]
port 11 nsew signal output
flabel metal2 s 39224 0 39304 80 0 FreeSans 320 0 0 0 output_no[100]
port 12 nsew signal output
flabel metal2 s 39608 0 39688 80 0 FreeSans 320 0 0 0 output_no[101]
port 13 nsew signal output
flabel metal2 s 39992 0 40072 80 0 FreeSans 320 0 0 0 output_no[102]
port 14 nsew signal output
flabel metal2 s 40376 0 40456 80 0 FreeSans 320 0 0 0 output_no[103]
port 15 nsew signal output
flabel metal2 s 40760 0 40840 80 0 FreeSans 320 0 0 0 output_no[104]
port 16 nsew signal output
flabel metal2 s 41144 0 41224 80 0 FreeSans 320 0 0 0 output_no[105]
port 17 nsew signal output
flabel metal2 s 41528 0 41608 80 0 FreeSans 320 0 0 0 output_no[106]
port 18 nsew signal output
flabel metal2 s 41912 0 41992 80 0 FreeSans 320 0 0 0 output_no[107]
port 19 nsew signal output
flabel metal2 s 42296 0 42376 80 0 FreeSans 320 0 0 0 output_no[108]
port 20 nsew signal output
flabel metal2 s 42680 0 42760 80 0 FreeSans 320 0 0 0 output_no[109]
port 21 nsew signal output
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 output_no[10]
port 22 nsew signal output
flabel metal2 s 43064 0 43144 80 0 FreeSans 320 0 0 0 output_no[110]
port 23 nsew signal output
flabel metal2 s 43448 0 43528 80 0 FreeSans 320 0 0 0 output_no[111]
port 24 nsew signal output
flabel metal2 s 43832 0 43912 80 0 FreeSans 320 0 0 0 output_no[112]
port 25 nsew signal output
flabel metal2 s 44216 0 44296 80 0 FreeSans 320 0 0 0 output_no[113]
port 26 nsew signal output
flabel metal2 s 44600 0 44680 80 0 FreeSans 320 0 0 0 output_no[114]
port 27 nsew signal output
flabel metal2 s 44984 0 45064 80 0 FreeSans 320 0 0 0 output_no[115]
port 28 nsew signal output
flabel metal2 s 45368 0 45448 80 0 FreeSans 320 0 0 0 output_no[116]
port 29 nsew signal output
flabel metal2 s 45752 0 45832 80 0 FreeSans 320 0 0 0 output_no[117]
port 30 nsew signal output
flabel metal2 s 46136 0 46216 80 0 FreeSans 320 0 0 0 output_no[118]
port 31 nsew signal output
flabel metal2 s 46520 0 46600 80 0 FreeSans 320 0 0 0 output_no[119]
port 32 nsew signal output
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 output_no[11]
port 33 nsew signal output
flabel metal2 s 46904 0 46984 80 0 FreeSans 320 0 0 0 output_no[120]
port 34 nsew signal output
flabel metal2 s 47288 0 47368 80 0 FreeSans 320 0 0 0 output_no[121]
port 35 nsew signal output
flabel metal2 s 47672 0 47752 80 0 FreeSans 320 0 0 0 output_no[122]
port 36 nsew signal output
flabel metal2 s 48056 0 48136 80 0 FreeSans 320 0 0 0 output_no[123]
port 37 nsew signal output
flabel metal2 s 48440 0 48520 80 0 FreeSans 320 0 0 0 output_no[124]
port 38 nsew signal output
flabel metal2 s 48824 0 48904 80 0 FreeSans 320 0 0 0 output_no[125]
port 39 nsew signal output
flabel metal2 s 49208 0 49288 80 0 FreeSans 320 0 0 0 output_no[126]
port 40 nsew signal output
flabel metal2 s 49592 0 49672 80 0 FreeSans 320 0 0 0 output_no[127]
port 41 nsew signal output
flabel metal2 s 49976 0 50056 80 0 FreeSans 320 0 0 0 output_no[128]
port 42 nsew signal output
flabel metal2 s 50360 0 50440 80 0 FreeSans 320 0 0 0 output_no[129]
port 43 nsew signal output
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 output_no[12]
port 44 nsew signal output
flabel metal2 s 50744 0 50824 80 0 FreeSans 320 0 0 0 output_no[130]
port 45 nsew signal output
flabel metal2 s 51128 0 51208 80 0 FreeSans 320 0 0 0 output_no[131]
port 46 nsew signal output
flabel metal2 s 51512 0 51592 80 0 FreeSans 320 0 0 0 output_no[132]
port 47 nsew signal output
flabel metal2 s 51896 0 51976 80 0 FreeSans 320 0 0 0 output_no[133]
port 48 nsew signal output
flabel metal2 s 52280 0 52360 80 0 FreeSans 320 0 0 0 output_no[134]
port 49 nsew signal output
flabel metal2 s 52664 0 52744 80 0 FreeSans 320 0 0 0 output_no[135]
port 50 nsew signal output
flabel metal2 s 53048 0 53128 80 0 FreeSans 320 0 0 0 output_no[136]
port 51 nsew signal output
flabel metal2 s 53432 0 53512 80 0 FreeSans 320 0 0 0 output_no[137]
port 52 nsew signal output
flabel metal2 s 53816 0 53896 80 0 FreeSans 320 0 0 0 output_no[138]
port 53 nsew signal output
flabel metal2 s 54200 0 54280 80 0 FreeSans 320 0 0 0 output_no[139]
port 54 nsew signal output
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 output_no[13]
port 55 nsew signal output
flabel metal2 s 54584 0 54664 80 0 FreeSans 320 0 0 0 output_no[140]
port 56 nsew signal output
flabel metal2 s 54968 0 55048 80 0 FreeSans 320 0 0 0 output_no[141]
port 57 nsew signal output
flabel metal2 s 55352 0 55432 80 0 FreeSans 320 0 0 0 output_no[142]
port 58 nsew signal output
flabel metal2 s 55736 0 55816 80 0 FreeSans 320 0 0 0 output_no[143]
port 59 nsew signal output
flabel metal2 s 56120 0 56200 80 0 FreeSans 320 0 0 0 output_no[144]
port 60 nsew signal output
flabel metal2 s 56504 0 56584 80 0 FreeSans 320 0 0 0 output_no[145]
port 61 nsew signal output
flabel metal2 s 56888 0 56968 80 0 FreeSans 320 0 0 0 output_no[146]
port 62 nsew signal output
flabel metal2 s 57272 0 57352 80 0 FreeSans 320 0 0 0 output_no[147]
port 63 nsew signal output
flabel metal2 s 57656 0 57736 80 0 FreeSans 320 0 0 0 output_no[148]
port 64 nsew signal output
flabel metal2 s 58040 0 58120 80 0 FreeSans 320 0 0 0 output_no[149]
port 65 nsew signal output
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 output_no[14]
port 66 nsew signal output
flabel metal2 s 58424 0 58504 80 0 FreeSans 320 0 0 0 output_no[150]
port 67 nsew signal output
flabel metal2 s 58808 0 58888 80 0 FreeSans 320 0 0 0 output_no[151]
port 68 nsew signal output
flabel metal2 s 59192 0 59272 80 0 FreeSans 320 0 0 0 output_no[152]
port 69 nsew signal output
flabel metal2 s 59576 0 59656 80 0 FreeSans 320 0 0 0 output_no[153]
port 70 nsew signal output
flabel metal2 s 59960 0 60040 80 0 FreeSans 320 0 0 0 output_no[154]
port 71 nsew signal output
flabel metal2 s 60344 0 60424 80 0 FreeSans 320 0 0 0 output_no[155]
port 72 nsew signal output
flabel metal2 s 60728 0 60808 80 0 FreeSans 320 0 0 0 output_no[156]
port 73 nsew signal output
flabel metal2 s 61112 0 61192 80 0 FreeSans 320 0 0 0 output_no[157]
port 74 nsew signal output
flabel metal2 s 61496 0 61576 80 0 FreeSans 320 0 0 0 output_no[158]
port 75 nsew signal output
flabel metal2 s 61880 0 61960 80 0 FreeSans 320 0 0 0 output_no[159]
port 76 nsew signal output
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 output_no[15]
port 77 nsew signal output
flabel metal2 s 62264 0 62344 80 0 FreeSans 320 0 0 0 output_no[160]
port 78 nsew signal output
flabel metal2 s 62648 0 62728 80 0 FreeSans 320 0 0 0 output_no[161]
port 79 nsew signal output
flabel metal2 s 63032 0 63112 80 0 FreeSans 320 0 0 0 output_no[162]
port 80 nsew signal output
flabel metal2 s 63416 0 63496 80 0 FreeSans 320 0 0 0 output_no[163]
port 81 nsew signal output
flabel metal2 s 63800 0 63880 80 0 FreeSans 320 0 0 0 output_no[164]
port 82 nsew signal output
flabel metal2 s 64184 0 64264 80 0 FreeSans 320 0 0 0 output_no[165]
port 83 nsew signal output
flabel metal2 s 64568 0 64648 80 0 FreeSans 320 0 0 0 output_no[166]
port 84 nsew signal output
flabel metal2 s 64952 0 65032 80 0 FreeSans 320 0 0 0 output_no[167]
port 85 nsew signal output
flabel metal2 s 65336 0 65416 80 0 FreeSans 320 0 0 0 output_no[168]
port 86 nsew signal output
flabel metal2 s 65720 0 65800 80 0 FreeSans 320 0 0 0 output_no[169]
port 87 nsew signal output
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 output_no[16]
port 88 nsew signal output
flabel metal2 s 66104 0 66184 80 0 FreeSans 320 0 0 0 output_no[170]
port 89 nsew signal output
flabel metal2 s 66488 0 66568 80 0 FreeSans 320 0 0 0 output_no[171]
port 90 nsew signal output
flabel metal2 s 66872 0 66952 80 0 FreeSans 320 0 0 0 output_no[172]
port 91 nsew signal output
flabel metal2 s 67256 0 67336 80 0 FreeSans 320 0 0 0 output_no[173]
port 92 nsew signal output
flabel metal2 s 67640 0 67720 80 0 FreeSans 320 0 0 0 output_no[174]
port 93 nsew signal output
flabel metal2 s 68024 0 68104 80 0 FreeSans 320 0 0 0 output_no[175]
port 94 nsew signal output
flabel metal2 s 68408 0 68488 80 0 FreeSans 320 0 0 0 output_no[176]
port 95 nsew signal output
flabel metal2 s 68792 0 68872 80 0 FreeSans 320 0 0 0 output_no[177]
port 96 nsew signal output
flabel metal2 s 69176 0 69256 80 0 FreeSans 320 0 0 0 output_no[178]
port 97 nsew signal output
flabel metal2 s 69560 0 69640 80 0 FreeSans 320 0 0 0 output_no[179]
port 98 nsew signal output
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 output_no[17]
port 99 nsew signal output
flabel metal2 s 69944 0 70024 80 0 FreeSans 320 0 0 0 output_no[180]
port 100 nsew signal output
flabel metal2 s 70328 0 70408 80 0 FreeSans 320 0 0 0 output_no[181]
port 101 nsew signal output
flabel metal2 s 70712 0 70792 80 0 FreeSans 320 0 0 0 output_no[182]
port 102 nsew signal output
flabel metal2 s 71096 0 71176 80 0 FreeSans 320 0 0 0 output_no[183]
port 103 nsew signal output
flabel metal2 s 71480 0 71560 80 0 FreeSans 320 0 0 0 output_no[184]
port 104 nsew signal output
flabel metal2 s 71864 0 71944 80 0 FreeSans 320 0 0 0 output_no[185]
port 105 nsew signal output
flabel metal2 s 72248 0 72328 80 0 FreeSans 320 0 0 0 output_no[186]
port 106 nsew signal output
flabel metal2 s 72632 0 72712 80 0 FreeSans 320 0 0 0 output_no[187]
port 107 nsew signal output
flabel metal2 s 73016 0 73096 80 0 FreeSans 320 0 0 0 output_no[188]
port 108 nsew signal output
flabel metal2 s 73400 0 73480 80 0 FreeSans 320 0 0 0 output_no[189]
port 109 nsew signal output
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 output_no[18]
port 110 nsew signal output
flabel metal2 s 73784 0 73864 80 0 FreeSans 320 0 0 0 output_no[190]
port 111 nsew signal output
flabel metal2 s 74168 0 74248 80 0 FreeSans 320 0 0 0 output_no[191]
port 112 nsew signal output
flabel metal2 s 74552 0 74632 80 0 FreeSans 320 0 0 0 output_no[192]
port 113 nsew signal output
flabel metal2 s 74936 0 75016 80 0 FreeSans 320 0 0 0 output_no[193]
port 114 nsew signal output
flabel metal2 s 75320 0 75400 80 0 FreeSans 320 0 0 0 output_no[194]
port 115 nsew signal output
flabel metal2 s 75704 0 75784 80 0 FreeSans 320 0 0 0 output_no[195]
port 116 nsew signal output
flabel metal2 s 76088 0 76168 80 0 FreeSans 320 0 0 0 output_no[196]
port 117 nsew signal output
flabel metal2 s 76472 0 76552 80 0 FreeSans 320 0 0 0 output_no[197]
port 118 nsew signal output
flabel metal2 s 76856 0 76936 80 0 FreeSans 320 0 0 0 output_no[198]
port 119 nsew signal output
flabel metal2 s 77240 0 77320 80 0 FreeSans 320 0 0 0 output_no[199]
port 120 nsew signal output
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 output_no[19]
port 121 nsew signal output
flabel metal2 s 1208 0 1288 80 0 FreeSans 320 0 0 0 output_no[1]
port 122 nsew signal output
flabel metal2 s 77624 0 77704 80 0 FreeSans 320 0 0 0 output_no[200]
port 123 nsew signal output
flabel metal2 s 78008 0 78088 80 0 FreeSans 320 0 0 0 output_no[201]
port 124 nsew signal output
flabel metal2 s 78392 0 78472 80 0 FreeSans 320 0 0 0 output_no[202]
port 125 nsew signal output
flabel metal2 s 78776 0 78856 80 0 FreeSans 320 0 0 0 output_no[203]
port 126 nsew signal output
flabel metal2 s 79160 0 79240 80 0 FreeSans 320 0 0 0 output_no[204]
port 127 nsew signal output
flabel metal2 s 79544 0 79624 80 0 FreeSans 320 0 0 0 output_no[205]
port 128 nsew signal output
flabel metal2 s 79928 0 80008 80 0 FreeSans 320 0 0 0 output_no[206]
port 129 nsew signal output
flabel metal2 s 80312 0 80392 80 0 FreeSans 320 0 0 0 output_no[207]
port 130 nsew signal output
flabel metal2 s 80696 0 80776 80 0 FreeSans 320 0 0 0 output_no[208]
port 131 nsew signal output
flabel metal2 s 81080 0 81160 80 0 FreeSans 320 0 0 0 output_no[209]
port 132 nsew signal output
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 output_no[20]
port 133 nsew signal output
flabel metal2 s 81464 0 81544 80 0 FreeSans 320 0 0 0 output_no[210]
port 134 nsew signal output
flabel metal2 s 81848 0 81928 80 0 FreeSans 320 0 0 0 output_no[211]
port 135 nsew signal output
flabel metal2 s 82232 0 82312 80 0 FreeSans 320 0 0 0 output_no[212]
port 136 nsew signal output
flabel metal2 s 82616 0 82696 80 0 FreeSans 320 0 0 0 output_no[213]
port 137 nsew signal output
flabel metal2 s 83000 0 83080 80 0 FreeSans 320 0 0 0 output_no[214]
port 138 nsew signal output
flabel metal2 s 83384 0 83464 80 0 FreeSans 320 0 0 0 output_no[215]
port 139 nsew signal output
flabel metal2 s 83768 0 83848 80 0 FreeSans 320 0 0 0 output_no[216]
port 140 nsew signal output
flabel metal2 s 84152 0 84232 80 0 FreeSans 320 0 0 0 output_no[217]
port 141 nsew signal output
flabel metal2 s 84536 0 84616 80 0 FreeSans 320 0 0 0 output_no[218]
port 142 nsew signal output
flabel metal2 s 84920 0 85000 80 0 FreeSans 320 0 0 0 output_no[219]
port 143 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 output_no[21]
port 144 nsew signal output
flabel metal2 s 85304 0 85384 80 0 FreeSans 320 0 0 0 output_no[220]
port 145 nsew signal output
flabel metal2 s 85688 0 85768 80 0 FreeSans 320 0 0 0 output_no[221]
port 146 nsew signal output
flabel metal2 s 86072 0 86152 80 0 FreeSans 320 0 0 0 output_no[222]
port 147 nsew signal output
flabel metal2 s 86456 0 86536 80 0 FreeSans 320 0 0 0 output_no[223]
port 148 nsew signal output
flabel metal2 s 86840 0 86920 80 0 FreeSans 320 0 0 0 output_no[224]
port 149 nsew signal output
flabel metal2 s 87224 0 87304 80 0 FreeSans 320 0 0 0 output_no[225]
port 150 nsew signal output
flabel metal2 s 87608 0 87688 80 0 FreeSans 320 0 0 0 output_no[226]
port 151 nsew signal output
flabel metal2 s 87992 0 88072 80 0 FreeSans 320 0 0 0 output_no[227]
port 152 nsew signal output
flabel metal2 s 88376 0 88456 80 0 FreeSans 320 0 0 0 output_no[228]
port 153 nsew signal output
flabel metal2 s 88760 0 88840 80 0 FreeSans 320 0 0 0 output_no[229]
port 154 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 output_no[22]
port 155 nsew signal output
flabel metal2 s 89144 0 89224 80 0 FreeSans 320 0 0 0 output_no[230]
port 156 nsew signal output
flabel metal2 s 89528 0 89608 80 0 FreeSans 320 0 0 0 output_no[231]
port 157 nsew signal output
flabel metal2 s 89912 0 89992 80 0 FreeSans 320 0 0 0 output_no[232]
port 158 nsew signal output
flabel metal2 s 90296 0 90376 80 0 FreeSans 320 0 0 0 output_no[233]
port 159 nsew signal output
flabel metal2 s 90680 0 90760 80 0 FreeSans 320 0 0 0 output_no[234]
port 160 nsew signal output
flabel metal2 s 91064 0 91144 80 0 FreeSans 320 0 0 0 output_no[235]
port 161 nsew signal output
flabel metal2 s 91448 0 91528 80 0 FreeSans 320 0 0 0 output_no[236]
port 162 nsew signal output
flabel metal2 s 91832 0 91912 80 0 FreeSans 320 0 0 0 output_no[237]
port 163 nsew signal output
flabel metal2 s 92216 0 92296 80 0 FreeSans 320 0 0 0 output_no[238]
port 164 nsew signal output
flabel metal2 s 92600 0 92680 80 0 FreeSans 320 0 0 0 output_no[239]
port 165 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 output_no[23]
port 166 nsew signal output
flabel metal2 s 92984 0 93064 80 0 FreeSans 320 0 0 0 output_no[240]
port 167 nsew signal output
flabel metal2 s 93368 0 93448 80 0 FreeSans 320 0 0 0 output_no[241]
port 168 nsew signal output
flabel metal2 s 93752 0 93832 80 0 FreeSans 320 0 0 0 output_no[242]
port 169 nsew signal output
flabel metal2 s 94136 0 94216 80 0 FreeSans 320 0 0 0 output_no[243]
port 170 nsew signal output
flabel metal2 s 94520 0 94600 80 0 FreeSans 320 0 0 0 output_no[244]
port 171 nsew signal output
flabel metal2 s 94904 0 94984 80 0 FreeSans 320 0 0 0 output_no[245]
port 172 nsew signal output
flabel metal2 s 95288 0 95368 80 0 FreeSans 320 0 0 0 output_no[246]
port 173 nsew signal output
flabel metal2 s 95672 0 95752 80 0 FreeSans 320 0 0 0 output_no[247]
port 174 nsew signal output
flabel metal2 s 96056 0 96136 80 0 FreeSans 320 0 0 0 output_no[248]
port 175 nsew signal output
flabel metal2 s 96440 0 96520 80 0 FreeSans 320 0 0 0 output_no[249]
port 176 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 output_no[24]
port 177 nsew signal output
flabel metal2 s 96824 0 96904 80 0 FreeSans 320 0 0 0 output_no[250]
port 178 nsew signal output
flabel metal2 s 97208 0 97288 80 0 FreeSans 320 0 0 0 output_no[251]
port 179 nsew signal output
flabel metal2 s 97592 0 97672 80 0 FreeSans 320 0 0 0 output_no[252]
port 180 nsew signal output
flabel metal2 s 97976 0 98056 80 0 FreeSans 320 0 0 0 output_no[253]
port 181 nsew signal output
flabel metal2 s 98360 0 98440 80 0 FreeSans 320 0 0 0 output_no[254]
port 182 nsew signal output
flabel metal2 s 98744 0 98824 80 0 FreeSans 320 0 0 0 output_no[255]
port 183 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 output_no[25]
port 184 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 output_no[26]
port 185 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 output_no[27]
port 186 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 output_no[28]
port 187 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 output_no[29]
port 188 nsew signal output
flabel metal2 s 1592 0 1672 80 0 FreeSans 320 0 0 0 output_no[2]
port 189 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 output_no[30]
port 190 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 output_no[31]
port 191 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 output_no[32]
port 192 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 output_no[33]
port 193 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 output_no[34]
port 194 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 output_no[35]
port 195 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 output_no[36]
port 196 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 output_no[37]
port 197 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 output_no[38]
port 198 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 output_no[39]
port 199 nsew signal output
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 output_no[3]
port 200 nsew signal output
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 output_no[40]
port 201 nsew signal output
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 output_no[41]
port 202 nsew signal output
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 output_no[42]
port 203 nsew signal output
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 output_no[43]
port 204 nsew signal output
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 output_no[44]
port 205 nsew signal output
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 output_no[45]
port 206 nsew signal output
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 output_no[46]
port 207 nsew signal output
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 output_no[47]
port 208 nsew signal output
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 output_no[48]
port 209 nsew signal output
flabel metal2 s 19640 0 19720 80 0 FreeSans 320 0 0 0 output_no[49]
port 210 nsew signal output
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 output_no[4]
port 211 nsew signal output
flabel metal2 s 20024 0 20104 80 0 FreeSans 320 0 0 0 output_no[50]
port 212 nsew signal output
flabel metal2 s 20408 0 20488 80 0 FreeSans 320 0 0 0 output_no[51]
port 213 nsew signal output
flabel metal2 s 20792 0 20872 80 0 FreeSans 320 0 0 0 output_no[52]
port 214 nsew signal output
flabel metal2 s 21176 0 21256 80 0 FreeSans 320 0 0 0 output_no[53]
port 215 nsew signal output
flabel metal2 s 21560 0 21640 80 0 FreeSans 320 0 0 0 output_no[54]
port 216 nsew signal output
flabel metal2 s 21944 0 22024 80 0 FreeSans 320 0 0 0 output_no[55]
port 217 nsew signal output
flabel metal2 s 22328 0 22408 80 0 FreeSans 320 0 0 0 output_no[56]
port 218 nsew signal output
flabel metal2 s 22712 0 22792 80 0 FreeSans 320 0 0 0 output_no[57]
port 219 nsew signal output
flabel metal2 s 23096 0 23176 80 0 FreeSans 320 0 0 0 output_no[58]
port 220 nsew signal output
flabel metal2 s 23480 0 23560 80 0 FreeSans 320 0 0 0 output_no[59]
port 221 nsew signal output
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 output_no[5]
port 222 nsew signal output
flabel metal2 s 23864 0 23944 80 0 FreeSans 320 0 0 0 output_no[60]
port 223 nsew signal output
flabel metal2 s 24248 0 24328 80 0 FreeSans 320 0 0 0 output_no[61]
port 224 nsew signal output
flabel metal2 s 24632 0 24712 80 0 FreeSans 320 0 0 0 output_no[62]
port 225 nsew signal output
flabel metal2 s 25016 0 25096 80 0 FreeSans 320 0 0 0 output_no[63]
port 226 nsew signal output
flabel metal2 s 25400 0 25480 80 0 FreeSans 320 0 0 0 output_no[64]
port 227 nsew signal output
flabel metal2 s 25784 0 25864 80 0 FreeSans 320 0 0 0 output_no[65]
port 228 nsew signal output
flabel metal2 s 26168 0 26248 80 0 FreeSans 320 0 0 0 output_no[66]
port 229 nsew signal output
flabel metal2 s 26552 0 26632 80 0 FreeSans 320 0 0 0 output_no[67]
port 230 nsew signal output
flabel metal2 s 26936 0 27016 80 0 FreeSans 320 0 0 0 output_no[68]
port 231 nsew signal output
flabel metal2 s 27320 0 27400 80 0 FreeSans 320 0 0 0 output_no[69]
port 232 nsew signal output
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 output_no[6]
port 233 nsew signal output
flabel metal2 s 27704 0 27784 80 0 FreeSans 320 0 0 0 output_no[70]
port 234 nsew signal output
flabel metal2 s 28088 0 28168 80 0 FreeSans 320 0 0 0 output_no[71]
port 235 nsew signal output
flabel metal2 s 28472 0 28552 80 0 FreeSans 320 0 0 0 output_no[72]
port 236 nsew signal output
flabel metal2 s 28856 0 28936 80 0 FreeSans 320 0 0 0 output_no[73]
port 237 nsew signal output
flabel metal2 s 29240 0 29320 80 0 FreeSans 320 0 0 0 output_no[74]
port 238 nsew signal output
flabel metal2 s 29624 0 29704 80 0 FreeSans 320 0 0 0 output_no[75]
port 239 nsew signal output
flabel metal2 s 30008 0 30088 80 0 FreeSans 320 0 0 0 output_no[76]
port 240 nsew signal output
flabel metal2 s 30392 0 30472 80 0 FreeSans 320 0 0 0 output_no[77]
port 241 nsew signal output
flabel metal2 s 30776 0 30856 80 0 FreeSans 320 0 0 0 output_no[78]
port 242 nsew signal output
flabel metal2 s 31160 0 31240 80 0 FreeSans 320 0 0 0 output_no[79]
port 243 nsew signal output
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 output_no[7]
port 244 nsew signal output
flabel metal2 s 31544 0 31624 80 0 FreeSans 320 0 0 0 output_no[80]
port 245 nsew signal output
flabel metal2 s 31928 0 32008 80 0 FreeSans 320 0 0 0 output_no[81]
port 246 nsew signal output
flabel metal2 s 32312 0 32392 80 0 FreeSans 320 0 0 0 output_no[82]
port 247 nsew signal output
flabel metal2 s 32696 0 32776 80 0 FreeSans 320 0 0 0 output_no[83]
port 248 nsew signal output
flabel metal2 s 33080 0 33160 80 0 FreeSans 320 0 0 0 output_no[84]
port 249 nsew signal output
flabel metal2 s 33464 0 33544 80 0 FreeSans 320 0 0 0 output_no[85]
port 250 nsew signal output
flabel metal2 s 33848 0 33928 80 0 FreeSans 320 0 0 0 output_no[86]
port 251 nsew signal output
flabel metal2 s 34232 0 34312 80 0 FreeSans 320 0 0 0 output_no[87]
port 252 nsew signal output
flabel metal2 s 34616 0 34696 80 0 FreeSans 320 0 0 0 output_no[88]
port 253 nsew signal output
flabel metal2 s 35000 0 35080 80 0 FreeSans 320 0 0 0 output_no[89]
port 254 nsew signal output
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 output_no[8]
port 255 nsew signal output
flabel metal2 s 35384 0 35464 80 0 FreeSans 320 0 0 0 output_no[90]
port 256 nsew signal output
flabel metal2 s 35768 0 35848 80 0 FreeSans 320 0 0 0 output_no[91]
port 257 nsew signal output
flabel metal2 s 36152 0 36232 80 0 FreeSans 320 0 0 0 output_no[92]
port 258 nsew signal output
flabel metal2 s 36536 0 36616 80 0 FreeSans 320 0 0 0 output_no[93]
port 259 nsew signal output
flabel metal2 s 36920 0 37000 80 0 FreeSans 320 0 0 0 output_no[94]
port 260 nsew signal output
flabel metal2 s 37304 0 37384 80 0 FreeSans 320 0 0 0 output_no[95]
port 261 nsew signal output
flabel metal2 s 37688 0 37768 80 0 FreeSans 320 0 0 0 output_no[96]
port 262 nsew signal output
flabel metal2 s 38072 0 38152 80 0 FreeSans 320 0 0 0 output_no[97]
port 263 nsew signal output
flabel metal2 s 38456 0 38536 80 0 FreeSans 320 0 0 0 output_no[98]
port 264 nsew signal output
flabel metal2 s 38840 0 38920 80 0 FreeSans 320 0 0 0 output_no[99]
port 265 nsew signal output
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 output_no[9]
port 266 nsew signal output
flabel metal2 s 1016 0 1096 80 0 FreeSans 320 0 0 0 output_o[0]
port 267 nsew signal output
flabel metal2 s 39416 0 39496 80 0 FreeSans 320 0 0 0 output_o[100]
port 268 nsew signal output
flabel metal2 s 39800 0 39880 80 0 FreeSans 320 0 0 0 output_o[101]
port 269 nsew signal output
flabel metal2 s 40184 0 40264 80 0 FreeSans 320 0 0 0 output_o[102]
port 270 nsew signal output
flabel metal2 s 40568 0 40648 80 0 FreeSans 320 0 0 0 output_o[103]
port 271 nsew signal output
flabel metal2 s 40952 0 41032 80 0 FreeSans 320 0 0 0 output_o[104]
port 272 nsew signal output
flabel metal2 s 41336 0 41416 80 0 FreeSans 320 0 0 0 output_o[105]
port 273 nsew signal output
flabel metal2 s 41720 0 41800 80 0 FreeSans 320 0 0 0 output_o[106]
port 274 nsew signal output
flabel metal2 s 42104 0 42184 80 0 FreeSans 320 0 0 0 output_o[107]
port 275 nsew signal output
flabel metal2 s 42488 0 42568 80 0 FreeSans 320 0 0 0 output_o[108]
port 276 nsew signal output
flabel metal2 s 42872 0 42952 80 0 FreeSans 320 0 0 0 output_o[109]
port 277 nsew signal output
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 output_o[10]
port 278 nsew signal output
flabel metal2 s 43256 0 43336 80 0 FreeSans 320 0 0 0 output_o[110]
port 279 nsew signal output
flabel metal2 s 43640 0 43720 80 0 FreeSans 320 0 0 0 output_o[111]
port 280 nsew signal output
flabel metal2 s 44024 0 44104 80 0 FreeSans 320 0 0 0 output_o[112]
port 281 nsew signal output
flabel metal2 s 44408 0 44488 80 0 FreeSans 320 0 0 0 output_o[113]
port 282 nsew signal output
flabel metal2 s 44792 0 44872 80 0 FreeSans 320 0 0 0 output_o[114]
port 283 nsew signal output
flabel metal2 s 45176 0 45256 80 0 FreeSans 320 0 0 0 output_o[115]
port 284 nsew signal output
flabel metal2 s 45560 0 45640 80 0 FreeSans 320 0 0 0 output_o[116]
port 285 nsew signal output
flabel metal2 s 45944 0 46024 80 0 FreeSans 320 0 0 0 output_o[117]
port 286 nsew signal output
flabel metal2 s 46328 0 46408 80 0 FreeSans 320 0 0 0 output_o[118]
port 287 nsew signal output
flabel metal2 s 46712 0 46792 80 0 FreeSans 320 0 0 0 output_o[119]
port 288 nsew signal output
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 output_o[11]
port 289 nsew signal output
flabel metal2 s 47096 0 47176 80 0 FreeSans 320 0 0 0 output_o[120]
port 290 nsew signal output
flabel metal2 s 47480 0 47560 80 0 FreeSans 320 0 0 0 output_o[121]
port 291 nsew signal output
flabel metal2 s 47864 0 47944 80 0 FreeSans 320 0 0 0 output_o[122]
port 292 nsew signal output
flabel metal2 s 48248 0 48328 80 0 FreeSans 320 0 0 0 output_o[123]
port 293 nsew signal output
flabel metal2 s 48632 0 48712 80 0 FreeSans 320 0 0 0 output_o[124]
port 294 nsew signal output
flabel metal2 s 49016 0 49096 80 0 FreeSans 320 0 0 0 output_o[125]
port 295 nsew signal output
flabel metal2 s 49400 0 49480 80 0 FreeSans 320 0 0 0 output_o[126]
port 296 nsew signal output
flabel metal2 s 49784 0 49864 80 0 FreeSans 320 0 0 0 output_o[127]
port 297 nsew signal output
flabel metal2 s 50168 0 50248 80 0 FreeSans 320 0 0 0 output_o[128]
port 298 nsew signal output
flabel metal2 s 50552 0 50632 80 0 FreeSans 320 0 0 0 output_o[129]
port 299 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 output_o[12]
port 300 nsew signal output
flabel metal2 s 50936 0 51016 80 0 FreeSans 320 0 0 0 output_o[130]
port 301 nsew signal output
flabel metal2 s 51320 0 51400 80 0 FreeSans 320 0 0 0 output_o[131]
port 302 nsew signal output
flabel metal2 s 51704 0 51784 80 0 FreeSans 320 0 0 0 output_o[132]
port 303 nsew signal output
flabel metal2 s 52088 0 52168 80 0 FreeSans 320 0 0 0 output_o[133]
port 304 nsew signal output
flabel metal2 s 52472 0 52552 80 0 FreeSans 320 0 0 0 output_o[134]
port 305 nsew signal output
flabel metal2 s 52856 0 52936 80 0 FreeSans 320 0 0 0 output_o[135]
port 306 nsew signal output
flabel metal2 s 53240 0 53320 80 0 FreeSans 320 0 0 0 output_o[136]
port 307 nsew signal output
flabel metal2 s 53624 0 53704 80 0 FreeSans 320 0 0 0 output_o[137]
port 308 nsew signal output
flabel metal2 s 54008 0 54088 80 0 FreeSans 320 0 0 0 output_o[138]
port 309 nsew signal output
flabel metal2 s 54392 0 54472 80 0 FreeSans 320 0 0 0 output_o[139]
port 310 nsew signal output
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 output_o[13]
port 311 nsew signal output
flabel metal2 s 54776 0 54856 80 0 FreeSans 320 0 0 0 output_o[140]
port 312 nsew signal output
flabel metal2 s 55160 0 55240 80 0 FreeSans 320 0 0 0 output_o[141]
port 313 nsew signal output
flabel metal2 s 55544 0 55624 80 0 FreeSans 320 0 0 0 output_o[142]
port 314 nsew signal output
flabel metal2 s 55928 0 56008 80 0 FreeSans 320 0 0 0 output_o[143]
port 315 nsew signal output
flabel metal2 s 56312 0 56392 80 0 FreeSans 320 0 0 0 output_o[144]
port 316 nsew signal output
flabel metal2 s 56696 0 56776 80 0 FreeSans 320 0 0 0 output_o[145]
port 317 nsew signal output
flabel metal2 s 57080 0 57160 80 0 FreeSans 320 0 0 0 output_o[146]
port 318 nsew signal output
flabel metal2 s 57464 0 57544 80 0 FreeSans 320 0 0 0 output_o[147]
port 319 nsew signal output
flabel metal2 s 57848 0 57928 80 0 FreeSans 320 0 0 0 output_o[148]
port 320 nsew signal output
flabel metal2 s 58232 0 58312 80 0 FreeSans 320 0 0 0 output_o[149]
port 321 nsew signal output
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 output_o[14]
port 322 nsew signal output
flabel metal2 s 58616 0 58696 80 0 FreeSans 320 0 0 0 output_o[150]
port 323 nsew signal output
flabel metal2 s 59000 0 59080 80 0 FreeSans 320 0 0 0 output_o[151]
port 324 nsew signal output
flabel metal2 s 59384 0 59464 80 0 FreeSans 320 0 0 0 output_o[152]
port 325 nsew signal output
flabel metal2 s 59768 0 59848 80 0 FreeSans 320 0 0 0 output_o[153]
port 326 nsew signal output
flabel metal2 s 60152 0 60232 80 0 FreeSans 320 0 0 0 output_o[154]
port 327 nsew signal output
flabel metal2 s 60536 0 60616 80 0 FreeSans 320 0 0 0 output_o[155]
port 328 nsew signal output
flabel metal2 s 60920 0 61000 80 0 FreeSans 320 0 0 0 output_o[156]
port 329 nsew signal output
flabel metal2 s 61304 0 61384 80 0 FreeSans 320 0 0 0 output_o[157]
port 330 nsew signal output
flabel metal2 s 61688 0 61768 80 0 FreeSans 320 0 0 0 output_o[158]
port 331 nsew signal output
flabel metal2 s 62072 0 62152 80 0 FreeSans 320 0 0 0 output_o[159]
port 332 nsew signal output
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 output_o[15]
port 333 nsew signal output
flabel metal2 s 62456 0 62536 80 0 FreeSans 320 0 0 0 output_o[160]
port 334 nsew signal output
flabel metal2 s 62840 0 62920 80 0 FreeSans 320 0 0 0 output_o[161]
port 335 nsew signal output
flabel metal2 s 63224 0 63304 80 0 FreeSans 320 0 0 0 output_o[162]
port 336 nsew signal output
flabel metal2 s 63608 0 63688 80 0 FreeSans 320 0 0 0 output_o[163]
port 337 nsew signal output
flabel metal2 s 63992 0 64072 80 0 FreeSans 320 0 0 0 output_o[164]
port 338 nsew signal output
flabel metal2 s 64376 0 64456 80 0 FreeSans 320 0 0 0 output_o[165]
port 339 nsew signal output
flabel metal2 s 64760 0 64840 80 0 FreeSans 320 0 0 0 output_o[166]
port 340 nsew signal output
flabel metal2 s 65144 0 65224 80 0 FreeSans 320 0 0 0 output_o[167]
port 341 nsew signal output
flabel metal2 s 65528 0 65608 80 0 FreeSans 320 0 0 0 output_o[168]
port 342 nsew signal output
flabel metal2 s 65912 0 65992 80 0 FreeSans 320 0 0 0 output_o[169]
port 343 nsew signal output
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 output_o[16]
port 344 nsew signal output
flabel metal2 s 66296 0 66376 80 0 FreeSans 320 0 0 0 output_o[170]
port 345 nsew signal output
flabel metal2 s 66680 0 66760 80 0 FreeSans 320 0 0 0 output_o[171]
port 346 nsew signal output
flabel metal2 s 67064 0 67144 80 0 FreeSans 320 0 0 0 output_o[172]
port 347 nsew signal output
flabel metal2 s 67448 0 67528 80 0 FreeSans 320 0 0 0 output_o[173]
port 348 nsew signal output
flabel metal2 s 67832 0 67912 80 0 FreeSans 320 0 0 0 output_o[174]
port 349 nsew signal output
flabel metal2 s 68216 0 68296 80 0 FreeSans 320 0 0 0 output_o[175]
port 350 nsew signal output
flabel metal2 s 68600 0 68680 80 0 FreeSans 320 0 0 0 output_o[176]
port 351 nsew signal output
flabel metal2 s 68984 0 69064 80 0 FreeSans 320 0 0 0 output_o[177]
port 352 nsew signal output
flabel metal2 s 69368 0 69448 80 0 FreeSans 320 0 0 0 output_o[178]
port 353 nsew signal output
flabel metal2 s 69752 0 69832 80 0 FreeSans 320 0 0 0 output_o[179]
port 354 nsew signal output
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 output_o[17]
port 355 nsew signal output
flabel metal2 s 70136 0 70216 80 0 FreeSans 320 0 0 0 output_o[180]
port 356 nsew signal output
flabel metal2 s 70520 0 70600 80 0 FreeSans 320 0 0 0 output_o[181]
port 357 nsew signal output
flabel metal2 s 70904 0 70984 80 0 FreeSans 320 0 0 0 output_o[182]
port 358 nsew signal output
flabel metal2 s 71288 0 71368 80 0 FreeSans 320 0 0 0 output_o[183]
port 359 nsew signal output
flabel metal2 s 71672 0 71752 80 0 FreeSans 320 0 0 0 output_o[184]
port 360 nsew signal output
flabel metal2 s 72056 0 72136 80 0 FreeSans 320 0 0 0 output_o[185]
port 361 nsew signal output
flabel metal2 s 72440 0 72520 80 0 FreeSans 320 0 0 0 output_o[186]
port 362 nsew signal output
flabel metal2 s 72824 0 72904 80 0 FreeSans 320 0 0 0 output_o[187]
port 363 nsew signal output
flabel metal2 s 73208 0 73288 80 0 FreeSans 320 0 0 0 output_o[188]
port 364 nsew signal output
flabel metal2 s 73592 0 73672 80 0 FreeSans 320 0 0 0 output_o[189]
port 365 nsew signal output
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 output_o[18]
port 366 nsew signal output
flabel metal2 s 73976 0 74056 80 0 FreeSans 320 0 0 0 output_o[190]
port 367 nsew signal output
flabel metal2 s 74360 0 74440 80 0 FreeSans 320 0 0 0 output_o[191]
port 368 nsew signal output
flabel metal2 s 74744 0 74824 80 0 FreeSans 320 0 0 0 output_o[192]
port 369 nsew signal output
flabel metal2 s 75128 0 75208 80 0 FreeSans 320 0 0 0 output_o[193]
port 370 nsew signal output
flabel metal2 s 75512 0 75592 80 0 FreeSans 320 0 0 0 output_o[194]
port 371 nsew signal output
flabel metal2 s 75896 0 75976 80 0 FreeSans 320 0 0 0 output_o[195]
port 372 nsew signal output
flabel metal2 s 76280 0 76360 80 0 FreeSans 320 0 0 0 output_o[196]
port 373 nsew signal output
flabel metal2 s 76664 0 76744 80 0 FreeSans 320 0 0 0 output_o[197]
port 374 nsew signal output
flabel metal2 s 77048 0 77128 80 0 FreeSans 320 0 0 0 output_o[198]
port 375 nsew signal output
flabel metal2 s 77432 0 77512 80 0 FreeSans 320 0 0 0 output_o[199]
port 376 nsew signal output
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 output_o[19]
port 377 nsew signal output
flabel metal2 s 1400 0 1480 80 0 FreeSans 320 0 0 0 output_o[1]
port 378 nsew signal output
flabel metal2 s 77816 0 77896 80 0 FreeSans 320 0 0 0 output_o[200]
port 379 nsew signal output
flabel metal2 s 78200 0 78280 80 0 FreeSans 320 0 0 0 output_o[201]
port 380 nsew signal output
flabel metal2 s 78584 0 78664 80 0 FreeSans 320 0 0 0 output_o[202]
port 381 nsew signal output
flabel metal2 s 78968 0 79048 80 0 FreeSans 320 0 0 0 output_o[203]
port 382 nsew signal output
flabel metal2 s 79352 0 79432 80 0 FreeSans 320 0 0 0 output_o[204]
port 383 nsew signal output
flabel metal2 s 79736 0 79816 80 0 FreeSans 320 0 0 0 output_o[205]
port 384 nsew signal output
flabel metal2 s 80120 0 80200 80 0 FreeSans 320 0 0 0 output_o[206]
port 385 nsew signal output
flabel metal2 s 80504 0 80584 80 0 FreeSans 320 0 0 0 output_o[207]
port 386 nsew signal output
flabel metal2 s 80888 0 80968 80 0 FreeSans 320 0 0 0 output_o[208]
port 387 nsew signal output
flabel metal2 s 81272 0 81352 80 0 FreeSans 320 0 0 0 output_o[209]
port 388 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 output_o[20]
port 389 nsew signal output
flabel metal2 s 81656 0 81736 80 0 FreeSans 320 0 0 0 output_o[210]
port 390 nsew signal output
flabel metal2 s 82040 0 82120 80 0 FreeSans 320 0 0 0 output_o[211]
port 391 nsew signal output
flabel metal2 s 82424 0 82504 80 0 FreeSans 320 0 0 0 output_o[212]
port 392 nsew signal output
flabel metal2 s 82808 0 82888 80 0 FreeSans 320 0 0 0 output_o[213]
port 393 nsew signal output
flabel metal2 s 83192 0 83272 80 0 FreeSans 320 0 0 0 output_o[214]
port 394 nsew signal output
flabel metal2 s 83576 0 83656 80 0 FreeSans 320 0 0 0 output_o[215]
port 395 nsew signal output
flabel metal2 s 83960 0 84040 80 0 FreeSans 320 0 0 0 output_o[216]
port 396 nsew signal output
flabel metal2 s 84344 0 84424 80 0 FreeSans 320 0 0 0 output_o[217]
port 397 nsew signal output
flabel metal2 s 84728 0 84808 80 0 FreeSans 320 0 0 0 output_o[218]
port 398 nsew signal output
flabel metal2 s 85112 0 85192 80 0 FreeSans 320 0 0 0 output_o[219]
port 399 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 output_o[21]
port 400 nsew signal output
flabel metal2 s 85496 0 85576 80 0 FreeSans 320 0 0 0 output_o[220]
port 401 nsew signal output
flabel metal2 s 85880 0 85960 80 0 FreeSans 320 0 0 0 output_o[221]
port 402 nsew signal output
flabel metal2 s 86264 0 86344 80 0 FreeSans 320 0 0 0 output_o[222]
port 403 nsew signal output
flabel metal2 s 86648 0 86728 80 0 FreeSans 320 0 0 0 output_o[223]
port 404 nsew signal output
flabel metal2 s 87032 0 87112 80 0 FreeSans 320 0 0 0 output_o[224]
port 405 nsew signal output
flabel metal2 s 87416 0 87496 80 0 FreeSans 320 0 0 0 output_o[225]
port 406 nsew signal output
flabel metal2 s 87800 0 87880 80 0 FreeSans 320 0 0 0 output_o[226]
port 407 nsew signal output
flabel metal2 s 88184 0 88264 80 0 FreeSans 320 0 0 0 output_o[227]
port 408 nsew signal output
flabel metal2 s 88568 0 88648 80 0 FreeSans 320 0 0 0 output_o[228]
port 409 nsew signal output
flabel metal2 s 88952 0 89032 80 0 FreeSans 320 0 0 0 output_o[229]
port 410 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 output_o[22]
port 411 nsew signal output
flabel metal2 s 89336 0 89416 80 0 FreeSans 320 0 0 0 output_o[230]
port 412 nsew signal output
flabel metal2 s 89720 0 89800 80 0 FreeSans 320 0 0 0 output_o[231]
port 413 nsew signal output
flabel metal2 s 90104 0 90184 80 0 FreeSans 320 0 0 0 output_o[232]
port 414 nsew signal output
flabel metal2 s 90488 0 90568 80 0 FreeSans 320 0 0 0 output_o[233]
port 415 nsew signal output
flabel metal2 s 90872 0 90952 80 0 FreeSans 320 0 0 0 output_o[234]
port 416 nsew signal output
flabel metal2 s 91256 0 91336 80 0 FreeSans 320 0 0 0 output_o[235]
port 417 nsew signal output
flabel metal2 s 91640 0 91720 80 0 FreeSans 320 0 0 0 output_o[236]
port 418 nsew signal output
flabel metal2 s 92024 0 92104 80 0 FreeSans 320 0 0 0 output_o[237]
port 419 nsew signal output
flabel metal2 s 92408 0 92488 80 0 FreeSans 320 0 0 0 output_o[238]
port 420 nsew signal output
flabel metal2 s 92792 0 92872 80 0 FreeSans 320 0 0 0 output_o[239]
port 421 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 output_o[23]
port 422 nsew signal output
flabel metal2 s 93176 0 93256 80 0 FreeSans 320 0 0 0 output_o[240]
port 423 nsew signal output
flabel metal2 s 93560 0 93640 80 0 FreeSans 320 0 0 0 output_o[241]
port 424 nsew signal output
flabel metal2 s 93944 0 94024 80 0 FreeSans 320 0 0 0 output_o[242]
port 425 nsew signal output
flabel metal2 s 94328 0 94408 80 0 FreeSans 320 0 0 0 output_o[243]
port 426 nsew signal output
flabel metal2 s 94712 0 94792 80 0 FreeSans 320 0 0 0 output_o[244]
port 427 nsew signal output
flabel metal2 s 95096 0 95176 80 0 FreeSans 320 0 0 0 output_o[245]
port 428 nsew signal output
flabel metal2 s 95480 0 95560 80 0 FreeSans 320 0 0 0 output_o[246]
port 429 nsew signal output
flabel metal2 s 95864 0 95944 80 0 FreeSans 320 0 0 0 output_o[247]
port 430 nsew signal output
flabel metal2 s 96248 0 96328 80 0 FreeSans 320 0 0 0 output_o[248]
port 431 nsew signal output
flabel metal2 s 96632 0 96712 80 0 FreeSans 320 0 0 0 output_o[249]
port 432 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 output_o[24]
port 433 nsew signal output
flabel metal2 s 97016 0 97096 80 0 FreeSans 320 0 0 0 output_o[250]
port 434 nsew signal output
flabel metal2 s 97400 0 97480 80 0 FreeSans 320 0 0 0 output_o[251]
port 435 nsew signal output
flabel metal2 s 97784 0 97864 80 0 FreeSans 320 0 0 0 output_o[252]
port 436 nsew signal output
flabel metal2 s 98168 0 98248 80 0 FreeSans 320 0 0 0 output_o[253]
port 437 nsew signal output
flabel metal2 s 98552 0 98632 80 0 FreeSans 320 0 0 0 output_o[254]
port 438 nsew signal output
flabel metal2 s 98936 0 99016 80 0 FreeSans 320 0 0 0 output_o[255]
port 439 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 output_o[25]
port 440 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 output_o[26]
port 441 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 output_o[27]
port 442 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 output_o[28]
port 443 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 output_o[29]
port 444 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 output_o[2]
port 445 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 output_o[30]
port 446 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 output_o[31]
port 447 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 output_o[32]
port 448 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 output_o[33]
port 449 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 output_o[34]
port 450 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 output_o[35]
port 451 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 output_o[36]
port 452 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 output_o[37]
port 453 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 output_o[38]
port 454 nsew signal output
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 output_o[39]
port 455 nsew signal output
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 output_o[3]
port 456 nsew signal output
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 output_o[40]
port 457 nsew signal output
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 output_o[41]
port 458 nsew signal output
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 output_o[42]
port 459 nsew signal output
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 output_o[43]
port 460 nsew signal output
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 output_o[44]
port 461 nsew signal output
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 output_o[45]
port 462 nsew signal output
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 output_o[46]
port 463 nsew signal output
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 output_o[47]
port 464 nsew signal output
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 output_o[48]
port 465 nsew signal output
flabel metal2 s 19832 0 19912 80 0 FreeSans 320 0 0 0 output_o[49]
port 466 nsew signal output
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 output_o[4]
port 467 nsew signal output
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 output_o[50]
port 468 nsew signal output
flabel metal2 s 20600 0 20680 80 0 FreeSans 320 0 0 0 output_o[51]
port 469 nsew signal output
flabel metal2 s 20984 0 21064 80 0 FreeSans 320 0 0 0 output_o[52]
port 470 nsew signal output
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 output_o[53]
port 471 nsew signal output
flabel metal2 s 21752 0 21832 80 0 FreeSans 320 0 0 0 output_o[54]
port 472 nsew signal output
flabel metal2 s 22136 0 22216 80 0 FreeSans 320 0 0 0 output_o[55]
port 473 nsew signal output
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 output_o[56]
port 474 nsew signal output
flabel metal2 s 22904 0 22984 80 0 FreeSans 320 0 0 0 output_o[57]
port 475 nsew signal output
flabel metal2 s 23288 0 23368 80 0 FreeSans 320 0 0 0 output_o[58]
port 476 nsew signal output
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 output_o[59]
port 477 nsew signal output
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 output_o[5]
port 478 nsew signal output
flabel metal2 s 24056 0 24136 80 0 FreeSans 320 0 0 0 output_o[60]
port 479 nsew signal output
flabel metal2 s 24440 0 24520 80 0 FreeSans 320 0 0 0 output_o[61]
port 480 nsew signal output
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 output_o[62]
port 481 nsew signal output
flabel metal2 s 25208 0 25288 80 0 FreeSans 320 0 0 0 output_o[63]
port 482 nsew signal output
flabel metal2 s 25592 0 25672 80 0 FreeSans 320 0 0 0 output_o[64]
port 483 nsew signal output
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 output_o[65]
port 484 nsew signal output
flabel metal2 s 26360 0 26440 80 0 FreeSans 320 0 0 0 output_o[66]
port 485 nsew signal output
flabel metal2 s 26744 0 26824 80 0 FreeSans 320 0 0 0 output_o[67]
port 486 nsew signal output
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 output_o[68]
port 487 nsew signal output
flabel metal2 s 27512 0 27592 80 0 FreeSans 320 0 0 0 output_o[69]
port 488 nsew signal output
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 output_o[6]
port 489 nsew signal output
flabel metal2 s 27896 0 27976 80 0 FreeSans 320 0 0 0 output_o[70]
port 490 nsew signal output
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 output_o[71]
port 491 nsew signal output
flabel metal2 s 28664 0 28744 80 0 FreeSans 320 0 0 0 output_o[72]
port 492 nsew signal output
flabel metal2 s 29048 0 29128 80 0 FreeSans 320 0 0 0 output_o[73]
port 493 nsew signal output
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 output_o[74]
port 494 nsew signal output
flabel metal2 s 29816 0 29896 80 0 FreeSans 320 0 0 0 output_o[75]
port 495 nsew signal output
flabel metal2 s 30200 0 30280 80 0 FreeSans 320 0 0 0 output_o[76]
port 496 nsew signal output
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 output_o[77]
port 497 nsew signal output
flabel metal2 s 30968 0 31048 80 0 FreeSans 320 0 0 0 output_o[78]
port 498 nsew signal output
flabel metal2 s 31352 0 31432 80 0 FreeSans 320 0 0 0 output_o[79]
port 499 nsew signal output
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 output_o[7]
port 500 nsew signal output
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 output_o[80]
port 501 nsew signal output
flabel metal2 s 32120 0 32200 80 0 FreeSans 320 0 0 0 output_o[81]
port 502 nsew signal output
flabel metal2 s 32504 0 32584 80 0 FreeSans 320 0 0 0 output_o[82]
port 503 nsew signal output
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 output_o[83]
port 504 nsew signal output
flabel metal2 s 33272 0 33352 80 0 FreeSans 320 0 0 0 output_o[84]
port 505 nsew signal output
flabel metal2 s 33656 0 33736 80 0 FreeSans 320 0 0 0 output_o[85]
port 506 nsew signal output
flabel metal2 s 34040 0 34120 80 0 FreeSans 320 0 0 0 output_o[86]
port 507 nsew signal output
flabel metal2 s 34424 0 34504 80 0 FreeSans 320 0 0 0 output_o[87]
port 508 nsew signal output
flabel metal2 s 34808 0 34888 80 0 FreeSans 320 0 0 0 output_o[88]
port 509 nsew signal output
flabel metal2 s 35192 0 35272 80 0 FreeSans 320 0 0 0 output_o[89]
port 510 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 output_o[8]
port 511 nsew signal output
flabel metal2 s 35576 0 35656 80 0 FreeSans 320 0 0 0 output_o[90]
port 512 nsew signal output
flabel metal2 s 35960 0 36040 80 0 FreeSans 320 0 0 0 output_o[91]
port 513 nsew signal output
flabel metal2 s 36344 0 36424 80 0 FreeSans 320 0 0 0 output_o[92]
port 514 nsew signal output
flabel metal2 s 36728 0 36808 80 0 FreeSans 320 0 0 0 output_o[93]
port 515 nsew signal output
flabel metal2 s 37112 0 37192 80 0 FreeSans 320 0 0 0 output_o[94]
port 516 nsew signal output
flabel metal2 s 37496 0 37576 80 0 FreeSans 320 0 0 0 output_o[95]
port 517 nsew signal output
flabel metal2 s 37880 0 37960 80 0 FreeSans 320 0 0 0 output_o[96]
port 518 nsew signal output
flabel metal2 s 38264 0 38344 80 0 FreeSans 320 0 0 0 output_o[97]
port 519 nsew signal output
flabel metal2 s 38648 0 38728 80 0 FreeSans 320 0 0 0 output_o[98]
port 520 nsew signal output
flabel metal2 s 39032 0 39112 80 0 FreeSans 320 0 0 0 output_o[99]
port 521 nsew signal output
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 output_o[9]
port 522 nsew signal output
rlabel metal1 49968 10584 49968 10584 0 VGND
rlabel metal1 49968 11340 49968 11340 0 VPWR
rlabel metal2 38304 8400 38304 8400 0 _000_
rlabel metal2 37728 5964 37728 5964 0 _001_
rlabel metal2 32304 8736 32304 8736 0 _002_
rlabel metal2 31200 6384 31200 6384 0 _003_
rlabel metal2 37344 6300 37344 6300 0 _004_
rlabel metal2 51648 7980 51648 7980 0 _005_
rlabel metal2 49440 6384 49440 6384 0 _006_
rlabel metal2 50976 6510 50976 6510 0 _007_
rlabel metal3 66960 6384 66960 6384 0 _008_
rlabel metal3 62496 6384 62496 6384 0 _009_
rlabel metal3 60816 6972 60816 6972 0 _010_
rlabel metal2 46368 6258 46368 6258 0 _011_
rlabel metal2 50496 8778 50496 8778 0 _012_
rlabel metal2 55392 5082 55392 5082 0 _013_
rlabel metal4 41568 6216 41568 6216 0 _014_
rlabel metal2 61344 5166 61344 5166 0 _015_
rlabel metal2 59424 7308 59424 7308 0 _016_
rlabel metal2 48768 8232 48768 8232 0 _017_
rlabel metal2 49632 4746 49632 4746 0 _018_
rlabel metal2 48288 8820 48288 8820 0 _019_
rlabel metal3 50304 4788 50304 4788 0 _020_
rlabel metal3 52272 4200 52272 4200 0 _021_
rlabel metal2 51360 7686 51360 7686 0 _022_
rlabel metal3 54144 5712 54144 5712 0 _023_
rlabel metal2 56784 8568 56784 8568 0 _024_
rlabel metal2 54864 8904 54864 8904 0 _025_
rlabel metal3 57024 7896 57024 7896 0 _026_
rlabel metal3 52128 7224 52128 7224 0 _027_
rlabel metal2 56736 6342 56736 6342 0 _028_
rlabel metal3 56352 5712 56352 5712 0 _029_
rlabel metal3 56352 4032 56352 4032 0 _030_
rlabel via1 56448 4957 56448 4957 0 _031_
rlabel metal3 57312 9576 57312 9576 0 _032_
rlabel metal2 58656 9870 58656 9870 0 _033_
rlabel metal2 57600 10290 57600 10290 0 _034_
rlabel via2 35901 6384 35901 6384 0 _035_
rlabel metal2 72096 8022 72096 8022 0 _036_
rlabel metal2 67584 6468 67584 6468 0 _037_
rlabel metal2 44928 8778 44928 8778 0 _038_
rlabel metal2 44352 4746 44352 4746 0 _039_
rlabel metal3 43728 7896 43728 7896 0 _040_
rlabel metal2 45600 4998 45600 4998 0 _041_
rlabel metal2 45216 7938 45216 7938 0 _042_
rlabel metal3 45744 4704 45744 4704 0 _043_
rlabel metal2 44352 7434 44352 7434 0 _044_
rlabel metal2 44256 5250 44256 5250 0 _045_
rlabel metal2 40896 8190 40896 8190 0 _046_
rlabel metal2 48528 4200 48528 4200 0 _047_
rlabel metal2 46272 8904 46272 8904 0 _048_
rlabel metal2 45984 4284 45984 4284 0 _049_
rlabel metal2 41376 7476 41376 7476 0 _050_
rlabel metal2 47520 3150 47520 3150 0 _051_
rlabel metal4 46368 7098 46368 7098 0 _052_
rlabel metal3 48144 4200 48144 4200 0 _053_
rlabel metal2 40320 9366 40320 9366 0 _054_
rlabel metal2 40224 6510 40224 6510 0 _055_
rlabel metal2 41568 10332 41568 10332 0 _056_
rlabel metal2 42624 5544 42624 5544 0 _057_
rlabel metal2 48672 10122 48672 10122 0 _058_
rlabel metal2 44352 6216 44352 6216 0 _059_
rlabel metal2 41568 9198 41568 9198 0 _060_
rlabel metal3 43152 6384 43152 6384 0 _061_
rlabel metal2 51168 9996 51168 9996 0 _062_
rlabel metal2 51456 6720 51456 6720 0 _063_
rlabel metal2 53472 9744 53472 9744 0 _064_
rlabel metal2 42864 6384 42864 6384 0 _065_
rlabel metal2 53088 10374 53088 10374 0 _066_
rlabel metal4 51840 7140 51840 7140 0 _067_
rlabel metal2 44640 8568 44640 8568 0 _068_
rlabel metal2 46656 5460 46656 5460 0 _069_
rlabel metal2 37920 6342 37920 6342 0 _070_
rlabel metal3 75504 8148 75504 8148 0 _071_
rlabel metal2 72768 6132 72768 6132 0 _072_
rlabel metal2 84672 6720 84672 6720 0 _073_
rlabel metal2 78624 8652 78624 8652 0 _074_
rlabel metal3 77712 4872 77712 4872 0 _075_
rlabel metal3 87552 7266 87552 7266 0 _076_
rlabel metal2 78432 4830 78432 4830 0 _077_
rlabel metal2 86688 6342 86688 6342 0 _078_
rlabel metal2 84576 5166 84576 5166 0 _079_
rlabel metal2 85632 7308 85632 7308 0 _080_
rlabel metal3 74736 5712 74736 5712 0 _081_
rlabel metal2 17184 7560 17184 7560 0 _082_
rlabel metal2 17184 4494 17184 4494 0 _083_
rlabel metal2 15744 8652 15744 8652 0 _084_
rlabel metal2 18240 4998 18240 4998 0 _085_
rlabel metal2 20640 7854 20640 7854 0 _086_
rlabel metal2 24288 6300 24288 6300 0 _087_
rlabel metal2 33888 8736 33888 8736 0 _088_
rlabel metal2 34080 8568 34080 8568 0 _089_
rlabel metal2 29184 6090 29184 6090 0 _090_
rlabel metal3 29904 8736 29904 8736 0 _091_
rlabel metal2 30144 6132 30144 6132 0 _092_
rlabel metal2 37104 8148 37104 8148 0 _093_
rlabel metal2 35712 5712 35712 5712 0 _094_
rlabel metal2 6240 13430 6240 13430 0 ena_i
rlabel metal2 17184 13136 17184 13136 0 input_ni[0]
rlabel metal2 28128 13136 28128 13136 0 input_ni[1]
rlabel metal2 39072 12926 39072 12926 0 input_ni[2]
rlabel metal2 50016 13136 50016 13136 0 input_ni[3]
rlabel metal2 60960 13136 60960 13136 0 input_ni[4]
rlabel metal2 71904 13136 71904 13136 0 input_ni[5]
rlabel metal2 82848 13136 82848 13136 0 input_ni[6]
rlabel metal2 93792 13430 93792 13430 0 input_ni[7]
rlabel metal2 19968 4452 19968 4452 0 net1
rlabel metal3 37008 9408 37008 9408 0 net10
rlabel metal2 60384 9240 60384 9240 0 net100
rlabel metal2 54816 4536 54816 4536 0 net101
rlabel metal2 58464 7980 58464 7980 0 net102
rlabel via1 57600 4193 57600 4193 0 net103
rlabel metal2 58176 10416 58176 10416 0 net104
rlabel metal2 58944 7140 58944 7140 0 net105
rlabel metal2 52608 6930 52608 6930 0 net106
rlabel metal2 53280 5628 53280 5628 0 net107
rlabel metal2 46560 4116 46560 4116 0 net108
rlabel metal2 55008 9114 55008 9114 0 net109
rlabel metal2 31104 5796 31104 5796 0 net11
rlabel metal2 46176 4914 46176 4914 0 net110
rlabel metal2 51744 7182 51744 7182 0 net111
rlabel metal2 56544 9114 56544 9114 0 net112
rlabel metal2 49344 9408 49344 9408 0 net113
rlabel metal2 45120 7602 45120 7602 0 net114
rlabel metal2 50784 8190 50784 8190 0 net115
rlabel metal2 45216 5754 45216 5754 0 net116
rlabel metal2 49920 5166 49920 5166 0 net117
rlabel metal2 44640 7098 44640 7098 0 net118
rlabel metal2 52560 8736 52560 8736 0 net119
rlabel metal3 31248 5712 31248 5712 0 net12
rlabel metal2 29760 7371 29760 7371 0 net120
rlabel metal3 36432 6972 36432 6972 0 net121
rlabel metal2 39456 7392 39456 7392 0 net122
rlabel metal3 44736 6300 44736 6300 0 net123
rlabel metal2 45408 5586 45408 5586 0 net124
rlabel metal2 47328 4914 47328 4914 0 net125
rlabel metal2 45984 7308 45984 7308 0 net126
rlabel metal3 51744 9240 51744 9240 0 net127
rlabel metal2 62016 6174 62016 6174 0 net128
rlabel metal2 50688 6552 50688 6552 0 net129
rlabel metal3 28416 8736 28416 8736 0 net13
rlabel metal3 38016 4200 38016 4200 0 net130
rlabel metal3 38784 5670 38784 5670 0 net131
rlabel metal3 41376 5880 41376 5880 0 net132
rlabel metal2 68928 5670 68928 5670 0 net133
rlabel metal2 37920 9534 37920 9534 0 net134
rlabel metal2 66240 7770 66240 7770 0 net135
rlabel via1 38401 4200 38401 4200 0 net136
rlabel metal2 69120 4116 69120 4116 0 net137
rlabel metal2 39120 4200 39120 4200 0 net138
rlabel metal2 68352 4830 68352 4830 0 net139
rlabel metal2 30432 9408 30432 9408 0 net14
rlabel metal2 39840 5040 39840 5040 0 net140
rlabel metal2 68544 4368 68544 4368 0 net141
rlabel metal2 35232 4284 35232 4284 0 net142
rlabel metal2 66912 4494 66912 4494 0 net143
rlabel metal2 38688 4830 38688 4830 0 net144
rlabel metal2 67200 4914 67200 4914 0 net145
rlabel metal2 38304 3948 38304 3948 0 net146
rlabel metal2 53664 4326 53664 4326 0 net147
rlabel metal2 38016 3948 38016 3948 0 net148
rlabel metal2 55008 4578 55008 4578 0 net149
rlabel metal3 28752 5712 28752 5712 0 net15
rlabel metal2 67344 4872 67344 4872 0 net150
rlabel metal3 68400 7224 68400 7224 0 net151
rlabel metal2 29952 6405 29952 6405 0 net152
rlabel metal2 81888 5670 81888 5670 0 net153
rlabel metal3 78432 2016 78432 2016 0 net154
rlabel metal4 17472 10164 17472 10164 0 net155
rlabel metal3 39168 11424 39168 11424 0 net156
rlabel metal2 39264 9198 39264 9198 0 net157
rlabel metal2 51264 9324 51264 9324 0 net158
rlabel metal2 39744 7980 39744 7980 0 net159
rlabel metal3 28032 6384 28032 6384 0 net16
rlabel metal2 39552 7602 39552 7602 0 net160
rlabel metal4 45696 6468 45696 6468 0 net161
rlabel metal2 10176 6720 10176 6720 0 net162
rlabel metal2 37248 3738 37248 3738 0 net163
rlabel metal2 37584 3444 37584 3444 0 net164
rlabel metal2 38352 5040 38352 5040 0 net165
rlabel metal2 40272 4956 40272 4956 0 net166
rlabel metal2 39600 5208 39600 5208 0 net167
rlabel metal2 40608 6846 40608 6846 0 net168
rlabel metal2 39984 4116 39984 4116 0 net169
rlabel metal3 24480 8736 24480 8736 0 net17
rlabel metal4 37824 3822 37824 3822 0 net170
rlabel metal2 41376 5628 41376 5628 0 net171
rlabel metal2 40752 8148 40752 8148 0 net172
rlabel metal2 18720 9744 18720 9744 0 net173
rlabel metal5 39504 3780 39504 3780 0 net174
rlabel metal2 42912 5964 42912 5964 0 net175
rlabel metal4 41472 5922 41472 5922 0 net176
rlabel metal4 39936 5628 39936 5628 0 net177
rlabel metal4 30912 6720 30912 6720 0 net178
rlabel metal2 42192 4116 42192 4116 0 net179
rlabel metal3 24912 9408 24912 9408 0 net18
rlabel metal4 42624 6048 42624 6048 0 net180
rlabel metal4 36672 4956 36672 4956 0 net181
rlabel metal4 43392 5964 43392 5964 0 net182
rlabel metal5 42280 3486 42280 3486 0 net183
rlabel metal4 16224 9114 16224 9114 0 net184
rlabel metal2 38880 9198 38880 9198 0 net185
rlabel metal2 37536 9744 37536 9744 0 net186
rlabel metal3 38496 9282 38496 9282 0 net187
rlabel metal2 39072 9072 39072 9072 0 net188
rlabel metal2 38688 9156 38688 9156 0 net189
rlabel metal2 24960 5292 24960 5292 0 net19
rlabel metal2 38208 8568 38208 8568 0 net190
rlabel metal4 48384 7518 48384 7518 0 net191
rlabel metal2 38112 9240 38112 9240 0 net192
rlabel metal2 48384 3108 48384 3108 0 net193
rlabel metal2 51264 4074 51264 4074 0 net194
rlabel metal2 7392 8148 7392 8148 0 net195
rlabel metal2 50496 3486 50496 3486 0 net196
rlabel metal2 51456 3486 51456 3486 0 net197
rlabel metal2 52224 3570 52224 3570 0 net198
rlabel metal2 55392 6258 55392 6258 0 net199
rlabel metal3 30432 5586 30432 5586 0 net2
rlabel via1 24970 6384 24970 6384 0 net20
rlabel metal2 53904 3444 53904 3444 0 net200
rlabel metal2 53952 4452 53952 4452 0 net201
rlabel metal2 55296 3612 55296 3612 0 net202
rlabel metal2 56064 3528 56064 3528 0 net203
rlabel metal2 56448 3696 56448 3696 0 net204
rlabel metal2 56832 3318 56832 3318 0 net205
rlabel metal2 12288 7602 12288 7602 0 net206
rlabel metal2 55776 4746 55776 4746 0 net207
rlabel metal3 57888 10080 57888 10080 0 net208
rlabel metal2 58032 9996 58032 9996 0 net209
rlabel metal2 19968 7847 19968 7847 0 net21
rlabel metal2 58944 3276 58944 3276 0 net210
rlabel metal2 58848 4662 58848 4662 0 net211
rlabel metal4 58272 4452 58272 4452 0 net212
rlabel metal2 49872 3612 49872 3612 0 net213
rlabel metal2 53184 4746 53184 4746 0 net214
rlabel metal2 54624 6090 54624 6090 0 net215
rlabel metal2 59520 6300 59520 6300 0 net216
rlabel metal2 12528 9996 12528 9996 0 net217
rlabel metal3 57552 9072 57552 9072 0 net218
rlabel metal2 59856 5628 59856 5628 0 net219
rlabel metal3 19680 9408 19680 9408 0 net22
rlabel metal2 62304 3486 62304 3486 0 net220
rlabel metal2 60288 5586 60288 5586 0 net221
rlabel metal2 56736 4410 56736 4410 0 net222
rlabel metal3 62502 3444 62502 3444 0 net223
rlabel metal2 63696 3444 63696 3444 0 net224
rlabel metal2 62784 4998 62784 4998 0 net225
rlabel metal2 62448 5628 62448 5628 0 net226
rlabel metal2 61824 5166 61824 5166 0 net227
rlabel metal4 9024 9366 9024 9366 0 net228
rlabel metal2 69984 6090 69984 6090 0 net229
rlabel metal2 19008 4746 19008 4746 0 net23
rlabel metal2 65568 3906 65568 3906 0 net230
rlabel metal2 70080 9030 70080 9030 0 net231
rlabel metal2 65280 5040 65280 5040 0 net232
rlabel metal2 66336 3486 66336 3486 0 net233
rlabel metal2 66720 3402 66720 3402 0 net234
rlabel metal2 67104 3402 67104 3402 0 net235
rlabel metal3 70752 8820 70752 8820 0 net236
rlabel metal2 67872 3612 67872 3612 0 net237
rlabel metal2 68256 3192 68256 3192 0 net238
rlabel metal2 6528 5544 6528 5544 0 net239
rlabel metal2 19440 5712 19440 5712 0 net24
rlabel metal2 66912 7224 66912 7224 0 net240
rlabel metal2 69024 3780 69024 3780 0 net241
rlabel metal2 71424 8190 71424 8190 0 net242
rlabel metal2 67872 5712 67872 5712 0 net243
rlabel metal4 69504 6888 69504 6888 0 net244
rlabel metal2 70570 3353 70570 3353 0 net245
rlabel metal2 70080 6048 70080 6048 0 net246
rlabel metal2 71808 3444 71808 3444 0 net247
rlabel metal2 71232 7602 71232 7602 0 net248
rlabel metal4 72960 5880 72960 5880 0 net249
rlabel metal2 12000 8022 12000 8022 0 net25
rlabel metal2 6912 5208 6912 5208 0 net250
rlabel metal2 71904 5376 71904 5376 0 net251
rlabel metal3 73824 8988 73824 8988 0 net252
rlabel via2 73068 8904 73068 8904 0 net253
rlabel metal2 73632 4158 73632 4158 0 net254
rlabel metal2 74400 3780 74400 3780 0 net255
rlabel metal2 74112 4368 74112 4368 0 net256
rlabel metal2 73728 6930 73728 6930 0 net257
rlabel metal2 75552 3612 75552 3612 0 net258
rlabel metal4 75264 6846 75264 6846 0 net259
rlabel metal2 11808 10836 11808 10836 0 net26
rlabel metal4 75648 7056 75648 7056 0 net260
rlabel metal3 8928 4116 8928 4116 0 net261
rlabel metal2 76992 3444 76992 3444 0 net262
rlabel metal2 77472 4284 77472 4284 0 net263
rlabel metal2 77904 3444 77904 3444 0 net264
rlabel metal2 76320 6720 76320 6720 0 net265
rlabel metal2 75744 6972 75744 6972 0 net266
rlabel metal2 79008 3612 79008 3612 0 net267
rlabel metal3 77712 5628 77712 5628 0 net268
rlabel metal2 79776 3402 79776 3402 0 net269
rlabel metal2 18576 4872 18576 4872 0 net27
rlabel metal2 79392 4410 79392 4410 0 net270
rlabel metal2 78960 4956 78960 4956 0 net271
rlabel metal2 7680 4200 7680 4200 0 net272
rlabel metal2 9600 6510 9600 6510 0 net273
rlabel metal3 80832 3444 80832 3444 0 net274
rlabel metal2 82272 7938 82272 7938 0 net275
rlabel metal2 82656 6426 82656 6426 0 net276
rlabel metal4 82272 7770 82272 7770 0 net277
rlabel metal3 82464 3444 82464 3444 0 net278
rlabel metal2 83280 3444 83280 3444 0 net279
rlabel metal2 16896 5754 16896 5754 0 net28
rlabel metal2 83904 8736 83904 8736 0 net280
rlabel metal2 82176 4830 82176 4830 0 net281
rlabel metal3 82080 5922 82080 5922 0 net282
rlabel metal3 83136 6678 83136 6678 0 net283
rlabel metal3 11526 7812 11526 7812 0 net284
rlabel metal2 84912 6048 84912 6048 0 net285
rlabel metal3 83139 6216 83139 6216 0 net286
rlabel metal2 86256 3444 86256 3444 0 net287
rlabel metal2 86016 8190 86016 8190 0 net288
rlabel metal2 86784 8904 86784 8904 0 net289
rlabel metal2 12096 7098 12096 7098 0 net29
rlabel metal2 85920 6636 85920 6636 0 net290
rlabel metal2 87504 3444 87504 3444 0 net291
rlabel metal2 86256 4956 86256 4956 0 net292
rlabel metal2 87840 3486 87840 3486 0 net293
rlabel metal2 86592 5250 86592 5250 0 net294
rlabel metal2 8448 6174 8448 6174 0 net295
rlabel metal2 88224 3696 88224 3696 0 net296
rlabel metal2 86976 4998 86976 4998 0 net297
rlabel metal2 89376 9240 89376 9240 0 net298
rlabel metal2 87360 5964 87360 5964 0 net299
rlabel metal3 11712 8736 11712 8736 0 net3
rlabel metal2 15360 9240 15360 9240 0 net30
rlabel metal2 88992 3738 88992 3738 0 net300
rlabel metal2 88608 5418 88608 5418 0 net301
rlabel metal3 88224 4956 88224 4956 0 net302
rlabel metal2 89904 3444 89904 3444 0 net303
rlabel metal2 89376 5838 89376 5838 0 net304
rlabel metal2 89760 4200 89760 4200 0 net305
rlabel metal2 12000 6006 12000 6006 0 net306
rlabel metal2 90144 6258 90144 6258 0 net307
rlabel metal2 90528 5586 90528 5586 0 net308
rlabel metal2 89568 7056 89568 7056 0 net309
rlabel metal2 87072 8442 87072 8442 0 net31
rlabel metal2 89760 6762 89760 6762 0 net310
rlabel metal2 89856 6342 89856 6342 0 net311
rlabel metal2 87744 8904 87744 8904 0 net312
rlabel metal2 92448 7182 92448 7182 0 net313
rlabel metal2 88320 10416 88320 10416 0 net314
rlabel metal2 93216 7098 93216 7098 0 net315
rlabel metal2 86880 4704 86880 4704 0 net316
rlabel metal2 12672 5838 12672 5838 0 net317
rlabel metal2 93984 6090 93984 6090 0 net318
rlabel metal2 94272 6552 94272 6552 0 net319
rlabel metal2 86832 7896 86832 7896 0 net32
rlabel metal4 86880 5712 86880 5712 0 net320
rlabel metal3 86112 4158 86112 4158 0 net321
rlabel metal2 87648 7476 87648 7476 0 net322
rlabel metal2 86592 6384 86592 6384 0 net323
rlabel metal2 84096 7686 84096 7686 0 net324
rlabel metal2 96672 5964 96672 5964 0 net325
rlabel metal2 89184 7728 89184 7728 0 net326
rlabel metal2 97440 6474 97440 6474 0 net327
rlabel metal2 9216 7308 9216 7308 0 net328
rlabel metal2 89856 9240 89856 9240 0 net329
rlabel metal2 84480 4116 84480 4116 0 net33
rlabel metal2 86976 8862 86976 8862 0 net330
rlabel metal2 97248 6762 97248 6762 0 net331
rlabel metal2 88704 5880 88704 5880 0 net332
rlabel metal2 97920 7476 97920 7476 0 net333
rlabel metal2 85728 7350 85728 7350 0 net334
rlabel metal2 9600 8526 9600 8526 0 net335
rlabel metal2 15264 7728 15264 7728 0 net336
rlabel metal3 13248 10836 13248 10836 0 net337
rlabel metal2 12096 10416 12096 10416 0 net338
rlabel metal3 11568 9576 11568 9576 0 net339
rlabel metal3 83904 4872 83904 4872 0 net34
rlabel metal2 1728 4872 1728 4872 0 net340
rlabel metal2 11808 8694 11808 8694 0 net341
rlabel metal2 12288 5334 12288 5334 0 net342
rlabel metal2 13056 8442 13056 8442 0 net343
rlabel metal2 13728 5544 13728 5544 0 net344
rlabel metal2 12384 4032 12384 4032 0 net345
rlabel metal2 13344 5880 13344 5880 0 net346
rlabel metal2 14304 6384 14304 6384 0 net347
rlabel metal2 13152 5292 13152 5292 0 net348
rlabel metal2 14208 5754 14208 5754 0 net349
rlabel metal2 88809 7847 88809 7847 0 net35
rlabel metal2 15072 5670 15072 5670 0 net350
rlabel metal2 1632 4494 1632 4494 0 net351
rlabel metal2 13920 4116 13920 4116 0 net352
rlabel metal2 14976 5586 14976 5586 0 net353
rlabel metal2 15264 4116 15264 4116 0 net354
rlabel metal2 16416 5460 16416 5460 0 net355
rlabel metal3 13104 9156 13104 9156 0 net356
rlabel metal2 16128 4578 16128 4578 0 net357
rlabel metal2 14496 10374 14496 10374 0 net358
rlabel metal4 16224 5082 16224 5082 0 net359
rlabel metal2 87840 7182 87840 7182 0 net36
rlabel metal2 19488 6510 19488 6510 0 net360
rlabel metal3 16896 3444 16896 3444 0 net361
rlabel metal2 1968 4116 1968 4116 0 net362
rlabel metal4 17472 5628 17472 5628 0 net363
rlabel metal2 20736 6720 20736 6720 0 net364
rlabel metal2 19488 7266 19488 7266 0 net365
rlabel metal2 19104 7434 19104 7434 0 net366
rlabel metal2 18912 3486 18912 3486 0 net367
rlabel metal4 19296 5418 19296 5418 0 net368
rlabel metal2 19680 4830 19680 4830 0 net369
rlabel metal3 71952 4872 71952 4872 0 net37
rlabel metal2 21504 5586 21504 5586 0 net370
rlabel metal2 21360 5040 21360 5040 0 net371
rlabel metal4 19872 7014 19872 7014 0 net372
rlabel metal2 2352 4116 2352 4116 0 net373
rlabel metal2 19488 9744 19488 9744 0 net374
rlabel metal3 21504 9324 21504 9324 0 net375
rlabel metal2 19104 10500 19104 10500 0 net376
rlabel metal2 19104 9072 19104 9072 0 net377
rlabel metal2 23808 3444 23808 3444 0 net378
rlabel metal2 24384 3444 24384 3444 0 net379
rlabel metal2 85488 4200 85488 4200 0 net38
rlabel metal2 26112 5670 26112 5670 0 net380
rlabel metal4 25728 5670 25728 5670 0 net381
rlabel metal2 24960 3444 24960 3444 0 net382
rlabel metal2 26880 6888 26880 6888 0 net383
rlabel metal2 2688 4158 2688 4158 0 net384
rlabel metal2 26544 4116 26544 4116 0 net385
rlabel metal2 25824 3738 25824 3738 0 net386
rlabel metal2 26880 4158 26880 4158 0 net387
rlabel metal2 26592 3528 26592 3528 0 net388
rlabel metal2 29568 6510 29568 6510 0 net389
rlabel via2 81119 7896 81119 7896 0 net39
rlabel metal2 29664 7560 29664 7560 0 net390
rlabel metal2 29280 8106 29280 8106 0 net391
rlabel metal2 28800 4158 28800 4158 0 net392
rlabel metal3 26208 9324 26208 9324 0 net393
rlabel metal2 28512 3570 28512 3570 0 net394
rlabel metal2 12384 8946 12384 8946 0 net395
rlabel metal2 29280 3612 29280 3612 0 net396
rlabel metal2 30048 3402 30048 3402 0 net397
rlabel metal4 31488 4536 31488 4536 0 net398
rlabel metal2 30816 3948 30816 3948 0 net399
rlabel metal2 18816 10332 18816 10332 0 net4
rlabel metal2 88800 9324 88800 9324 0 net40
rlabel metal2 32640 8316 32640 8316 0 net400
rlabel metal4 31680 6552 31680 6552 0 net401
rlabel metal2 33408 7560 33408 7560 0 net402
rlabel metal3 30048 5712 30048 5712 0 net403
rlabel metal3 31632 8064 31632 8064 0 net404
rlabel metal3 33696 4956 33696 4956 0 net405
rlabel metal2 3456 7056 3456 7056 0 net406
rlabel metal2 35712 7350 35712 7350 0 net407
rlabel metal2 34176 5040 34176 5040 0 net408
rlabel metal2 33120 3402 33120 3402 0 net409
rlabel metal2 77184 4158 77184 4158 0 net41
rlabel metal2 30240 9240 30240 9240 0 net410
rlabel metal2 35328 3612 35328 3612 0 net411
rlabel metal3 35952 8988 35952 8988 0 net412
rlabel metal2 36480 4542 36480 4542 0 net413
rlabel metal4 36096 4662 36096 4662 0 net414
rlabel metal2 37968 4956 37968 4956 0 net415
rlabel metal4 37248 6426 37248 6426 0 net416
rlabel metal2 7488 7518 7488 7518 0 net417
rlabel metal3 33852 1344 33852 1344 0 net418
rlabel metal2 35424 4872 35424 4872 0 net419
rlabel metal2 79440 4872 79440 4872 0 net42
rlabel metal2 40128 5124 40128 5124 0 net420
rlabel metal4 36576 3948 36576 3948 0 net421
rlabel metal2 38784 3612 38784 3612 0 net422
rlabel metal2 41280 5796 41280 5796 0 net423
rlabel metal2 39168 3276 39168 3276 0 net424
rlabel metal2 40992 4998 40992 4998 0 net425
rlabel metal3 40464 4116 40464 4116 0 net426
rlabel metal2 39936 3318 39936 3318 0 net427
rlabel metal2 41760 5208 41760 5208 0 net428
rlabel metal3 14304 5502 14304 5502 0 net429
rlabel metal2 78432 8904 78432 8904 0 net43
rlabel metal3 40992 4116 40992 4116 0 net430
rlabel metal4 39744 4074 39744 4074 0 net431
rlabel metal3 38448 3948 38448 3948 0 net432
rlabel metal2 41856 4410 41856 4410 0 net433
rlabel metal2 41472 3654 41472 3654 0 net434
rlabel metal2 38976 3696 38976 3696 0 net435
rlabel metal3 37824 3906 37824 3906 0 net436
rlabel metal2 39552 3822 39552 3822 0 net437
rlabel metal3 43008 3906 43008 3906 0 net438
rlabel metal3 40086 4032 40086 4032 0 net439
rlabel metal2 82080 9450 82080 9450 0 net44
rlabel metal3 15840 5670 15840 5670 0 net440
rlabel metal3 42912 5208 42912 5208 0 net441
rlabel metal2 44496 3444 44496 3444 0 net442
rlabel metal2 44928 2940 44928 2940 0 net443
rlabel metal2 39264 3570 39264 3570 0 net444
rlabel metal2 38112 5376 38112 5376 0 net445
rlabel metal3 38736 6048 38736 6048 0 net446
rlabel metal4 38208 5502 38208 5502 0 net447
rlabel metal5 41580 3402 41580 3402 0 net448
rlabel metal2 48768 3276 48768 3276 0 net449
rlabel metal3 70560 5712 70560 5712 0 net45
rlabel metal2 50880 4410 50880 4410 0 net450
rlabel metal4 6240 4872 6240 4872 0 net451
rlabel metal2 50832 3444 50832 3444 0 net452
rlabel metal3 52128 3444 52128 3444 0 net453
rlabel metal2 53232 3444 53232 3444 0 net454
rlabel metal2 52896 7056 52896 7056 0 net455
rlabel metal2 54288 3444 54288 3444 0 net456
rlabel metal2 54720 7518 54720 7518 0 net457
rlabel metal2 55728 3444 55728 3444 0 net458
rlabel metal3 56256 4116 56256 4116 0 net459
rlabel metal2 74064 5712 74064 5712 0 net46
rlabel metal2 56064 4200 56064 4200 0 net460
rlabel metal3 55176 5628 55176 5628 0 net461
rlabel metal3 16512 5418 16512 5418 0 net462
rlabel metal2 55296 5838 55296 5838 0 net463
rlabel metal4 58176 4368 58176 4368 0 net464
rlabel metal2 58560 3654 58560 3654 0 net465
rlabel metal2 62496 6888 62496 6888 0 net466
rlabel metal2 55200 4410 55200 4410 0 net467
rlabel metal4 49536 3738 49536 3738 0 net468
rlabel metal4 58080 4746 58080 4746 0 net469
rlabel metal3 75360 8736 75360 8736 0 net47
rlabel metal2 53376 3822 53376 3822 0 net470
rlabel metal4 54144 3570 54144 3570 0 net471
rlabel metal2 58848 7098 58848 7098 0 net472
rlabel metal2 5472 5292 5472 5292 0 net473
rlabel metal4 54912 5334 54912 5334 0 net474
rlabel metal2 60768 5502 60768 5502 0 net475
rlabel metal2 61632 4410 61632 4410 0 net476
rlabel metal4 62016 4998 62016 4998 0 net477
rlabel metal2 62400 4284 62400 4284 0 net478
rlabel metal2 62784 4368 62784 4368 0 net479
rlabel metal2 76416 8736 76416 8736 0 net48
rlabel metal2 60768 8400 60768 8400 0 net480
rlabel metal2 64320 3192 64320 3192 0 net481
rlabel metal2 64800 3360 64800 3360 0 net482
rlabel metal3 63552 3570 63552 3570 0 net483
rlabel metal3 8406 2436 8406 2436 0 net484
rlabel metal2 67584 5208 67584 5208 0 net485
rlabel metal3 67536 3948 67536 3948 0 net486
rlabel metal3 66480 3444 66480 3444 0 net487
rlabel metal2 67776 3906 67776 3906 0 net488
rlabel metal2 65664 4158 65664 4158 0 net489
rlabel metal3 38640 6384 38640 6384 0 net49
rlabel metal3 66144 4116 66144 4116 0 net490
rlabel metal3 67440 4116 67440 4116 0 net491
rlabel metal3 67536 4368 67536 4368 0 net492
rlabel metal2 66528 5208 66528 5208 0 net493
rlabel metal2 67632 4116 67632 4116 0 net494
rlabel metal3 6078 2352 6078 2352 0 net495
rlabel metal2 68544 3444 68544 3444 0 net496
rlabel metal3 67584 5628 67584 5628 0 net497
rlabel metal2 69792 4074 69792 4074 0 net498
rlabel metal2 70128 3444 70128 3444 0 net499
rlabel metal2 33120 7854 33120 7854 0 net5
rlabel metal2 68976 7224 68976 7224 0 net50
rlabel metal2 68928 5208 68928 5208 0 net500
rlabel metal2 69888 4326 69888 4326 0 net501
rlabel metal2 70944 3528 70944 3528 0 net502
rlabel metal3 70032 4032 70032 4032 0 net503
rlabel metal2 72096 3486 72096 3486 0 net504
rlabel metal3 70320 4956 70320 4956 0 net505
rlabel metal3 14400 2100 14400 2100 0 net506
rlabel metal2 70944 4536 70944 4536 0 net507
rlabel metal2 70560 5292 70560 5292 0 net508
rlabel metal3 71952 4116 71952 4116 0 net509
rlabel metal2 38016 10542 38016 10542 0 net51
rlabel metal2 69792 5376 69792 5376 0 net510
rlabel metal2 74784 4830 74784 4830 0 net511
rlabel metal3 74688 3444 74688 3444 0 net512
rlabel metal2 74544 4116 74544 4116 0 net513
rlabel metal2 75936 3491 75936 3491 0 net514
rlabel metal4 76320 5040 76320 5040 0 net515
rlabel metal2 76704 3528 76704 3528 0 net516
rlabel metal3 10560 1890 10560 1890 0 net517
rlabel metal3 76272 4116 76272 4116 0 net518
rlabel metal3 74544 5628 74544 5628 0 net519
rlabel metal2 83232 10290 83232 10290 0 net52
rlabel metal2 78240 3486 78240 3486 0 net520
rlabel metal2 72576 3612 72576 3612 0 net521
rlabel metal2 76704 5754 76704 5754 0 net522
rlabel metal2 72768 4368 72768 4368 0 net523
rlabel metal3 79104 3444 79104 3444 0 net524
rlabel metal2 78528 4998 78528 4998 0 net525
rlabel metal4 80160 4494 80160 4494 0 net526
rlabel metal2 79776 4788 79776 4788 0 net527
rlabel metal4 7008 3528 7008 3528 0 net528
rlabel metal4 35808 4536 35808 4536 0 net529
rlabel metal2 41952 6762 41952 6762 0 net53
rlabel metal2 80160 5292 80160 5292 0 net530
rlabel metal2 79872 4998 79872 4998 0 net531
rlabel metal2 80592 4956 80592 4956 0 net532
rlabel metal2 79152 5544 79152 5544 0 net533
rlabel metal2 79392 5964 79392 5964 0 net534
rlabel metal2 82656 4662 82656 4662 0 net535
rlabel metal3 78720 5418 78720 5418 0 net536
rlabel metal2 83040 4578 83040 4578 0 net537
rlabel metal2 82560 4536 82560 4536 0 net538
rlabel metal3 80352 2142 80352 2142 0 net539
rlabel metal2 68256 7182 68256 7182 0 net54
rlabel metal3 8352 2940 8352 2940 0 net540
rlabel metal3 71808 5040 71808 5040 0 net541
rlabel metal2 81312 1638 81312 1638 0 net542
rlabel metal2 85920 3990 85920 3990 0 net543
rlabel metal4 73728 4620 73728 4620 0 net544
rlabel metal2 85056 5208 85056 5208 0 net545
rlabel metal2 86592 4368 86592 4368 0 net546
rlabel metal2 85440 6090 85440 6090 0 net547
rlabel metal3 86112 3612 86112 3612 0 net548
rlabel metal2 85824 5586 85824 5586 0 net549
rlabel metal2 38400 10332 38400 10332 0 net55
rlabel metal2 87456 4284 87456 4284 0 net550
rlabel metal3 14016 3150 14016 3150 0 net551
rlabel metal3 84432 5628 84432 5628 0 net552
rlabel metal2 87840 5166 87840 5166 0 net553
rlabel metal2 85440 4452 85440 4452 0 net554
rlabel metal3 86112 4914 86112 4914 0 net555
rlabel metal4 72576 4872 72576 4872 0 net556
rlabel metal3 81312 1722 81312 1722 0 net557
rlabel metal2 88992 4416 88992 4416 0 net558
rlabel metal4 88512 4872 88512 4872 0 net559
rlabel metal3 83136 10248 83136 10248 0 net56
rlabel metal3 85584 2100 85584 2100 0 net560
rlabel metal3 81312 2352 81312 2352 0 net561
rlabel metal2 18624 4116 18624 4116 0 net562
rlabel metal2 86688 2772 86688 2772 0 net563
rlabel metal3 81792 2814 81792 2814 0 net564
rlabel metal3 87936 3486 87936 3486 0 net565
rlabel metal2 86880 3444 86880 3444 0 net566
rlabel metal2 83136 5334 83136 5334 0 net567
rlabel metal3 88704 3024 88704 3024 0 net568
rlabel metal3 82368 5418 82368 5418 0 net569
rlabel metal2 37920 5586 37920 5586 0 net57
rlabel metal3 84768 6132 84768 6132 0 net570
rlabel metal2 89664 5838 89664 5838 0 net571
rlabel metal3 89280 3234 89280 3234 0 net572
rlabel metal3 13344 2982 13344 2982 0 net573
rlabel metal4 60288 3402 60288 3402 0 net574
rlabel metal5 75120 3192 75120 3192 0 net575
rlabel metal4 64800 3780 64800 3780 0 net576
rlabel metal4 67104 3696 67104 3696 0 net577
rlabel metal2 88608 2856 88608 2856 0 net578
rlabel metal5 64260 3486 64260 3486 0 net579
rlabel metal2 69696 6468 69696 6468 0 net58
rlabel metal4 81888 3234 81888 3234 0 net580
rlabel metal3 68640 3654 68640 3654 0 net581
rlabel metal4 97824 4872 97824 4872 0 net582
rlabel metal2 83424 3822 83424 3822 0 net583
rlabel metal2 16128 5376 16128 5376 0 net584
rlabel metal4 82368 6468 82368 6468 0 net585
rlabel metal4 80640 5208 80640 5208 0 net586
rlabel metal4 81888 5166 81888 5166 0 net587
rlabel metal2 98496 5544 98496 5544 0 net588
rlabel metal2 83808 4620 83808 4620 0 net589
rlabel metal2 38784 10374 38784 10374 0 net59
rlabel metal5 82608 5544 82608 5544 0 net590
rlabel metal2 15744 5292 15744 5292 0 net591
rlabel metal2 9696 4662 9696 4662 0 net592
rlabel metal3 15744 3360 15744 3360 0 net593
rlabel metal2 13920 2982 13920 2982 0 net594
rlabel metal2 15168 3528 15168 3528 0 net595
rlabel metal2 34416 4032 34416 4032 0 net596
rlabel metal2 15360 5250 15360 5250 0 net597
rlabel metal2 11616 4326 11616 4326 0 net598
rlabel metal2 12000 3528 12000 3528 0 net599
rlabel metal2 38400 9072 38400 9072 0 net6
rlabel metal2 71328 10332 71328 10332 0 net60
rlabel metal4 17376 4368 17376 4368 0 net600
rlabel metal3 17760 3990 17760 3990 0 net601
rlabel metal3 12960 1680 12960 1680 0 net602
rlabel metal2 13824 4242 13824 4242 0 net603
rlabel metal3 15792 4956 15792 4956 0 net604
rlabel metal2 13536 3234 13536 3234 0 net605
rlabel metal2 14592 4158 14592 4158 0 net606
rlabel via6 2152 4426 2152 4426 0 net607
rlabel metal2 15456 4914 15456 4914 0 net608
rlabel metal2 14304 3570 14304 3570 0 net609
rlabel metal3 39984 5712 39984 5712 0 net61
rlabel metal2 14688 3990 14688 3990 0 net610
rlabel metal2 15744 4200 15744 4200 0 net611
rlabel metal2 16800 4998 16800 4998 0 net612
rlabel metal2 15456 3318 15456 3318 0 net613
rlabel metal2 16512 4620 16512 4620 0 net614
rlabel metal2 16224 3948 16224 3948 0 net615
rlabel metal2 16608 3066 16608 3066 0 net616
rlabel metal2 17760 3990 17760 3990 0 net617
rlabel metal4 1248 3360 1248 3360 0 net618
rlabel metal3 21792 4074 21792 4074 0 net619
rlabel metal2 68064 6594 68064 6594 0 net62
rlabel metal2 18528 4410 18528 4410 0 net620
rlabel metal4 25440 3528 25440 3528 0 net621
rlabel metal3 22512 4956 22512 4956 0 net622
rlabel metal4 24000 4620 24000 4620 0 net623
rlabel metal2 20352 4200 20352 4200 0 net624
rlabel metal2 20736 4326 20736 4326 0 net625
rlabel metal3 20064 3402 20064 3402 0 net626
rlabel metal2 20880 3444 20880 3444 0 net627
rlabel metal2 21600 3486 21600 3486 0 net628
rlabel via6 1696 3522 1696 3522 0 net629
rlabel metal2 39168 10206 39168 10206 0 net63
rlabel metal2 23040 4620 23040 4620 0 net630
rlabel metal2 22416 3444 22416 3444 0 net631
rlabel metal2 22752 3528 22752 3528 0 net632
rlabel metal4 23520 5208 23520 5208 0 net633
rlabel metal2 25920 4998 25920 4998 0 net634
rlabel metal2 25344 4410 25344 4410 0 net635
rlabel metal2 24672 3612 24672 3612 0 net636
rlabel metal3 28224 4746 28224 4746 0 net637
rlabel metal2 26112 4074 26112 4074 0 net638
rlabel metal3 26448 3444 26448 3444 0 net639
rlabel metal3 71280 9408 71280 9408 0 net64
rlabel metal5 2152 3486 2152 3486 0 net640
rlabel metal2 27264 5208 27264 5208 0 net641
rlabel metal2 27840 5208 27840 5208 0 net642
rlabel metal2 26208 3402 26208 3402 0 net643
rlabel metal2 26976 4158 26976 4158 0 net644
rlabel metal2 27360 4536 27360 4536 0 net645
rlabel metal3 28080 4116 28080 4116 0 net646
rlabel metal2 27744 3360 27744 3360 0 net647
rlabel metal2 29568 5040 29568 5040 0 net648
rlabel metal2 29856 6216 29856 6216 0 net649
rlabel metal3 37920 6426 37920 6426 0 net65
rlabel metal2 28896 3906 28896 3906 0 net650
rlabel metal4 16416 3528 16416 3528 0 net651
rlabel metal3 30000 3444 30000 3444 0 net652
rlabel metal2 30432 4452 30432 4452 0 net653
rlabel metal2 32256 5208 32256 5208 0 net654
rlabel metal2 31872 4074 31872 4074 0 net655
rlabel metal2 31200 3780 31200 3780 0 net656
rlabel metal3 32352 4956 32352 4956 0 net657
rlabel metal2 31584 4074 31584 4074 0 net658
rlabel metal2 30192 3948 30192 3948 0 net659
rlabel metal2 69120 6426 69120 6426 0 net66
rlabel metal3 32976 4116 32976 4116 0 net660
rlabel metal2 32352 4116 32352 4116 0 net661
rlabel metal3 13734 6300 13734 6300 0 net662
rlabel metal2 33408 4452 33408 4452 0 net663
rlabel metal2 32736 3780 32736 3780 0 net664
rlabel metal2 33504 4368 33504 4368 0 net665
rlabel metal2 34272 3528 34272 3528 0 net666
rlabel metal2 36096 4200 36096 4200 0 net667
rlabel metal3 34704 3444 34704 3444 0 net668
rlabel metal3 37104 4956 37104 4956 0 net669
rlabel metal2 38592 9660 38592 9660 0 net67
rlabel metal2 36864 4788 36864 4788 0 net670
rlabel metal2 36480 3738 36480 3738 0 net671
rlabel metal2 36864 3612 36864 3612 0 net672
rlabel metal2 3168 5040 3168 5040 0 net673
rlabel metal2 82560 10290 82560 10290 0 net68
rlabel metal2 38688 6594 38688 6594 0 net69
rlabel metal3 36096 4872 36096 4872 0 net7
rlabel metal2 68592 7224 68592 7224 0 net70
rlabel metal2 40608 10500 40608 10500 0 net71
rlabel metal2 66144 9240 66144 9240 0 net72
rlabel metal2 39360 6720 39360 6720 0 net73
rlabel metal3 68208 5712 68208 5712 0 net74
rlabel metal3 38640 9408 38640 9408 0 net75
rlabel metal2 72192 9198 72192 9198 0 net76
rlabel metal2 13344 7980 13344 7980 0 net77
rlabel metal2 71040 8652 71040 8652 0 net78
rlabel metal3 38400 8064 38400 8064 0 net79
rlabel metal3 35088 5712 35088 5712 0 net8
rlabel metal2 71136 8064 71136 8064 0 net80
rlabel metal2 19200 8022 19200 8022 0 net81
rlabel metal2 64992 8274 64992 8274 0 net82
rlabel metal2 31104 4242 31104 4242 0 net83
rlabel metal2 67968 4914 67968 4914 0 net84
rlabel metal2 39936 8232 39936 8232 0 net85
rlabel metal2 70752 7980 70752 7980 0 net86
rlabel metal2 18912 7392 18912 7392 0 net87
rlabel metal2 70752 7476 70752 7476 0 net88
rlabel metal2 42336 9576 42336 9576 0 net89
rlabel metal3 36288 8736 36288 8736 0 net9
rlabel metal3 68688 8736 68688 8736 0 net90
rlabel metal3 39744 8442 39744 8442 0 net91
rlabel metal2 70368 7938 70368 7938 0 net92
rlabel metal2 18432 7686 18432 7686 0 net93
rlabel metal2 69792 7728 69792 7728 0 net94
rlabel metal3 71328 7896 71328 7896 0 net95
rlabel metal2 72000 9114 72000 9114 0 net96
rlabel metal2 53760 5838 53760 5838 0 net97
rlabel metal2 54432 6342 54432 6342 0 net98
rlabel metal2 56544 6594 56544 6594 0 net99
rlabel metal2 1056 6216 1056 6216 0 output_no[0]
rlabel metal2 39264 828 39264 828 0 output_no[100]
rlabel metal2 39648 576 39648 576 0 output_no[101]
rlabel metal2 40032 912 40032 912 0 output_no[102]
rlabel metal2 40416 2382 40416 2382 0 output_no[103]
rlabel metal2 40800 660 40800 660 0 output_no[104]
rlabel metal2 41184 1206 41184 1206 0 output_no[105]
rlabel metal2 41568 618 41568 618 0 output_no[106]
rlabel metal2 39744 2394 39744 2394 0 output_no[107]
rlabel metal2 42336 72 42336 72 0 output_no[108]
rlabel metal2 41376 2772 41376 2772 0 output_no[109]
rlabel metal2 4704 828 4704 828 0 output_no[10]
rlabel metal2 40512 1974 40512 1974 0 output_no[110]
rlabel metal2 43488 1500 43488 1500 0 output_no[111]
rlabel metal2 43872 1332 43872 1332 0 output_no[112]
rlabel metal2 41280 1764 41280 1764 0 output_no[113]
rlabel metal2 44640 1710 44640 1710 0 output_no[114]
rlabel metal2 45024 156 45024 156 0 output_no[115]
rlabel metal2 45408 2046 45408 2046 0 output_no[116]
rlabel metal2 45792 2004 45792 2004 0 output_no[117]
rlabel metal2 46176 1920 46176 1920 0 output_no[118]
rlabel metal2 46560 1458 46560 1458 0 output_no[119]
rlabel metal2 5088 1038 5088 1038 0 output_no[11]
rlabel metal2 43968 3066 43968 3066 0 output_no[120]
rlabel metal2 47376 3696 47376 3696 0 output_no[121]
rlabel metal2 47712 576 47712 576 0 output_no[122]
rlabel metal2 48096 660 48096 660 0 output_no[123]
rlabel metal2 48384 3696 48384 3696 0 output_no[124]
rlabel metal2 48672 5460 48672 5460 0 output_no[125]
rlabel metal3 48960 3024 48960 3024 0 output_no[126]
rlabel metal2 49632 1206 49632 1206 0 output_no[127]
rlabel metal2 50016 786 50016 786 0 output_no[128]
rlabel metal2 50448 420 50448 420 0 output_no[129]
rlabel metal2 5472 1038 5472 1038 0 output_no[12]
rlabel metal2 50736 3192 50736 3192 0 output_no[130]
rlabel metal2 51168 1290 51168 1290 0 output_no[131]
rlabel metal2 51552 828 51552 828 0 output_no[132]
rlabel metal2 51936 870 51936 870 0 output_no[133]
rlabel metal2 52320 828 52320 828 0 output_no[134]
rlabel metal2 52704 1038 52704 1038 0 output_no[135]
rlabel metal2 53088 744 53088 744 0 output_no[136]
rlabel metal2 53472 1626 53472 1626 0 output_no[137]
rlabel metal2 53856 702 53856 702 0 output_no[138]
rlabel metal2 54240 828 54240 828 0 output_no[139]
rlabel metal2 5856 996 5856 996 0 output_no[13]
rlabel metal2 54624 1206 54624 1206 0 output_no[140]
rlabel metal2 55008 786 55008 786 0 output_no[141]
rlabel metal2 55392 1164 55392 1164 0 output_no[142]
rlabel metal2 55776 408 55776 408 0 output_no[143]
rlabel metal2 56160 534 56160 534 0 output_no[144]
rlabel metal2 56544 576 56544 576 0 output_no[145]
rlabel metal2 56928 1752 56928 1752 0 output_no[146]
rlabel metal2 57312 1122 57312 1122 0 output_no[147]
rlabel metal3 58272 2688 58272 2688 0 output_no[148]
rlabel metal2 58080 1164 58080 1164 0 output_no[149]
rlabel metal2 6240 1038 6240 1038 0 output_no[14]
rlabel metal2 58464 1122 58464 1122 0 output_no[150]
rlabel metal2 58848 1290 58848 1290 0 output_no[151]
rlabel metal2 59232 576 59232 576 0 output_no[152]
rlabel metal2 59616 1290 59616 1290 0 output_no[153]
rlabel metal2 60000 1290 60000 1290 0 output_no[154]
rlabel metal2 60384 954 60384 954 0 output_no[155]
rlabel metal3 62112 3192 62112 3192 0 output_no[156]
rlabel metal2 61152 1248 61152 1248 0 output_no[157]
rlabel metal2 61536 1290 61536 1290 0 output_no[158]
rlabel metal2 61920 1458 61920 1458 0 output_no[159]
rlabel metal2 6624 1038 6624 1038 0 output_no[15]
rlabel metal2 62304 1206 62304 1206 0 output_no[160]
rlabel metal2 62688 618 62688 618 0 output_no[161]
rlabel metal2 63024 3024 63024 3024 0 output_no[162]
rlabel metal2 63456 1038 63456 1038 0 output_no[163]
rlabel metal2 66144 2982 66144 2982 0 output_no[164]
rlabel metal2 64224 828 64224 828 0 output_no[165]
rlabel metal3 65712 2856 65712 2856 0 output_no[166]
rlabel metal3 66144 2940 66144 2940 0 output_no[167]
rlabel metal3 66528 2604 66528 2604 0 output_no[168]
rlabel metal2 65760 744 65760 744 0 output_no[169]
rlabel metal2 7008 1038 7008 1038 0 output_no[16]
rlabel metal2 66144 1206 66144 1206 0 output_no[170]
rlabel metal3 67680 2772 67680 2772 0 output_no[171]
rlabel metal2 66912 702 66912 702 0 output_no[172]
rlabel metal2 67296 1290 67296 1290 0 output_no[173]
rlabel metal2 67680 450 67680 450 0 output_no[174]
rlabel metal2 68064 828 68064 828 0 output_no[175]
rlabel metal2 68448 1206 68448 1206 0 output_no[176]
rlabel metal3 69984 2604 69984 2604 0 output_no[177]
rlabel metal2 69216 534 69216 534 0 output_no[178]
rlabel metal2 69600 1290 69600 1290 0 output_no[179]
rlabel metal2 7392 996 7392 996 0 output_no[17]
rlabel metal2 69984 492 69984 492 0 output_no[180]
rlabel metal2 70368 282 70368 282 0 output_no[181]
rlabel metal2 70752 534 70752 534 0 output_no[182]
rlabel metal2 71136 828 71136 828 0 output_no[183]
rlabel metal2 71520 450 71520 450 0 output_no[184]
rlabel metal2 71904 576 71904 576 0 output_no[185]
rlabel metal2 72288 408 72288 408 0 output_no[186]
rlabel metal2 72672 198 72672 198 0 output_no[187]
rlabel metal2 73056 618 73056 618 0 output_no[188]
rlabel metal2 73440 1290 73440 1290 0 output_no[189]
rlabel metal2 7776 1038 7776 1038 0 output_no[18]
rlabel metal2 73824 744 73824 744 0 output_no[190]
rlabel metal2 74208 870 74208 870 0 output_no[191]
rlabel metal2 74592 576 74592 576 0 output_no[192]
rlabel metal2 74976 1290 74976 1290 0 output_no[193]
rlabel metal2 75360 1290 75360 1290 0 output_no[194]
rlabel metal2 75744 534 75744 534 0 output_no[195]
rlabel metal2 76128 1290 76128 1290 0 output_no[196]
rlabel metal3 78048 2856 78048 2856 0 output_no[197]
rlabel metal2 76896 660 76896 660 0 output_no[198]
rlabel metal2 77280 786 77280 786 0 output_no[199]
rlabel metal2 8160 1038 8160 1038 0 output_no[19]
rlabel metal2 1248 1416 1248 1416 0 output_no[1]
rlabel metal2 77664 492 77664 492 0 output_no[200]
rlabel metal2 78048 1038 78048 1038 0 output_no[201]
rlabel metal2 78432 1164 78432 1164 0 output_no[202]
rlabel metal2 78816 366 78816 366 0 output_no[203]
rlabel metal2 79200 534 79200 534 0 output_no[204]
rlabel metal2 79584 576 79584 576 0 output_no[205]
rlabel metal2 79968 660 79968 660 0 output_no[206]
rlabel metal2 80352 408 80352 408 0 output_no[207]
rlabel metal2 80736 240 80736 240 0 output_no[208]
rlabel metal2 81120 1626 81120 1626 0 output_no[209]
rlabel metal2 8544 786 8544 786 0 output_no[20]
rlabel metal2 81504 786 81504 786 0 output_no[210]
rlabel metal2 81888 870 81888 870 0 output_no[211]
rlabel metal2 82272 702 82272 702 0 output_no[212]
rlabel metal2 82656 744 82656 744 0 output_no[213]
rlabel metal2 83040 828 83040 828 0 output_no[214]
rlabel metal2 83424 534 83424 534 0 output_no[215]
rlabel metal2 83808 282 83808 282 0 output_no[216]
rlabel metal2 84192 618 84192 618 0 output_no[217]
rlabel metal2 84576 366 84576 366 0 output_no[218]
rlabel metal2 84960 1248 84960 1248 0 output_no[219]
rlabel metal2 8928 1038 8928 1038 0 output_no[21]
rlabel metal2 85344 534 85344 534 0 output_no[220]
rlabel metal2 85728 576 85728 576 0 output_no[221]
rlabel metal2 86112 786 86112 786 0 output_no[222]
rlabel metal2 86496 660 86496 660 0 output_no[223]
rlabel metal2 86880 576 86880 576 0 output_no[224]
rlabel metal2 87264 744 87264 744 0 output_no[225]
rlabel metal2 87648 660 87648 660 0 output_no[226]
rlabel metal2 88032 828 88032 828 0 output_no[227]
rlabel metal2 88416 702 88416 702 0 output_no[228]
rlabel via2 88800 72 88800 72 0 output_no[229]
rlabel metal2 9264 3192 9264 3192 0 output_no[22]
rlabel metal2 89184 660 89184 660 0 output_no[230]
rlabel metal2 89568 576 89568 576 0 output_no[231]
rlabel metal2 89952 660 89952 660 0 output_no[232]
rlabel metal2 90336 702 90336 702 0 output_no[233]
rlabel metal2 90720 240 90720 240 0 output_no[234]
rlabel metal2 91104 828 91104 828 0 output_no[235]
rlabel metal2 91488 744 91488 744 0 output_no[236]
rlabel metal2 91872 702 91872 702 0 output_no[237]
rlabel metal2 92256 786 92256 786 0 output_no[238]
rlabel metal2 92640 828 92640 828 0 output_no[239]
rlabel metal2 9696 534 9696 534 0 output_no[23]
rlabel metal2 93024 744 93024 744 0 output_no[240]
rlabel metal2 93408 702 93408 702 0 output_no[241]
rlabel metal2 93792 786 93792 786 0 output_no[242]
rlabel metal2 94176 828 94176 828 0 output_no[243]
rlabel metal2 94560 1038 94560 1038 0 output_no[244]
rlabel metal2 94944 744 94944 744 0 output_no[245]
rlabel metal2 95328 786 95328 786 0 output_no[246]
rlabel metal3 96048 2856 96048 2856 0 output_no[247]
rlabel metal2 96096 828 96096 828 0 output_no[248]
rlabel metal2 96480 744 96480 744 0 output_no[249]
rlabel metal2 10080 660 10080 660 0 output_no[24]
rlabel metal2 96864 618 96864 618 0 output_no[250]
rlabel metal2 97248 786 97248 786 0 output_no[251]
rlabel metal2 97632 702 97632 702 0 output_no[252]
rlabel metal2 98016 1206 98016 1206 0 output_no[253]
rlabel metal3 98256 3024 98256 3024 0 output_no[254]
rlabel metal2 98784 618 98784 618 0 output_no[255]
rlabel metal2 10464 1038 10464 1038 0 output_no[25]
rlabel metal2 10848 1038 10848 1038 0 output_no[26]
rlabel metal2 11232 1038 11232 1038 0 output_no[27]
rlabel metal2 11616 1290 11616 1290 0 output_no[28]
rlabel metal2 12000 1290 12000 1290 0 output_no[29]
rlabel metal2 1632 1206 1632 1206 0 output_no[2]
rlabel metal2 12384 1290 12384 1290 0 output_no[30]
rlabel metal2 12768 660 12768 660 0 output_no[31]
rlabel metal2 13152 324 13152 324 0 output_no[32]
rlabel metal2 13536 1290 13536 1290 0 output_no[33]
rlabel metal2 13920 282 13920 282 0 output_no[34]
rlabel metal2 14304 1248 14304 1248 0 output_no[35]
rlabel metal2 14688 1290 14688 1290 0 output_no[36]
rlabel metal2 15072 828 15072 828 0 output_no[37]
rlabel metal2 15456 660 15456 660 0 output_no[38]
rlabel metal2 15840 1290 15840 1290 0 output_no[39]
rlabel metal2 2016 1038 2016 1038 0 output_no[3]
rlabel metal2 16224 576 16224 576 0 output_no[40]
rlabel metal2 16608 618 16608 618 0 output_no[41]
rlabel metal2 16992 1248 16992 1248 0 output_no[42]
rlabel metal2 17376 618 17376 618 0 output_no[43]
rlabel metal2 17760 828 17760 828 0 output_no[44]
rlabel metal2 18144 660 18144 660 0 output_no[45]
rlabel metal2 18528 1290 18528 1290 0 output_no[46]
rlabel metal2 18912 198 18912 198 0 output_no[47]
rlabel metal2 19296 1290 19296 1290 0 output_no[48]
rlabel metal3 18432 3192 18432 3192 0 output_no[49]
rlabel metal2 2400 996 2400 996 0 output_no[4]
rlabel metal2 20064 1248 20064 1248 0 output_no[50]
rlabel metal2 20448 1290 20448 1290 0 output_no[51]
rlabel metal4 20832 4242 20832 4242 0 output_no[52]
rlabel metal2 21216 1290 21216 1290 0 output_no[53]
rlabel metal2 19104 2394 19104 2394 0 output_no[54]
rlabel metal2 19488 2352 19488 2352 0 output_no[55]
rlabel metal2 19872 2268 19872 2268 0 output_no[56]
rlabel metal2 22752 1206 22752 1206 0 output_no[57]
rlabel metal2 23136 618 23136 618 0 output_no[58]
rlabel metal2 23520 534 23520 534 0 output_no[59]
rlabel metal2 2496 3234 2496 3234 0 output_no[5]
rlabel metal2 23904 786 23904 786 0 output_no[60]
rlabel metal2 24288 1290 24288 1290 0 output_no[61]
rlabel metal2 24672 660 24672 660 0 output_no[62]
rlabel metal2 25056 828 25056 828 0 output_no[63]
rlabel metal2 25440 702 25440 702 0 output_no[64]
rlabel metal2 25824 786 25824 786 0 output_no[65]
rlabel metal2 26208 1290 26208 1290 0 output_no[66]
rlabel metal2 26592 618 26592 618 0 output_no[67]
rlabel metal3 26112 3192 26112 3192 0 output_no[68]
rlabel metal2 27360 1290 27360 1290 0 output_no[69]
rlabel metal2 3168 618 3168 618 0 output_no[6]
rlabel metal2 27744 1290 27744 1290 0 output_no[70]
rlabel metal2 28128 912 28128 912 0 output_no[71]
rlabel metal3 27792 2688 27792 2688 0 output_no[72]
rlabel metal2 28896 786 28896 786 0 output_no[73]
rlabel metal2 29280 1290 29280 1290 0 output_no[74]
rlabel metal2 29664 1290 29664 1290 0 output_no[75]
rlabel metal2 30048 1206 30048 1206 0 output_no[76]
rlabel metal2 30432 618 30432 618 0 output_no[77]
rlabel metal2 30816 534 30816 534 0 output_no[78]
rlabel metal2 31200 1374 31200 1374 0 output_no[79]
rlabel metal3 3408 3108 3408 3108 0 output_no[7]
rlabel metal2 31584 660 31584 660 0 output_no[80]
rlabel metal2 31968 828 31968 828 0 output_no[81]
rlabel metal2 32352 1038 32352 1038 0 output_no[82]
rlabel metal2 32736 828 32736 828 0 output_no[83]
rlabel metal2 33120 1206 33120 1206 0 output_no[84]
rlabel metal2 33504 660 33504 660 0 output_no[85]
rlabel metal2 33888 1458 33888 1458 0 output_no[86]
rlabel metal2 34272 912 34272 912 0 output_no[87]
rlabel metal3 33408 2940 33408 2940 0 output_no[88]
rlabel metal2 35040 1164 35040 1164 0 output_no[89]
rlabel metal2 3936 1038 3936 1038 0 output_no[8]
rlabel metal2 35424 618 35424 618 0 output_no[90]
rlabel metal2 35808 660 35808 660 0 output_no[91]
rlabel metal2 36192 492 36192 492 0 output_no[92]
rlabel metal2 36576 576 36576 576 0 output_no[93]
rlabel metal3 36960 3150 36960 3150 0 output_no[94]
rlabel metal2 37344 2382 37344 2382 0 output_no[95]
rlabel metal2 37728 1038 37728 1038 0 output_no[96]
rlabel via2 38112 72 38112 72 0 output_no[97]
rlabel metal2 38496 1206 38496 1206 0 output_no[98]
rlabel metal2 38880 1710 38880 1710 0 output_no[99]
rlabel metal2 4320 1038 4320 1038 0 output_no[9]
rlabel metal2 1056 1710 1056 1710 0 output_o[0]
rlabel metal2 39456 2760 39456 2760 0 output_o[100]
rlabel metal2 39840 2172 39840 2172 0 output_o[101]
rlabel metal2 40224 786 40224 786 0 output_o[102]
rlabel metal2 40608 576 40608 576 0 output_o[103]
rlabel metal2 40992 2172 40992 2172 0 output_o[104]
rlabel metal2 41376 324 41376 324 0 output_o[105]
rlabel metal2 41184 3612 41184 3612 0 output_o[106]
rlabel metal2 40512 3654 40512 3654 0 output_o[107]
rlabel metal2 40128 2436 40128 2436 0 output_o[108]
rlabel metal2 42912 1290 42912 1290 0 output_o[109]
rlabel metal2 4896 786 4896 786 0 output_o[10]
rlabel metal2 41280 3864 41280 3864 0 output_o[110]
rlabel metal2 40896 2310 40896 2310 0 output_o[111]
rlabel metal2 44064 1416 44064 1416 0 output_o[112]
rlabel metal2 44448 1710 44448 1710 0 output_o[113]
rlabel metal2 44832 492 44832 492 0 output_o[114]
rlabel metal2 45216 534 45216 534 0 output_o[115]
rlabel metal2 45600 828 45600 828 0 output_o[116]
rlabel metal2 45984 660 45984 660 0 output_o[117]
rlabel metal2 46368 1542 46368 1542 0 output_o[118]
rlabel metal2 46848 3444 46848 3444 0 output_o[119]
rlabel metal2 5280 828 5280 828 0 output_o[11]
rlabel metal2 44352 2982 44352 2982 0 output_o[120]
rlabel metal2 44736 2898 44736 2898 0 output_o[121]
rlabel metal2 47904 618 47904 618 0 output_o[122]
rlabel metal2 45504 2856 45504 2856 0 output_o[123]
rlabel metal2 48672 828 48672 828 0 output_o[124]
rlabel metal3 48624 3528 48624 3528 0 output_o[125]
rlabel metal3 49200 3612 49200 3612 0 output_o[126]
rlabel metal2 49824 828 49824 828 0 output_o[127]
rlabel metal3 49584 3192 49584 3192 0 output_o[128]
rlabel metal2 50592 1038 50592 1038 0 output_o[129]
rlabel metal2 5664 870 5664 870 0 output_o[12]
rlabel metal2 50976 1290 50976 1290 0 output_o[130]
rlabel metal2 51360 1290 51360 1290 0 output_o[131]
rlabel metal2 51744 660 51744 660 0 output_o[132]
rlabel metal2 52128 1206 52128 1206 0 output_o[133]
rlabel metal2 52512 912 52512 912 0 output_o[134]
rlabel metal3 53520 3780 53520 3780 0 output_o[135]
rlabel metal2 53280 660 53280 660 0 output_o[136]
rlabel metal2 53664 1710 53664 1710 0 output_o[137]
rlabel metal2 54048 2004 54048 2004 0 output_o[138]
rlabel metal2 54432 1290 54432 1290 0 output_o[139]
rlabel metal2 6048 912 6048 912 0 output_o[13]
rlabel metal2 54816 450 54816 450 0 output_o[140]
rlabel metal2 55200 870 55200 870 0 output_o[141]
rlabel metal2 55584 156 55584 156 0 output_o[142]
rlabel metal2 55920 4704 55920 4704 0 output_o[143]
rlabel metal2 56304 4704 56304 4704 0 output_o[144]
rlabel metal2 56736 912 56736 912 0 output_o[145]
rlabel metal2 57120 1416 57120 1416 0 output_o[146]
rlabel metal2 57504 828 57504 828 0 output_o[147]
rlabel metal2 57888 744 57888 744 0 output_o[148]
rlabel metal3 58512 3780 58512 3780 0 output_o[149]
rlabel metal2 6432 1038 6432 1038 0 output_o[14]
rlabel metal2 58656 660 58656 660 0 output_o[150]
rlabel metal2 59040 1206 59040 1206 0 output_o[151]
rlabel metal2 59424 1038 59424 1038 0 output_o[152]
rlabel metal2 59808 618 59808 618 0 output_o[153]
rlabel metal2 60192 450 60192 450 0 output_o[154]
rlabel metal2 60576 828 60576 828 0 output_o[155]
rlabel metal2 60960 534 60960 534 0 output_o[156]
rlabel metal2 61344 492 61344 492 0 output_o[157]
rlabel metal2 61728 576 61728 576 0 output_o[158]
rlabel metal2 62112 492 62112 492 0 output_o[159]
rlabel metal2 6816 954 6816 954 0 output_o[15]
rlabel metal3 62784 4536 62784 4536 0 output_o[160]
rlabel metal3 63504 4704 63504 4704 0 output_o[161]
rlabel metal2 63264 870 63264 870 0 output_o[162]
rlabel metal2 63696 3276 63696 3276 0 output_o[163]
rlabel metal2 64032 660 64032 660 0 output_o[164]
rlabel metal2 64416 1038 64416 1038 0 output_o[165]
rlabel metal2 64800 1038 64800 1038 0 output_o[166]
rlabel metal2 65184 1206 65184 1206 0 output_o[167]
rlabel metal2 65568 1206 65568 1206 0 output_o[168]
rlabel metal2 65952 660 65952 660 0 output_o[169]
rlabel metal2 7200 996 7200 996 0 output_o[16]
rlabel metal3 67392 3192 67392 3192 0 output_o[170]
rlabel metal2 66720 1290 66720 1290 0 output_o[171]
rlabel metal2 67104 828 67104 828 0 output_o[172]
rlabel metal2 67488 576 67488 576 0 output_o[173]
rlabel metal2 67872 1206 67872 1206 0 output_o[174]
rlabel metal2 68256 954 68256 954 0 output_o[175]
rlabel metal2 68640 618 68640 618 0 output_o[176]
rlabel metal2 69024 1290 69024 1290 0 output_o[177]
rlabel metal2 69408 660 69408 660 0 output_o[178]
rlabel metal2 69792 1206 69792 1206 0 output_o[179]
rlabel metal2 7584 870 7584 870 0 output_o[17]
rlabel metal2 70176 1290 70176 1290 0 output_o[180]
rlabel metal2 70560 1290 70560 1290 0 output_o[181]
rlabel metal2 70944 1038 70944 1038 0 output_o[182]
rlabel metal2 71328 870 71328 870 0 output_o[183]
rlabel metal2 71712 786 71712 786 0 output_o[184]
rlabel metal2 72096 1374 72096 1374 0 output_o[185]
rlabel metal2 72480 1080 72480 1080 0 output_o[186]
rlabel metal2 72864 912 72864 912 0 output_o[187]
rlabel metal2 73248 660 73248 660 0 output_o[188]
rlabel metal2 73632 492 73632 492 0 output_o[189]
rlabel metal2 7968 1038 7968 1038 0 output_o[18]
rlabel metal2 74016 450 74016 450 0 output_o[190]
rlabel metal3 74832 3024 74832 3024 0 output_o[191]
rlabel metal3 76416 2940 76416 2940 0 output_o[192]
rlabel metal3 76800 2772 76800 2772 0 output_o[193]
rlabel metal2 75552 1248 75552 1248 0 output_o[194]
rlabel metal2 75936 1164 75936 1164 0 output_o[195]
rlabel metal2 76320 618 76320 618 0 output_o[196]
rlabel metal2 76704 1206 76704 1206 0 output_o[197]
rlabel metal2 77088 534 77088 534 0 output_o[198]
rlabel metal2 77472 660 77472 660 0 output_o[199]
rlabel metal2 8352 1122 8352 1122 0 output_o[19]
rlabel metal2 1440 1416 1440 1416 0 output_o[1]
rlabel metal2 77856 408 77856 408 0 output_o[200]
rlabel metal2 78240 1206 78240 1206 0 output_o[201]
rlabel metal2 78624 1122 78624 1122 0 output_o[202]
rlabel metal2 78960 3276 78960 3276 0 output_o[203]
rlabel metal2 79392 114 79392 114 0 output_o[204]
rlabel metal2 79776 366 79776 366 0 output_o[205]
rlabel metal2 80160 618 80160 618 0 output_o[206]
rlabel metal2 80544 660 80544 660 0 output_o[207]
rlabel metal2 80928 744 80928 744 0 output_o[208]
rlabel metal2 81312 534 81312 534 0 output_o[209]
rlabel metal2 8736 828 8736 828 0 output_o[20]
rlabel metal2 81696 1290 81696 1290 0 output_o[210]
rlabel metal2 82080 324 82080 324 0 output_o[211]
rlabel metal2 82464 450 82464 450 0 output_o[212]
rlabel metal2 82848 156 82848 156 0 output_o[213]
rlabel metal2 83232 576 83232 576 0 output_o[214]
rlabel metal2 83616 408 83616 408 0 output_o[215]
rlabel metal2 84000 660 84000 660 0 output_o[216]
rlabel metal2 84384 660 84384 660 0 output_o[217]
rlabel metal2 84768 1290 84768 1290 0 output_o[218]
rlabel metal2 85152 1290 85152 1290 0 output_o[219]
rlabel metal2 9120 1206 9120 1206 0 output_o[21]
rlabel metal2 85536 660 85536 660 0 output_o[220]
rlabel metal2 85920 1206 85920 1206 0 output_o[221]
rlabel metal2 86304 1290 86304 1290 0 output_o[222]
rlabel metal2 86688 702 86688 702 0 output_o[223]
rlabel metal2 87072 1290 87072 1290 0 output_o[224]
rlabel metal3 88320 3192 88320 3192 0 output_o[225]
rlabel metal2 87840 660 87840 660 0 output_o[226]
rlabel metal2 88224 1290 88224 1290 0 output_o[227]
rlabel metal2 88608 996 88608 996 0 output_o[228]
rlabel metal2 88992 786 88992 786 0 output_o[229]
rlabel metal2 9504 1290 9504 1290 0 output_o[22]
rlabel metal2 89376 1206 89376 1206 0 output_o[230]
rlabel metal3 90912 1764 90912 1764 0 output_o[231]
rlabel metal2 90144 828 90144 828 0 output_o[232]
rlabel metal2 90528 786 90528 786 0 output_o[233]
rlabel metal2 90912 870 90912 870 0 output_o[234]
rlabel metal2 91296 912 91296 912 0 output_o[235]
rlabel metal2 91680 828 91680 828 0 output_o[236]
rlabel metal2 92064 786 92064 786 0 output_o[237]
rlabel metal2 92448 870 92448 870 0 output_o[238]
rlabel metal2 92832 912 92832 912 0 output_o[239]
rlabel metal2 9888 618 9888 618 0 output_o[23]
rlabel metal3 93888 3192 93888 3192 0 output_o[240]
rlabel metal2 93600 828 93600 828 0 output_o[241]
rlabel metal2 93984 870 93984 870 0 output_o[242]
rlabel metal2 94368 786 94368 786 0 output_o[243]
rlabel metal2 94752 912 94752 912 0 output_o[244]
rlabel metal2 95136 828 95136 828 0 output_o[245]
rlabel metal2 95520 702 95520 702 0 output_o[246]
rlabel metal2 95904 870 95904 870 0 output_o[247]
rlabel metal2 96288 786 96288 786 0 output_o[248]
rlabel metal2 96672 1290 96672 1290 0 output_o[249]
rlabel metal2 10272 702 10272 702 0 output_o[24]
rlabel metal3 97728 3192 97728 3192 0 output_o[250]
rlabel metal2 97440 1206 97440 1206 0 output_o[251]
rlabel metal2 97824 1206 97824 1206 0 output_o[252]
rlabel metal2 98208 1290 98208 1290 0 output_o[253]
rlabel metal2 98592 1290 98592 1290 0 output_o[254]
rlabel metal3 98400 4284 98400 4284 0 output_o[255]
rlabel metal2 10656 828 10656 828 0 output_o[25]
rlabel metal2 11040 870 11040 870 0 output_o[26]
rlabel metal2 11424 786 11424 786 0 output_o[27]
rlabel metal2 11808 912 11808 912 0 output_o[28]
rlabel metal2 12192 954 12192 954 0 output_o[29]
rlabel metal2 1824 1206 1824 1206 0 output_o[2]
rlabel metal2 12576 870 12576 870 0 output_o[30]
rlabel metal2 12960 996 12960 996 0 output_o[31]
rlabel metal2 13344 1164 13344 1164 0 output_o[32]
rlabel metal2 13728 660 13728 660 0 output_o[33]
rlabel metal2 14112 1290 14112 1290 0 output_o[34]
rlabel metal2 14496 786 14496 786 0 output_o[35]
rlabel metal2 14880 702 14880 702 0 output_o[36]
rlabel metal2 15264 660 15264 660 0 output_o[37]
rlabel metal2 15648 534 15648 534 0 output_o[38]
rlabel metal2 16032 660 16032 660 0 output_o[39]
rlabel metal2 2208 1206 2208 1206 0 output_o[3]
rlabel metal2 16416 1248 16416 1248 0 output_o[40]
rlabel metal2 16800 240 16800 240 0 output_o[41]
rlabel metal2 17184 786 17184 786 0 output_o[42]
rlabel metal2 17568 1248 17568 1248 0 output_o[43]
rlabel metal2 17952 450 17952 450 0 output_o[44]
rlabel metal2 18336 576 18336 576 0 output_o[45]
rlabel metal2 18720 450 18720 450 0 output_o[46]
rlabel metal2 19104 492 19104 492 0 output_o[47]
rlabel metal2 19488 324 19488 324 0 output_o[48]
rlabel metal2 19872 366 19872 366 0 output_o[49]
rlabel metal2 2592 1206 2592 1206 0 output_o[4]
rlabel metal2 18336 2604 18336 2604 0 output_o[50]
rlabel metal2 18768 3360 18768 3360 0 output_o[51]
rlabel metal2 18720 2100 18720 2100 0 output_o[52]
rlabel metal2 21408 660 21408 660 0 output_o[53]
rlabel metal2 21792 1290 21792 1290 0 output_o[54]
rlabel metal2 22176 618 22176 618 0 output_o[55]
rlabel metal2 22560 492 22560 492 0 output_o[56]
rlabel metal2 22944 450 22944 450 0 output_o[57]
rlabel metal2 23328 660 23328 660 0 output_o[58]
rlabel metal2 23712 870 23712 870 0 output_o[59]
rlabel metal2 1824 2856 1824 2856 0 output_o[5]
rlabel metal2 24096 618 24096 618 0 output_o[60]
rlabel metal2 24480 576 24480 576 0 output_o[61]
rlabel metal2 24864 660 24864 660 0 output_o[62]
rlabel metal2 25248 1248 25248 1248 0 output_o[63]
rlabel metal2 25632 1206 25632 1206 0 output_o[64]
rlabel metal2 26016 660 26016 660 0 output_o[65]
rlabel metal2 26400 870 26400 870 0 output_o[66]
rlabel metal2 26784 1290 26784 1290 0 output_o[67]
rlabel metal2 27168 534 27168 534 0 output_o[68]
rlabel metal2 27552 1248 27552 1248 0 output_o[69]
rlabel metal2 3360 1080 3360 1080 0 output_o[6]
rlabel metal2 27936 1290 27936 1290 0 output_o[70]
rlabel metal2 28320 1290 28320 1290 0 output_o[71]
rlabel metal2 28704 954 28704 954 0 output_o[72]
rlabel metal2 29088 702 29088 702 0 output_o[73]
rlabel metal2 29472 828 29472 828 0 output_o[74]
rlabel metal2 29856 660 29856 660 0 output_o[75]
rlabel metal2 30240 576 30240 576 0 output_o[76]
rlabel metal2 30624 492 30624 492 0 output_o[77]
rlabel metal2 31008 576 31008 576 0 output_o[78]
rlabel metal2 31392 534 31392 534 0 output_o[79]
rlabel metal2 3744 702 3744 702 0 output_o[7]
rlabel metal2 31776 702 31776 702 0 output_o[80]
rlabel metal2 32160 828 32160 828 0 output_o[81]
rlabel metal2 32544 1206 32544 1206 0 output_o[82]
rlabel metal2 32928 408 32928 408 0 output_o[83]
rlabel metal2 33312 618 33312 618 0 output_o[84]
rlabel metal2 33696 1206 33696 1206 0 output_o[85]
rlabel metal3 32928 2772 32928 2772 0 output_o[86]
rlabel metal2 34464 1206 34464 1206 0 output_o[87]
rlabel metal2 34848 1038 34848 1038 0 output_o[88]
rlabel metal3 33888 2688 33888 2688 0 output_o[89]
rlabel metal2 4128 660 4128 660 0 output_o[8]
rlabel metal2 35616 1962 35616 1962 0 output_o[90]
rlabel metal2 36000 450 36000 450 0 output_o[91]
rlabel metal2 36384 534 36384 534 0 output_o[92]
rlabel metal2 36768 828 36768 828 0 output_o[93]
rlabel metal2 37152 660 37152 660 0 output_o[94]
rlabel metal2 37536 870 37536 870 0 output_o[95]
rlabel metal2 37920 1290 37920 1290 0 output_o[96]
rlabel metal2 38304 1080 38304 1080 0 output_o[97]
rlabel metal2 38688 744 38688 744 0 output_o[98]
rlabel metal2 39072 618 39072 618 0 output_o[99]
rlabel metal2 4512 618 4512 618 0 output_o[9]
<< properties >>
string FIXED_BBOX 0 0 100000 15000
<< end >>
