magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753774363
<< metal1 >>
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 45763 6656 45821 6657
rect 45763 6616 45772 6656
rect 45812 6616 45821 6656
rect 45763 6615 45821 6616
rect 48547 6656 48605 6657
rect 48547 6616 48556 6656
rect 48596 6616 48605 6656
rect 48547 6615 48605 6616
rect 41739 6488 41781 6497
rect 41739 6448 41740 6488
rect 41780 6448 41781 6488
rect 41739 6439 41781 6448
rect 42027 6488 42069 6497
rect 42027 6448 42028 6488
rect 42068 6448 42069 6488
rect 42027 6439 42069 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44715 6488 44757 6497
rect 44715 6448 44716 6488
rect 44756 6448 44757 6488
rect 44715 6439 44757 6448
rect 45859 6488 45917 6489
rect 45859 6448 45868 6488
rect 45908 6448 45917 6488
rect 45859 6447 45917 6448
rect 46435 6488 46493 6489
rect 46435 6448 46444 6488
rect 46484 6448 46493 6488
rect 46435 6447 46493 6448
rect 46539 6488 46581 6497
rect 46539 6448 46540 6488
rect 46580 6448 46581 6488
rect 46539 6439 46581 6448
rect 47595 6488 47637 6497
rect 47595 6448 47596 6488
rect 47636 6448 47637 6488
rect 47595 6439 47637 6448
rect 47883 6488 47925 6497
rect 47883 6448 47884 6488
rect 47924 6448 47925 6488
rect 47883 6439 47925 6448
rect 48451 6488 48509 6489
rect 48451 6448 48460 6488
rect 48500 6448 48509 6488
rect 48451 6447 48509 6448
rect 48747 6488 48789 6497
rect 48747 6448 48748 6488
rect 48788 6448 48789 6488
rect 48747 6439 48789 6448
rect 49035 6488 49077 6497
rect 49035 6448 49036 6488
rect 49076 6448 49077 6488
rect 49035 6439 49077 6448
rect 49227 6488 49269 6497
rect 49227 6448 49228 6488
rect 49268 6448 49269 6488
rect 49227 6439 49269 6448
rect 49419 6488 49461 6497
rect 49419 6448 49420 6488
rect 49460 6448 49461 6488
rect 49419 6439 49461 6448
rect 46635 6404 46677 6413
rect 46635 6364 46636 6404
rect 46676 6364 46677 6404
rect 46635 6355 46677 6364
rect 48843 6404 48885 6413
rect 48843 6364 48844 6404
rect 48884 6364 48885 6404
rect 48843 6355 48885 6364
rect 49323 6404 49365 6413
rect 49323 6364 49324 6404
rect 49364 6364 49365 6404
rect 49323 6355 49365 6364
rect 41739 6320 41781 6329
rect 41739 6280 41740 6320
rect 41780 6280 41781 6320
rect 41739 6271 41781 6280
rect 46731 6320 46773 6329
rect 46731 6280 46732 6320
rect 46772 6280 46773 6320
rect 46731 6271 46773 6280
rect 46827 6320 46869 6329
rect 46827 6280 46828 6320
rect 46868 6280 46869 6320
rect 46827 6271 46869 6280
rect 47595 6320 47637 6329
rect 47595 6280 47596 6320
rect 47636 6280 47637 6320
rect 47595 6271 47637 6280
rect 48259 6320 48317 6321
rect 48259 6280 48268 6320
rect 48308 6280 48317 6320
rect 48259 6279 48317 6280
rect 44523 6236 44565 6245
rect 44523 6196 44524 6236
rect 44564 6196 44565 6236
rect 44523 6187 44565 6196
rect 46051 6236 46109 6237
rect 46051 6196 46060 6236
rect 46100 6196 46109 6236
rect 46051 6195 46109 6196
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 53451 5900 53493 5909
rect 53451 5860 53452 5900
rect 53492 5860 53493 5900
rect 53451 5851 53493 5860
rect 41067 5648 41109 5657
rect 41067 5608 41068 5648
rect 41108 5608 41109 5648
rect 41067 5599 41109 5608
rect 41355 5648 41397 5657
rect 41355 5608 41356 5648
rect 41396 5608 41397 5648
rect 41355 5599 41397 5608
rect 41739 5648 41781 5657
rect 41739 5608 41740 5648
rect 41780 5608 41781 5648
rect 41739 5599 41781 5608
rect 41835 5648 41877 5657
rect 41835 5608 41836 5648
rect 41876 5608 41877 5648
rect 41835 5599 41877 5608
rect 44235 5648 44277 5657
rect 44235 5608 44236 5648
rect 44276 5608 44277 5648
rect 44235 5599 44277 5608
rect 44331 5648 44373 5657
rect 44331 5608 44332 5648
rect 44372 5608 44373 5648
rect 44331 5599 44373 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45003 5648 45045 5657
rect 45003 5608 45004 5648
rect 45044 5608 45045 5648
rect 45003 5599 45045 5608
rect 46051 5648 46109 5649
rect 46051 5608 46060 5648
rect 46100 5608 46109 5648
rect 46051 5607 46109 5608
rect 46251 5648 46293 5657
rect 46251 5608 46252 5648
rect 46292 5608 46293 5648
rect 46251 5599 46293 5608
rect 46339 5648 46397 5649
rect 46339 5608 46348 5648
rect 46388 5608 46397 5648
rect 46339 5607 46397 5608
rect 50467 5648 50525 5649
rect 50467 5608 50476 5648
rect 50516 5608 50525 5648
rect 50467 5607 50525 5608
rect 50667 5648 50709 5657
rect 50667 5608 50668 5648
rect 50708 5608 50709 5648
rect 50667 5599 50709 5608
rect 51915 5648 51957 5657
rect 51915 5608 51916 5648
rect 51956 5608 51957 5648
rect 51915 5599 51957 5608
rect 52099 5648 52157 5649
rect 52099 5608 52108 5648
rect 52148 5608 52157 5648
rect 52099 5607 52157 5608
rect 52491 5648 52533 5657
rect 52491 5608 52492 5648
rect 52532 5608 52533 5648
rect 52491 5599 52533 5608
rect 52587 5648 52629 5657
rect 52587 5608 52588 5648
rect 52628 5608 52629 5648
rect 52587 5599 52629 5608
rect 53643 5648 53685 5657
rect 53643 5608 53644 5648
rect 53684 5608 53685 5648
rect 53643 5599 53685 5608
rect 53739 5648 53781 5657
rect 53739 5608 53740 5648
rect 53780 5608 53781 5648
rect 53739 5599 53781 5608
rect 54315 5648 54357 5657
rect 54315 5608 54316 5648
rect 54356 5608 54357 5648
rect 54315 5599 54357 5608
rect 54499 5648 54557 5649
rect 54499 5608 54508 5648
rect 54548 5608 54557 5648
rect 54499 5607 54557 5608
rect 55467 5648 55509 5657
rect 55467 5608 55468 5648
rect 55508 5608 55509 5648
rect 55467 5599 55509 5608
rect 55563 5648 55605 5657
rect 55563 5608 55564 5648
rect 55604 5608 55605 5648
rect 55563 5599 55605 5608
rect 56323 5648 56381 5649
rect 56323 5608 56332 5648
rect 56372 5608 56381 5648
rect 56323 5607 56381 5608
rect 56611 5648 56669 5649
rect 56611 5608 56620 5648
rect 56660 5608 56669 5648
rect 56611 5607 56669 5608
rect 56811 5648 56853 5657
rect 56811 5608 56812 5648
rect 56852 5608 56853 5648
rect 56811 5599 56853 5608
rect 58155 5648 58197 5657
rect 58155 5608 58156 5648
rect 58196 5608 58197 5648
rect 58155 5599 58197 5608
rect 58347 5648 58389 5657
rect 58347 5608 58348 5648
rect 58388 5608 58389 5648
rect 58347 5599 58389 5608
rect 61227 5648 61269 5657
rect 61227 5608 61228 5648
rect 61268 5608 61269 5648
rect 61227 5599 61269 5608
rect 61323 5648 61365 5657
rect 61323 5608 61324 5648
rect 61364 5608 61365 5648
rect 61323 5599 61365 5608
rect 61707 5648 61749 5657
rect 61707 5608 61708 5648
rect 61748 5608 61749 5648
rect 61707 5599 61749 5608
rect 61803 5648 61845 5657
rect 61803 5608 61804 5648
rect 61844 5608 61845 5648
rect 61803 5599 61845 5608
rect 61899 5648 61941 5657
rect 61899 5608 61900 5648
rect 61940 5608 61941 5648
rect 61899 5599 61941 5608
rect 61995 5648 62037 5657
rect 61995 5608 61996 5648
rect 62036 5608 62037 5648
rect 61995 5599 62037 5608
rect 41539 5564 41597 5565
rect 41539 5524 41548 5564
rect 41588 5524 41597 5564
rect 41539 5523 41597 5524
rect 44035 5564 44093 5565
rect 44035 5524 44044 5564
rect 44084 5524 44093 5564
rect 44035 5523 44093 5524
rect 44707 5564 44765 5565
rect 44707 5524 44716 5564
rect 44756 5524 44765 5564
rect 44707 5523 44765 5524
rect 50571 5564 50613 5573
rect 50571 5524 50572 5564
rect 50612 5524 50613 5564
rect 50571 5515 50613 5524
rect 52011 5564 52053 5573
rect 52011 5524 52012 5564
rect 52052 5524 52053 5564
rect 52011 5515 52053 5524
rect 52291 5564 52349 5565
rect 52291 5524 52300 5564
rect 52340 5524 52349 5564
rect 52291 5523 52349 5524
rect 54411 5564 54453 5573
rect 54411 5524 54412 5564
rect 54452 5524 54453 5564
rect 54411 5515 54453 5524
rect 55267 5564 55325 5565
rect 55267 5524 55276 5564
rect 55316 5524 55325 5564
rect 55267 5523 55325 5524
rect 56715 5564 56757 5573
rect 56715 5524 56716 5564
rect 56756 5524 56757 5564
rect 56715 5515 56757 5524
rect 61123 5564 61181 5565
rect 61123 5524 61132 5564
rect 61172 5524 61181 5564
rect 61123 5523 61181 5524
rect 41259 5480 41301 5489
rect 41259 5440 41260 5480
rect 41300 5440 41301 5480
rect 41259 5431 41301 5440
rect 41827 5480 41885 5481
rect 41827 5440 41836 5480
rect 41876 5440 41885 5480
rect 41827 5439 41885 5440
rect 44323 5480 44381 5481
rect 44323 5440 44332 5480
rect 44372 5440 44381 5480
rect 44323 5439 44381 5440
rect 44995 5480 45053 5481
rect 44995 5440 45004 5480
rect 45044 5440 45053 5480
rect 44995 5439 45053 5440
rect 46059 5480 46101 5489
rect 46059 5440 46060 5480
rect 46100 5440 46101 5480
rect 46059 5431 46101 5440
rect 52579 5480 52637 5481
rect 52579 5440 52588 5480
rect 52628 5440 52637 5480
rect 52579 5439 52637 5440
rect 53731 5480 53789 5481
rect 53731 5440 53740 5480
rect 53780 5440 53789 5480
rect 53731 5439 53789 5440
rect 55555 5480 55613 5481
rect 55555 5440 55564 5480
rect 55604 5440 55613 5480
rect 55555 5439 55613 5440
rect 56131 5480 56189 5481
rect 56131 5440 56140 5480
rect 56180 5440 56189 5480
rect 56131 5439 56189 5440
rect 56419 5480 56477 5481
rect 56419 5440 56428 5480
rect 56468 5440 56477 5480
rect 56419 5439 56477 5440
rect 58251 5480 58293 5489
rect 58251 5440 58252 5480
rect 58292 5440 58293 5480
rect 58251 5431 58293 5440
rect 60939 5480 60981 5489
rect 60939 5440 60940 5480
rect 60980 5440 60981 5480
rect 60939 5431 60981 5440
rect 61027 5480 61085 5481
rect 61027 5440 61036 5480
rect 61076 5440 61085 5480
rect 61027 5439 61085 5440
rect 61507 5480 61565 5481
rect 61507 5440 61516 5480
rect 61556 5440 61565 5480
rect 61507 5439 61565 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 41443 5144 41501 5145
rect 41443 5104 41452 5144
rect 41492 5104 41501 5144
rect 41443 5103 41501 5104
rect 42115 5144 42173 5145
rect 42115 5104 42124 5144
rect 42164 5104 42173 5144
rect 42115 5103 42173 5104
rect 45859 5144 45917 5145
rect 45859 5104 45868 5144
rect 45908 5104 45917 5144
rect 45859 5103 45917 5104
rect 46627 5144 46685 5145
rect 46627 5104 46636 5144
rect 46676 5104 46685 5144
rect 46627 5103 46685 5104
rect 48067 5144 48125 5145
rect 48067 5104 48076 5144
rect 48116 5104 48125 5144
rect 48067 5103 48125 5104
rect 48835 5144 48893 5145
rect 48835 5104 48844 5144
rect 48884 5104 48893 5144
rect 48835 5103 48893 5104
rect 56611 5144 56669 5145
rect 56611 5104 56620 5144
rect 56660 5104 56669 5144
rect 56611 5103 56669 5104
rect 58051 5144 58109 5145
rect 58051 5104 58060 5144
rect 58100 5104 58109 5144
rect 58051 5103 58109 5104
rect 58723 5144 58781 5145
rect 58723 5104 58732 5144
rect 58772 5104 58781 5144
rect 58723 5103 58781 5104
rect 61891 5144 61949 5145
rect 61891 5104 61900 5144
rect 61940 5104 61949 5144
rect 61891 5103 61949 5104
rect 62179 5060 62237 5061
rect 62179 5020 62188 5060
rect 62228 5020 62237 5060
rect 62179 5019 62237 5020
rect 50859 4987 50901 4996
rect 22435 4976 22493 4977
rect 22435 4936 22444 4976
rect 22484 4936 22493 4976
rect 22435 4935 22493 4936
rect 41355 4976 41397 4985
rect 41355 4936 41356 4976
rect 41396 4936 41397 4976
rect 41355 4927 41397 4936
rect 41451 4976 41493 4985
rect 41451 4936 41452 4976
rect 41492 4936 41493 4976
rect 41451 4927 41493 4936
rect 42027 4976 42069 4985
rect 42027 4936 42028 4976
rect 42068 4936 42069 4976
rect 42027 4927 42069 4936
rect 42123 4976 42165 4985
rect 42123 4936 42124 4976
rect 42164 4936 42165 4976
rect 42123 4927 42165 4936
rect 45867 4976 45909 4985
rect 45867 4936 45868 4976
rect 45908 4936 45909 4976
rect 45867 4927 45909 4936
rect 45963 4976 46005 4985
rect 45963 4936 45964 4976
rect 46004 4936 46005 4976
rect 45963 4927 46005 4936
rect 46539 4976 46581 4985
rect 46539 4936 46540 4976
rect 46580 4936 46581 4976
rect 46539 4927 46581 4936
rect 46635 4976 46677 4985
rect 46635 4936 46636 4976
rect 46676 4936 46677 4976
rect 46635 4927 46677 4936
rect 48075 4976 48117 4985
rect 48075 4936 48076 4976
rect 48116 4936 48117 4976
rect 48075 4927 48117 4936
rect 48171 4976 48213 4985
rect 48171 4936 48172 4976
rect 48212 4936 48213 4976
rect 48171 4927 48213 4936
rect 48747 4976 48789 4985
rect 48747 4936 48748 4976
rect 48788 4936 48789 4976
rect 48747 4927 48789 4936
rect 48843 4976 48885 4985
rect 48843 4936 48844 4976
rect 48884 4936 48885 4976
rect 48843 4927 48885 4936
rect 49315 4976 49373 4977
rect 49315 4936 49324 4976
rect 49364 4936 49373 4976
rect 49315 4935 49373 4936
rect 49515 4976 49557 4985
rect 49515 4936 49516 4976
rect 49556 4936 49557 4976
rect 49515 4927 49557 4936
rect 49603 4976 49661 4977
rect 49603 4936 49612 4976
rect 49652 4936 49661 4976
rect 49603 4935 49661 4936
rect 50379 4976 50421 4985
rect 50379 4936 50380 4976
rect 50420 4936 50421 4976
rect 50379 4927 50421 4936
rect 50667 4976 50709 4985
rect 50667 4936 50668 4976
rect 50708 4936 50709 4976
rect 50859 4947 50860 4987
rect 50900 4947 50901 4987
rect 52676 4987 52734 4988
rect 50859 4938 50901 4947
rect 52395 4976 52437 4985
rect 50667 4927 50709 4936
rect 52395 4936 52396 4976
rect 52436 4936 52437 4976
rect 52676 4947 52685 4987
rect 52725 4947 52734 4987
rect 52676 4946 52734 4947
rect 52875 4976 52917 4985
rect 52395 4927 52437 4936
rect 52875 4936 52876 4976
rect 52916 4936 52917 4976
rect 52875 4927 52917 4936
rect 53539 4976 53597 4977
rect 53539 4936 53548 4976
rect 53588 4936 53597 4976
rect 53539 4935 53597 4936
rect 53739 4976 53781 4985
rect 53739 4936 53740 4976
rect 53780 4936 53781 4976
rect 53739 4927 53781 4936
rect 54891 4976 54933 4985
rect 54891 4936 54892 4976
rect 54932 4936 54933 4976
rect 54891 4927 54933 4936
rect 55179 4976 55221 4985
rect 55179 4936 55180 4976
rect 55220 4936 55221 4976
rect 55179 4927 55221 4936
rect 55371 4976 55413 4985
rect 55371 4936 55372 4976
rect 55412 4936 55413 4976
rect 55371 4927 55413 4936
rect 55947 4976 55989 4985
rect 55947 4936 55948 4976
rect 55988 4936 55989 4976
rect 55947 4927 55989 4936
rect 56139 4976 56181 4985
rect 56139 4936 56140 4976
rect 56180 4936 56181 4976
rect 56139 4927 56181 4936
rect 56331 4976 56373 4985
rect 56331 4936 56332 4976
rect 56372 4936 56373 4976
rect 56331 4927 56373 4936
rect 56427 4976 56469 4985
rect 56427 4936 56428 4976
rect 56468 4936 56469 4976
rect 56427 4927 56469 4936
rect 57963 4976 58005 4985
rect 57963 4936 57964 4976
rect 58004 4936 58005 4976
rect 57963 4927 58005 4936
rect 58059 4976 58101 4985
rect 58059 4936 58060 4976
rect 58100 4936 58101 4976
rect 58059 4927 58101 4936
rect 58635 4976 58677 4985
rect 58635 4936 58636 4976
rect 58676 4936 58677 4976
rect 58635 4927 58677 4936
rect 58731 4976 58773 4985
rect 58731 4936 58732 4976
rect 58772 4936 58773 4976
rect 58731 4927 58773 4936
rect 60459 4976 60501 4985
rect 60459 4936 60460 4976
rect 60500 4936 60501 4976
rect 60459 4927 60501 4936
rect 60843 4976 60885 4985
rect 60843 4936 60844 4976
rect 60884 4936 60885 4976
rect 60843 4927 60885 4936
rect 61035 4976 61077 4985
rect 61035 4936 61036 4976
rect 61076 4936 61077 4976
rect 61035 4927 61077 4936
rect 61219 4976 61277 4977
rect 61219 4936 61228 4976
rect 61268 4936 61277 4976
rect 61219 4935 61277 4936
rect 61323 4976 61365 4985
rect 61323 4936 61324 4976
rect 61364 4936 61365 4976
rect 61323 4927 61365 4936
rect 61507 4976 61565 4977
rect 61507 4936 61516 4976
rect 61556 4936 61565 4976
rect 61507 4935 61565 4936
rect 61899 4976 61941 4985
rect 61899 4936 61900 4976
rect 61940 4936 61941 4976
rect 61899 4927 61941 4936
rect 61995 4976 62037 4985
rect 61995 4936 61996 4976
rect 62036 4936 62037 4976
rect 61995 4927 62037 4936
rect 62371 4976 62429 4977
rect 62371 4936 62380 4976
rect 62420 4936 62429 4976
rect 62371 4935 62429 4936
rect 62571 4976 62613 4985
rect 62571 4936 62572 4976
rect 62612 4936 62613 4976
rect 62571 4927 62613 4936
rect 62659 4976 62717 4977
rect 62659 4936 62668 4976
rect 62708 4936 62717 4976
rect 62659 4935 62717 4936
rect 66891 4976 66933 4985
rect 66891 4936 66892 4976
rect 66932 4936 66933 4976
rect 66891 4927 66933 4936
rect 67179 4976 67221 4985
rect 67179 4936 67180 4976
rect 67220 4936 67221 4976
rect 67179 4927 67221 4936
rect 73323 4976 73365 4985
rect 73323 4936 73324 4976
rect 73364 4936 73365 4976
rect 73323 4927 73365 4936
rect 73611 4976 73653 4985
rect 73611 4936 73612 4976
rect 73652 4936 73653 4976
rect 73611 4927 73653 4936
rect 73803 4976 73845 4985
rect 73803 4936 73804 4976
rect 73844 4936 73845 4976
rect 73803 4927 73845 4936
rect 74091 4976 74133 4985
rect 74091 4936 74092 4976
rect 74132 4936 74133 4976
rect 74091 4927 74133 4936
rect 74283 4976 74325 4985
rect 74283 4936 74284 4976
rect 74324 4936 74325 4976
rect 74283 4927 74325 4936
rect 74475 4976 74517 4985
rect 74475 4936 74476 4976
rect 74516 4936 74517 4976
rect 74475 4927 74517 4936
rect 82155 4976 82197 4985
rect 82155 4936 82156 4976
rect 82196 4936 82197 4976
rect 82155 4927 82197 4936
rect 82347 4976 82389 4985
rect 82347 4936 82348 4976
rect 82388 4936 82389 4976
rect 82347 4927 82389 4936
rect 50763 4892 50805 4901
rect 50763 4852 50764 4892
rect 50804 4852 50805 4892
rect 50763 4843 50805 4852
rect 56043 4892 56085 4901
rect 56043 4852 56044 4892
rect 56084 4852 56085 4892
rect 56043 4843 56085 4852
rect 74379 4892 74421 4901
rect 74379 4852 74380 4892
rect 74420 4852 74421 4892
rect 74379 4843 74421 4852
rect 48555 4808 48597 4817
rect 48555 4768 48556 4808
rect 48596 4768 48597 4808
rect 48555 4759 48597 4768
rect 50379 4808 50421 4817
rect 50379 4768 50380 4808
rect 50420 4768 50421 4808
rect 50379 4759 50421 4768
rect 52395 4808 52437 4817
rect 52395 4768 52396 4808
rect 52436 4768 52437 4808
rect 52395 4759 52437 4768
rect 54891 4808 54933 4817
rect 54891 4768 54892 4808
rect 54932 4768 54933 4808
rect 54891 4759 54933 4768
rect 60459 4808 60501 4817
rect 60459 4768 60460 4808
rect 60500 4768 60501 4808
rect 60459 4759 60501 4768
rect 22347 4724 22389 4733
rect 22347 4684 22348 4724
rect 22388 4684 22389 4724
rect 22347 4675 22389 4684
rect 41163 4724 41205 4733
rect 41163 4684 41164 4724
rect 41204 4684 41205 4724
rect 41163 4675 41205 4684
rect 41835 4724 41877 4733
rect 41835 4684 41836 4724
rect 41876 4684 41877 4724
rect 41835 4675 41877 4684
rect 46155 4724 46197 4733
rect 46155 4684 46156 4724
rect 46196 4684 46197 4724
rect 46155 4675 46197 4684
rect 46347 4724 46389 4733
rect 46347 4684 46348 4724
rect 46388 4684 46389 4724
rect 46347 4675 46389 4684
rect 48363 4724 48405 4733
rect 48363 4684 48364 4724
rect 48404 4684 48405 4724
rect 48363 4675 48405 4684
rect 49515 4724 49557 4733
rect 49515 4684 49516 4724
rect 49556 4684 49557 4724
rect 49515 4675 49557 4684
rect 50187 4724 50229 4733
rect 50187 4684 50188 4724
rect 50228 4684 50229 4724
rect 50187 4675 50229 4684
rect 52203 4724 52245 4733
rect 52203 4684 52204 4724
rect 52244 4684 52245 4724
rect 52203 4675 52245 4684
rect 52683 4724 52725 4733
rect 52683 4684 52684 4724
rect 52724 4684 52725 4724
rect 52683 4675 52725 4684
rect 53643 4724 53685 4733
rect 53643 4684 53644 4724
rect 53684 4684 53685 4724
rect 53643 4675 53685 4684
rect 54699 4724 54741 4733
rect 54699 4684 54700 4724
rect 54740 4684 54741 4724
rect 54699 4675 54741 4684
rect 55179 4724 55221 4733
rect 55179 4684 55180 4724
rect 55220 4684 55221 4724
rect 55179 4675 55221 4684
rect 57771 4724 57813 4733
rect 57771 4684 57772 4724
rect 57812 4684 57813 4724
rect 57771 4675 57813 4684
rect 58443 4724 58485 4733
rect 58443 4684 58444 4724
rect 58484 4684 58485 4724
rect 58443 4675 58485 4684
rect 60651 4724 60693 4733
rect 60651 4684 60652 4724
rect 60692 4684 60693 4724
rect 60651 4675 60693 4684
rect 60843 4724 60885 4733
rect 60843 4684 60844 4724
rect 60884 4684 60885 4724
rect 60843 4675 60885 4684
rect 61323 4724 61365 4733
rect 61323 4684 61324 4724
rect 61364 4684 61365 4724
rect 61323 4675 61365 4684
rect 62379 4724 62421 4733
rect 62379 4684 62380 4724
rect 62420 4684 62421 4724
rect 62379 4675 62421 4684
rect 67179 4724 67221 4733
rect 67179 4684 67180 4724
rect 67220 4684 67221 4724
rect 67179 4675 67221 4684
rect 73323 4724 73365 4733
rect 73323 4684 73324 4724
rect 73364 4684 73365 4724
rect 73323 4675 73365 4684
rect 74091 4724 74133 4733
rect 74091 4684 74092 4724
rect 74132 4684 74133 4724
rect 74091 4675 74133 4684
rect 82155 4724 82197 4733
rect 82155 4684 82156 4724
rect 82196 4684 82197 4724
rect 82155 4675 82197 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 38667 4388 38709 4397
rect 38667 4348 38668 4388
rect 38708 4348 38709 4388
rect 38667 4339 38709 4348
rect 43083 4388 43125 4397
rect 43083 4348 43084 4388
rect 43124 4348 43125 4388
rect 43083 4339 43125 4348
rect 52299 4388 52341 4397
rect 52299 4348 52300 4388
rect 52340 4348 52341 4388
rect 52299 4339 52341 4348
rect 7563 4304 7605 4313
rect 7563 4264 7564 4304
rect 7604 4264 7605 4304
rect 7563 4255 7605 4264
rect 53355 4304 53397 4313
rect 53355 4264 53356 4304
rect 53396 4264 53397 4304
rect 53355 4255 53397 4264
rect 58155 4304 58197 4313
rect 58155 4264 58156 4304
rect 58196 4264 58197 4304
rect 58155 4255 58197 4264
rect 59019 4304 59061 4313
rect 59019 4264 59020 4304
rect 59060 4264 59061 4304
rect 59019 4255 59061 4264
rect 41539 4178 41597 4179
rect 19083 4167 19125 4176
rect 6987 4136 7029 4145
rect 6987 4096 6988 4136
rect 7028 4096 7029 4136
rect 6987 4087 7029 4096
rect 7179 4136 7221 4145
rect 7179 4096 7180 4136
rect 7220 4096 7221 4136
rect 7179 4087 7221 4096
rect 7563 4136 7605 4145
rect 7563 4096 7564 4136
rect 7604 4096 7605 4136
rect 7563 4087 7605 4096
rect 18315 4136 18357 4145
rect 18315 4096 18316 4136
rect 18356 4096 18357 4136
rect 18315 4087 18357 4096
rect 18411 4136 18453 4145
rect 18411 4096 18412 4136
rect 18452 4096 18453 4136
rect 18411 4087 18453 4096
rect 18987 4136 19029 4145
rect 18987 4096 18988 4136
rect 19028 4096 19029 4136
rect 19083 4127 19084 4167
rect 19124 4127 19125 4167
rect 19083 4118 19125 4127
rect 19459 4136 19517 4137
rect 18987 4087 19029 4096
rect 19459 4096 19468 4136
rect 19508 4096 19517 4136
rect 19459 4095 19517 4096
rect 19659 4136 19701 4145
rect 19659 4096 19660 4136
rect 19700 4096 19701 4136
rect 19659 4087 19701 4096
rect 19747 4136 19805 4137
rect 19747 4096 19756 4136
rect 19796 4096 19805 4136
rect 19747 4095 19805 4096
rect 24363 4136 24405 4145
rect 24363 4096 24364 4136
rect 24404 4096 24405 4136
rect 24363 4087 24405 4096
rect 24459 4136 24501 4145
rect 24459 4096 24460 4136
rect 24500 4096 24501 4136
rect 24459 4087 24501 4096
rect 24835 4136 24893 4137
rect 24835 4096 24844 4136
rect 24884 4096 24893 4136
rect 24835 4095 24893 4096
rect 25035 4136 25077 4145
rect 25035 4096 25036 4136
rect 25076 4096 25077 4136
rect 25035 4087 25077 4096
rect 25123 4136 25181 4137
rect 25123 4096 25132 4136
rect 25172 4096 25181 4136
rect 25123 4095 25181 4096
rect 25899 4136 25941 4145
rect 25899 4096 25900 4136
rect 25940 4096 25941 4136
rect 25899 4087 25941 4096
rect 26091 4136 26133 4145
rect 26091 4096 26092 4136
rect 26132 4096 26133 4136
rect 26091 4087 26133 4096
rect 27915 4136 27957 4145
rect 27915 4096 27916 4136
rect 27956 4096 27957 4136
rect 27915 4087 27957 4096
rect 28011 4136 28053 4145
rect 28011 4096 28012 4136
rect 28052 4096 28053 4136
rect 28011 4087 28053 4096
rect 32139 4136 32181 4145
rect 32139 4096 32140 4136
rect 32180 4096 32181 4136
rect 32139 4087 32181 4096
rect 32235 4136 32277 4145
rect 32235 4096 32236 4136
rect 32276 4096 32277 4136
rect 32235 4087 32277 4096
rect 32611 4136 32669 4137
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32611 4095 32669 4096
rect 32811 4136 32853 4145
rect 32811 4096 32812 4136
rect 32852 4096 32853 4136
rect 32811 4087 32853 4096
rect 32899 4136 32957 4137
rect 32899 4096 32908 4136
rect 32948 4096 32957 4136
rect 32899 4095 32957 4096
rect 37227 4136 37269 4145
rect 37227 4096 37228 4136
rect 37268 4096 37269 4136
rect 37227 4087 37269 4096
rect 37323 4136 37365 4145
rect 37323 4096 37324 4136
rect 37364 4096 37365 4136
rect 37323 4087 37365 4096
rect 37699 4136 37757 4137
rect 37699 4096 37708 4136
rect 37748 4096 37757 4136
rect 37699 4095 37757 4096
rect 37803 4136 37845 4145
rect 37803 4096 37804 4136
rect 37844 4096 37845 4136
rect 37803 4087 37845 4096
rect 37987 4136 38045 4137
rect 37987 4096 37996 4136
rect 38036 4096 38045 4136
rect 37987 4095 38045 4096
rect 38379 4136 38421 4145
rect 38379 4096 38380 4136
rect 38420 4096 38421 4136
rect 38379 4087 38421 4096
rect 38475 4136 38517 4145
rect 38475 4096 38476 4136
rect 38516 4096 38517 4136
rect 38475 4087 38517 4096
rect 41251 4136 41309 4137
rect 41251 4096 41260 4136
rect 41300 4096 41309 4136
rect 41251 4095 41309 4096
rect 41451 4136 41493 4145
rect 41539 4138 41548 4178
rect 41588 4138 41597 4178
rect 44611 4178 44669 4179
rect 41539 4137 41597 4138
rect 41451 4096 41452 4136
rect 41492 4096 41493 4136
rect 41451 4087 41493 4096
rect 41931 4136 41973 4145
rect 41931 4096 41932 4136
rect 41972 4096 41973 4136
rect 41931 4087 41973 4096
rect 42027 4136 42069 4145
rect 42027 4096 42028 4136
rect 42068 4096 42069 4136
rect 42027 4087 42069 4096
rect 42403 4136 42461 4137
rect 42403 4096 42412 4136
rect 42452 4096 42461 4136
rect 42403 4095 42461 4096
rect 42603 4136 42645 4145
rect 42603 4096 42604 4136
rect 42644 4096 42645 4136
rect 42603 4087 42645 4096
rect 42691 4136 42749 4137
rect 42691 4096 42700 4136
rect 42740 4096 42749 4136
rect 42691 4095 42749 4096
rect 42883 4136 42941 4137
rect 42883 4096 42892 4136
rect 42932 4096 42941 4136
rect 42883 4095 42941 4096
rect 43083 4136 43125 4145
rect 43083 4096 43084 4136
rect 43124 4096 43125 4136
rect 43083 4087 43125 4096
rect 43171 4136 43229 4137
rect 43171 4096 43180 4136
rect 43220 4096 43229 4136
rect 43171 4095 43229 4096
rect 44323 4136 44381 4137
rect 44323 4096 44332 4136
rect 44372 4096 44381 4136
rect 44323 4095 44381 4096
rect 44523 4136 44565 4145
rect 44611 4138 44620 4178
rect 44660 4138 44669 4178
rect 52395 4151 52437 4160
rect 44611 4137 44669 4138
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44803 4136 44861 4137
rect 44803 4096 44812 4136
rect 44852 4096 44861 4136
rect 44803 4095 44861 4096
rect 45003 4136 45045 4145
rect 45003 4096 45004 4136
rect 45044 4096 45045 4136
rect 45003 4087 45045 4096
rect 45091 4136 45149 4137
rect 45091 4096 45100 4136
rect 45140 4096 45149 4136
rect 45091 4095 45149 4096
rect 46051 4136 46109 4137
rect 46051 4096 46060 4136
rect 46100 4096 46109 4136
rect 46051 4095 46109 4096
rect 46251 4136 46293 4145
rect 46251 4096 46252 4136
rect 46292 4096 46293 4136
rect 46251 4087 46293 4096
rect 46339 4136 46397 4137
rect 46339 4096 46348 4136
rect 46388 4096 46397 4136
rect 46339 4095 46397 4096
rect 48163 4136 48221 4137
rect 48163 4096 48172 4136
rect 48212 4096 48221 4136
rect 48163 4095 48221 4096
rect 48363 4136 48405 4145
rect 48363 4096 48364 4136
rect 48404 4096 48405 4136
rect 48363 4087 48405 4096
rect 48451 4136 48509 4137
rect 48451 4096 48460 4136
rect 48500 4096 48509 4136
rect 48451 4095 48509 4096
rect 48643 4136 48701 4137
rect 48643 4096 48652 4136
rect 48692 4096 48701 4136
rect 48643 4095 48701 4096
rect 48843 4136 48885 4145
rect 48843 4096 48844 4136
rect 48884 4096 48885 4136
rect 48843 4087 48885 4096
rect 48931 4136 48989 4137
rect 48931 4096 48940 4136
rect 48980 4096 48989 4136
rect 48931 4095 48989 4096
rect 50187 4136 50229 4145
rect 50187 4096 50188 4136
rect 50228 4096 50229 4136
rect 50187 4087 50229 4096
rect 50371 4136 50429 4137
rect 50371 4096 50380 4136
rect 50420 4096 50429 4136
rect 50371 4095 50429 4096
rect 50563 4136 50621 4137
rect 50563 4096 50572 4136
rect 50612 4096 50621 4136
rect 50563 4095 50621 4096
rect 50763 4136 50805 4145
rect 50763 4096 50764 4136
rect 50804 4096 50805 4136
rect 50763 4087 50805 4096
rect 51235 4136 51293 4137
rect 51235 4096 51244 4136
rect 51284 4096 51293 4136
rect 51235 4095 51293 4096
rect 51435 4136 51477 4145
rect 51435 4096 51436 4136
rect 51476 4096 51477 4136
rect 51435 4087 51477 4096
rect 51523 4136 51581 4137
rect 51523 4096 51532 4136
rect 51572 4096 51581 4136
rect 51523 4095 51581 4096
rect 52195 4136 52253 4137
rect 52195 4096 52204 4136
rect 52244 4096 52253 4136
rect 52395 4111 52396 4151
rect 52436 4111 52437 4151
rect 52395 4102 52437 4111
rect 52587 4151 52629 4160
rect 52587 4111 52588 4151
rect 52628 4111 52629 4151
rect 52587 4102 52629 4111
rect 52771 4136 52829 4137
rect 52195 4095 52253 4096
rect 52771 4096 52780 4136
rect 52820 4096 52829 4136
rect 52771 4095 52829 4096
rect 53355 4136 53397 4145
rect 53355 4096 53356 4136
rect 53396 4096 53397 4136
rect 53355 4087 53397 4096
rect 53643 4136 53685 4145
rect 53643 4096 53644 4136
rect 53684 4096 53685 4136
rect 53643 4087 53685 4096
rect 53835 4136 53877 4145
rect 53835 4096 53836 4136
rect 53876 4096 53877 4136
rect 53835 4087 53877 4096
rect 55075 4136 55133 4137
rect 55075 4096 55084 4136
rect 55124 4096 55133 4136
rect 55075 4095 55133 4096
rect 55275 4136 55317 4145
rect 55275 4096 55276 4136
rect 55316 4096 55317 4136
rect 55275 4087 55317 4096
rect 55363 4136 55421 4137
rect 55363 4096 55372 4136
rect 55412 4096 55421 4136
rect 55363 4095 55421 4096
rect 58155 4136 58197 4145
rect 58155 4096 58156 4136
rect 58196 4096 58197 4136
rect 58155 4087 58197 4096
rect 58531 4136 58589 4137
rect 58531 4096 58540 4136
rect 58580 4096 58589 4136
rect 58531 4095 58589 4096
rect 58731 4136 58773 4145
rect 58731 4096 58732 4136
rect 58772 4096 58773 4136
rect 58731 4087 58773 4096
rect 59019 4136 59061 4145
rect 59019 4096 59020 4136
rect 59060 4096 59061 4136
rect 59019 4087 59061 4096
rect 59403 4136 59445 4145
rect 59403 4096 59404 4136
rect 59444 4096 59445 4136
rect 59403 4087 59445 4096
rect 59595 4136 59637 4145
rect 59595 4096 59596 4136
rect 59636 4096 59637 4136
rect 59595 4087 59637 4096
rect 61507 4136 61565 4137
rect 61507 4096 61516 4136
rect 61556 4096 61565 4136
rect 61507 4095 61565 4096
rect 61891 4136 61949 4137
rect 61891 4096 61900 4136
rect 61940 4096 61949 4136
rect 61891 4095 61949 4096
rect 62275 4136 62333 4137
rect 62275 4096 62284 4136
rect 62324 4096 62333 4136
rect 62275 4095 62333 4096
rect 62475 4136 62517 4145
rect 62475 4096 62476 4136
rect 62516 4096 62517 4136
rect 62475 4087 62517 4096
rect 66499 4136 66557 4137
rect 66499 4096 66508 4136
rect 66548 4096 66557 4136
rect 66499 4095 66557 4096
rect 66787 4136 66845 4137
rect 66787 4096 66796 4136
rect 66836 4096 66845 4136
rect 66787 4095 66845 4096
rect 66987 4136 67029 4145
rect 66987 4096 66988 4136
rect 67028 4096 67029 4136
rect 66987 4087 67029 4096
rect 68515 4136 68573 4137
rect 68515 4096 68524 4136
rect 68564 4096 68573 4136
rect 68515 4095 68573 4096
rect 68899 4136 68957 4137
rect 68899 4096 68908 4136
rect 68948 4096 68957 4136
rect 68899 4095 68957 4096
rect 69099 4136 69141 4145
rect 69099 4096 69100 4136
rect 69140 4096 69141 4136
rect 69099 4087 69141 4096
rect 74083 4136 74141 4137
rect 74083 4096 74092 4136
rect 74132 4096 74141 4136
rect 74083 4095 74141 4096
rect 74283 4136 74325 4145
rect 74283 4096 74284 4136
rect 74324 4096 74325 4136
rect 74283 4087 74325 4096
rect 74371 4136 74429 4137
rect 74371 4096 74380 4136
rect 74420 4096 74429 4136
rect 74371 4095 74429 4096
rect 74763 4136 74805 4145
rect 74763 4096 74764 4136
rect 74804 4096 74805 4136
rect 74763 4087 74805 4096
rect 74859 4136 74901 4145
rect 74859 4096 74860 4136
rect 74900 4096 74901 4136
rect 74859 4087 74901 4096
rect 80331 4136 80373 4145
rect 80331 4096 80332 4136
rect 80372 4096 80373 4136
rect 80331 4087 80373 4096
rect 80515 4136 80573 4137
rect 80515 4096 80524 4136
rect 80564 4096 80573 4136
rect 80515 4095 80573 4096
rect 80803 4136 80861 4137
rect 80803 4096 80812 4136
rect 80852 4096 80861 4136
rect 80803 4095 80861 4096
rect 86659 4136 86717 4137
rect 86659 4096 86668 4136
rect 86708 4096 86717 4136
rect 86659 4095 86717 4096
rect 87043 4136 87101 4137
rect 87043 4096 87052 4136
rect 87092 4096 87101 4136
rect 87043 4095 87101 4096
rect 87243 4136 87285 4145
rect 87243 4096 87244 4136
rect 87284 4096 87285 4136
rect 87243 4087 87285 4096
rect 91563 4136 91605 4145
rect 91563 4096 91564 4136
rect 91604 4096 91605 4136
rect 91563 4087 91605 4096
rect 91747 4136 91805 4137
rect 91747 4096 91756 4136
rect 91796 4096 91805 4136
rect 91747 4095 91805 4096
rect 92035 4136 92093 4137
rect 92035 4096 92044 4136
rect 92084 4096 92093 4136
rect 92035 4095 92093 4096
rect 18115 4052 18173 4053
rect 18115 4012 18124 4052
rect 18164 4012 18173 4052
rect 18115 4011 18173 4012
rect 18787 4052 18845 4053
rect 18787 4012 18796 4052
rect 18836 4012 18845 4052
rect 18787 4011 18845 4012
rect 24643 4052 24701 4053
rect 24643 4012 24652 4052
rect 24692 4012 24701 4052
rect 24643 4011 24701 4012
rect 31939 4052 31997 4053
rect 31939 4012 31948 4052
rect 31988 4012 31997 4052
rect 31939 4011 31997 4012
rect 37507 4052 37565 4053
rect 37507 4012 37516 4052
rect 37556 4012 37565 4052
rect 37507 4011 37565 4012
rect 41731 4052 41789 4053
rect 41731 4012 41740 4052
rect 41780 4012 41789 4052
rect 41731 4011 41789 4012
rect 50283 4052 50325 4061
rect 50283 4012 50284 4052
rect 50324 4012 50325 4052
rect 50283 4003 50325 4012
rect 50667 4052 50709 4061
rect 50667 4012 50668 4052
rect 50708 4012 50709 4052
rect 50667 4003 50709 4012
rect 52683 4052 52725 4061
rect 52683 4012 52684 4052
rect 52724 4012 52725 4052
rect 52683 4003 52725 4012
rect 58635 4052 58677 4061
rect 58635 4012 58636 4052
rect 58676 4012 58677 4052
rect 58635 4003 58677 4012
rect 62379 4052 62421 4061
rect 62379 4012 62380 4052
rect 62420 4012 62421 4052
rect 62379 4003 62421 4012
rect 66891 4052 66933 4061
rect 66891 4012 66892 4052
rect 66932 4012 66933 4052
rect 66891 4003 66933 4012
rect 69003 4052 69045 4061
rect 69003 4012 69004 4052
rect 69044 4012 69045 4052
rect 69003 4003 69045 4012
rect 75043 4052 75101 4053
rect 75043 4012 75052 4052
rect 75092 4012 75101 4052
rect 75043 4011 75101 4012
rect 80427 4052 80469 4061
rect 80427 4012 80428 4052
rect 80468 4012 80469 4052
rect 80427 4003 80469 4012
rect 87147 4052 87189 4061
rect 87147 4012 87148 4052
rect 87188 4012 87189 4052
rect 87147 4003 87189 4012
rect 91659 4052 91701 4061
rect 91659 4012 91660 4052
rect 91700 4012 91701 4052
rect 91659 4003 91701 4012
rect 7083 3968 7125 3977
rect 7083 3928 7084 3968
rect 7124 3928 7125 3968
rect 7083 3919 7125 3928
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 18403 3968 18461 3969
rect 18403 3928 18412 3968
rect 18452 3928 18461 3968
rect 18403 3927 18461 3928
rect 19075 3968 19133 3969
rect 19075 3928 19084 3968
rect 19124 3928 19133 3968
rect 19075 3927 19133 3928
rect 19467 3968 19509 3977
rect 19467 3928 19468 3968
rect 19508 3928 19509 3968
rect 19467 3919 19509 3928
rect 24355 3968 24413 3969
rect 24355 3928 24364 3968
rect 24404 3928 24413 3968
rect 24355 3927 24413 3928
rect 24843 3968 24885 3977
rect 24843 3928 24844 3968
rect 24884 3928 24885 3968
rect 24843 3919 24885 3928
rect 25995 3968 26037 3977
rect 25995 3928 25996 3968
rect 26036 3928 26037 3968
rect 25995 3919 26037 3928
rect 27715 3968 27773 3969
rect 27715 3928 27724 3968
rect 27764 3928 27773 3968
rect 27715 3927 27773 3928
rect 32227 3968 32285 3969
rect 32227 3928 32236 3968
rect 32276 3928 32285 3968
rect 32227 3927 32285 3928
rect 32619 3968 32661 3977
rect 32619 3928 32620 3968
rect 32660 3928 32661 3968
rect 32619 3919 32661 3928
rect 37219 3968 37277 3969
rect 37219 3928 37228 3968
rect 37268 3928 37277 3968
rect 37219 3927 37277 3928
rect 37995 3968 38037 3977
rect 37995 3928 37996 3968
rect 38036 3928 38037 3968
rect 37995 3919 38037 3928
rect 38371 3968 38429 3969
rect 38371 3928 38380 3968
rect 38420 3928 38429 3968
rect 38371 3927 38429 3928
rect 41259 3968 41301 3977
rect 41259 3928 41260 3968
rect 41300 3928 41301 3968
rect 41259 3919 41301 3928
rect 42019 3968 42077 3969
rect 42019 3928 42028 3968
rect 42068 3928 42077 3968
rect 42019 3927 42077 3928
rect 42411 3968 42453 3977
rect 42411 3928 42412 3968
rect 42452 3928 42453 3968
rect 42411 3919 42453 3928
rect 44331 3968 44373 3977
rect 44331 3928 44332 3968
rect 44372 3928 44373 3968
rect 44331 3919 44373 3928
rect 44811 3968 44853 3977
rect 44811 3928 44812 3968
rect 44852 3928 44853 3968
rect 44811 3919 44853 3928
rect 46059 3968 46101 3977
rect 46059 3928 46060 3968
rect 46100 3928 46101 3968
rect 46059 3919 46101 3928
rect 48171 3968 48213 3977
rect 48171 3928 48172 3968
rect 48212 3928 48213 3968
rect 48171 3919 48213 3928
rect 48651 3968 48693 3977
rect 48651 3928 48652 3968
rect 48692 3928 48693 3968
rect 48651 3919 48693 3928
rect 51243 3968 51285 3977
rect 51243 3928 51244 3968
rect 51284 3928 51285 3968
rect 51243 3919 51285 3928
rect 53163 3968 53205 3977
rect 53163 3928 53164 3968
rect 53204 3928 53205 3968
rect 53163 3919 53205 3928
rect 53739 3968 53781 3977
rect 53739 3928 53740 3968
rect 53780 3928 53781 3968
rect 53739 3919 53781 3928
rect 55083 3968 55125 3977
rect 55083 3928 55084 3968
rect 55124 3928 55125 3968
rect 55083 3919 55125 3928
rect 58347 3968 58389 3977
rect 58347 3928 58348 3968
rect 58388 3928 58389 3968
rect 58347 3919 58389 3928
rect 59211 3968 59253 3977
rect 59211 3928 59212 3968
rect 59252 3928 59253 3968
rect 59211 3919 59253 3928
rect 59499 3968 59541 3977
rect 59499 3928 59500 3968
rect 59540 3928 59541 3968
rect 59499 3919 59541 3928
rect 61315 3968 61373 3969
rect 61315 3928 61324 3968
rect 61364 3928 61373 3968
rect 61315 3927 61373 3928
rect 61603 3968 61661 3969
rect 61603 3928 61612 3968
rect 61652 3928 61661 3968
rect 61603 3927 61661 3928
rect 61795 3968 61853 3969
rect 61795 3928 61804 3968
rect 61844 3928 61853 3968
rect 61795 3927 61853 3928
rect 62083 3968 62141 3969
rect 62083 3928 62092 3968
rect 62132 3928 62141 3968
rect 62083 3927 62141 3928
rect 66307 3968 66365 3969
rect 66307 3928 66316 3968
rect 66356 3928 66365 3968
rect 66307 3927 66365 3928
rect 66595 3968 66653 3969
rect 66595 3928 66604 3968
rect 66644 3928 66653 3968
rect 66595 3927 66653 3928
rect 68419 3968 68477 3969
rect 68419 3928 68428 3968
rect 68468 3928 68477 3968
rect 68419 3927 68477 3928
rect 68707 3968 68765 3969
rect 68707 3928 68716 3968
rect 68756 3928 68765 3968
rect 68707 3927 68765 3928
rect 74091 3968 74133 3977
rect 74091 3928 74092 3968
rect 74132 3928 74133 3968
rect 74091 3919 74133 3928
rect 74755 3968 74813 3969
rect 74755 3928 74764 3968
rect 74804 3928 74813 3968
rect 74755 3927 74813 3928
rect 80707 3968 80765 3969
rect 80707 3928 80716 3968
rect 80756 3928 80765 3968
rect 80707 3927 80765 3928
rect 80995 3968 81053 3969
rect 80995 3928 81004 3968
rect 81044 3928 81053 3968
rect 80995 3927 81053 3928
rect 86563 3968 86621 3969
rect 86563 3928 86572 3968
rect 86612 3928 86621 3968
rect 86563 3927 86621 3928
rect 86851 3968 86909 3969
rect 86851 3928 86860 3968
rect 86900 3928 86909 3968
rect 86851 3927 86909 3928
rect 91939 3968 91997 3969
rect 91939 3928 91948 3968
rect 91988 3928 91997 3968
rect 91939 3927 91997 3928
rect 92227 3968 92285 3969
rect 92227 3928 92236 3968
rect 92276 3928 92285 3968
rect 92227 3927 92285 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 33675 3548 33717 3557
rect 33675 3508 33676 3548
rect 33716 3508 33717 3548
rect 33675 3499 33717 3508
rect 7267 3485 7325 3486
rect 1899 3464 1941 3473
rect 1899 3424 1900 3464
rect 1940 3424 1941 3464
rect 1899 3415 1941 3424
rect 2083 3464 2141 3465
rect 2083 3424 2092 3464
rect 2132 3424 2141 3464
rect 2083 3423 2141 3424
rect 4203 3464 4245 3473
rect 4203 3424 4204 3464
rect 4244 3424 4245 3464
rect 4203 3415 4245 3424
rect 4387 3464 4445 3465
rect 4387 3424 4396 3464
rect 4436 3424 4445 3464
rect 4387 3423 4445 3424
rect 4587 3464 4629 3473
rect 4587 3424 4588 3464
rect 4628 3424 4629 3464
rect 4587 3415 4629 3424
rect 4771 3464 4829 3465
rect 4771 3424 4780 3464
rect 4820 3424 4829 3464
rect 4771 3423 4829 3424
rect 4971 3464 5013 3473
rect 4971 3424 4972 3464
rect 5012 3424 5013 3464
rect 4971 3415 5013 3424
rect 5155 3464 5213 3465
rect 5155 3424 5164 3464
rect 5204 3424 5213 3464
rect 5155 3423 5213 3424
rect 5739 3464 5781 3473
rect 5739 3424 5740 3464
rect 5780 3424 5781 3464
rect 5739 3415 5781 3424
rect 5923 3464 5981 3465
rect 5923 3424 5932 3464
rect 5972 3424 5981 3464
rect 5923 3423 5981 3424
rect 6883 3464 6941 3465
rect 6883 3424 6892 3464
rect 6932 3424 6941 3464
rect 6883 3423 6941 3424
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7267 3445 7276 3485
rect 7316 3445 7325 3485
rect 7267 3444 7325 3445
rect 7467 3464 7509 3473
rect 7083 3415 7125 3424
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7651 3464 7709 3465
rect 7651 3424 7660 3464
rect 7700 3424 7709 3464
rect 7651 3423 7709 3424
rect 7851 3464 7893 3473
rect 7851 3424 7852 3464
rect 7892 3424 7893 3464
rect 7851 3415 7893 3424
rect 8419 3464 8477 3465
rect 8419 3424 8428 3464
rect 8468 3424 8477 3464
rect 8419 3423 8477 3424
rect 8619 3464 8661 3473
rect 8619 3424 8620 3464
rect 8660 3424 8661 3464
rect 8619 3415 8661 3424
rect 8803 3464 8861 3465
rect 8803 3424 8812 3464
rect 8852 3424 8861 3464
rect 8803 3423 8861 3424
rect 9003 3464 9045 3473
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9187 3464 9245 3465
rect 9187 3424 9196 3464
rect 9236 3424 9245 3464
rect 9187 3423 9245 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 9571 3464 9629 3465
rect 9571 3424 9580 3464
rect 9620 3424 9629 3464
rect 9571 3423 9629 3424
rect 9771 3464 9813 3473
rect 9771 3424 9772 3464
rect 9812 3424 9813 3464
rect 9771 3415 9813 3424
rect 9955 3464 10013 3465
rect 9955 3424 9964 3464
rect 10004 3424 10013 3464
rect 9955 3423 10013 3424
rect 10155 3464 10197 3473
rect 10155 3424 10156 3464
rect 10196 3424 10197 3464
rect 10155 3415 10197 3424
rect 10339 3464 10397 3465
rect 10339 3424 10348 3464
rect 10388 3424 10397 3464
rect 10339 3423 10397 3424
rect 10539 3464 10581 3473
rect 10539 3424 10540 3464
rect 10580 3424 10581 3464
rect 10539 3415 10581 3424
rect 10723 3464 10781 3465
rect 10723 3424 10732 3464
rect 10772 3424 10781 3464
rect 10723 3423 10781 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 11107 3464 11165 3465
rect 11107 3424 11116 3464
rect 11156 3424 11165 3464
rect 11107 3423 11165 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11491 3464 11549 3465
rect 11491 3424 11500 3464
rect 11540 3424 11549 3464
rect 11491 3423 11549 3424
rect 11691 3464 11733 3473
rect 11691 3424 11692 3464
rect 11732 3424 11733 3464
rect 11691 3415 11733 3424
rect 11875 3464 11933 3465
rect 11875 3424 11884 3464
rect 11924 3424 11933 3464
rect 11875 3423 11933 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 12259 3464 12317 3465
rect 12259 3424 12268 3464
rect 12308 3424 12317 3464
rect 12259 3423 12317 3424
rect 12459 3464 12501 3473
rect 12459 3424 12460 3464
rect 12500 3424 12501 3464
rect 12459 3415 12501 3424
rect 13027 3464 13085 3465
rect 13027 3424 13036 3464
rect 13076 3424 13085 3464
rect 13027 3423 13085 3424
rect 13227 3464 13269 3473
rect 13227 3424 13228 3464
rect 13268 3424 13269 3464
rect 13227 3415 13269 3424
rect 13411 3464 13469 3465
rect 13411 3424 13420 3464
rect 13460 3424 13469 3464
rect 13411 3423 13469 3424
rect 13611 3464 13653 3473
rect 13611 3424 13612 3464
rect 13652 3424 13653 3464
rect 13611 3415 13653 3424
rect 13795 3464 13853 3465
rect 13795 3424 13804 3464
rect 13844 3424 13853 3464
rect 13795 3423 13853 3424
rect 13995 3464 14037 3473
rect 13995 3424 13996 3464
rect 14036 3424 14037 3464
rect 13995 3415 14037 3424
rect 14283 3464 14325 3473
rect 14283 3424 14284 3464
rect 14324 3424 14325 3464
rect 14283 3415 14325 3424
rect 14467 3464 14525 3465
rect 14467 3424 14476 3464
rect 14516 3424 14525 3464
rect 14467 3423 14525 3424
rect 14667 3464 14709 3473
rect 14667 3424 14668 3464
rect 14708 3424 14709 3464
rect 14667 3415 14709 3424
rect 14851 3464 14909 3465
rect 14851 3424 14860 3464
rect 14900 3424 14909 3464
rect 14851 3423 14909 3424
rect 15051 3464 15093 3473
rect 15051 3424 15052 3464
rect 15092 3424 15093 3464
rect 15051 3415 15093 3424
rect 15235 3464 15293 3465
rect 15235 3424 15244 3464
rect 15284 3424 15293 3464
rect 15235 3423 15293 3424
rect 15435 3464 15477 3473
rect 15435 3424 15436 3464
rect 15476 3424 15477 3464
rect 15435 3415 15477 3424
rect 15619 3464 15677 3465
rect 15619 3424 15628 3464
rect 15668 3424 15677 3464
rect 15619 3423 15677 3424
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 16003 3464 16061 3465
rect 16003 3424 16012 3464
rect 16052 3424 16061 3464
rect 16003 3423 16061 3424
rect 16203 3464 16245 3473
rect 16203 3424 16204 3464
rect 16244 3424 16245 3464
rect 16203 3415 16245 3424
rect 16387 3464 16445 3465
rect 16387 3424 16396 3464
rect 16436 3424 16445 3464
rect 16387 3423 16445 3424
rect 16587 3464 16629 3473
rect 16587 3424 16588 3464
rect 16628 3424 16629 3464
rect 16587 3415 16629 3424
rect 16771 3464 16829 3465
rect 16771 3424 16780 3464
rect 16820 3424 16829 3464
rect 16771 3423 16829 3424
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 17155 3464 17213 3465
rect 17155 3424 17164 3464
rect 17204 3424 17213 3464
rect 17155 3423 17213 3424
rect 17355 3464 17397 3473
rect 17355 3424 17356 3464
rect 17396 3424 17397 3464
rect 17355 3415 17397 3424
rect 17539 3464 17597 3465
rect 17539 3424 17548 3464
rect 17588 3424 17597 3464
rect 17539 3423 17597 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 17923 3464 17981 3465
rect 17923 3424 17932 3464
rect 17972 3424 17981 3464
rect 17923 3423 17981 3424
rect 18123 3464 18165 3473
rect 18123 3424 18124 3464
rect 18164 3424 18165 3464
rect 18123 3415 18165 3424
rect 18307 3464 18365 3465
rect 18307 3424 18316 3464
rect 18356 3424 18365 3464
rect 18307 3423 18365 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18691 3464 18749 3465
rect 18691 3424 18700 3464
rect 18740 3424 18749 3464
rect 18691 3423 18749 3424
rect 18883 3464 18941 3465
rect 18883 3424 18892 3464
rect 18932 3424 18941 3464
rect 18883 3423 18941 3424
rect 19083 3464 19125 3473
rect 19083 3424 19084 3464
rect 19124 3424 19125 3464
rect 19083 3415 19125 3424
rect 19171 3464 19229 3465
rect 19171 3424 19180 3464
rect 19220 3424 19229 3464
rect 19171 3423 19229 3424
rect 19939 3464 19997 3465
rect 19939 3424 19948 3464
rect 19988 3424 19997 3464
rect 20707 3464 20765 3465
rect 19939 3423 19997 3424
rect 20148 3449 20190 3458
rect 20148 3409 20149 3449
rect 20189 3409 20190 3449
rect 20707 3424 20716 3464
rect 20756 3424 20765 3464
rect 20707 3423 20765 3424
rect 20907 3464 20949 3473
rect 20907 3424 20908 3464
rect 20948 3424 20949 3464
rect 20907 3415 20949 3424
rect 21091 3464 21149 3465
rect 21091 3424 21100 3464
rect 21140 3424 21149 3464
rect 21091 3423 21149 3424
rect 21291 3464 21333 3473
rect 21291 3424 21292 3464
rect 21332 3424 21333 3464
rect 21291 3415 21333 3424
rect 21475 3464 21533 3465
rect 21475 3424 21484 3464
rect 21524 3424 21533 3464
rect 21475 3423 21533 3424
rect 21675 3464 21717 3473
rect 21675 3424 21676 3464
rect 21716 3424 21717 3464
rect 21675 3415 21717 3424
rect 22155 3464 22197 3473
rect 22155 3424 22156 3464
rect 22196 3424 22197 3464
rect 22155 3415 22197 3424
rect 22339 3464 22397 3465
rect 22339 3424 22348 3464
rect 22388 3424 22397 3464
rect 22339 3423 22397 3424
rect 22539 3464 22581 3473
rect 22539 3424 22540 3464
rect 22580 3424 22581 3464
rect 22539 3415 22581 3424
rect 22723 3464 22781 3465
rect 22723 3424 22732 3464
rect 22772 3424 22781 3464
rect 22723 3423 22781 3424
rect 22923 3464 22965 3473
rect 22923 3424 22924 3464
rect 22964 3424 22965 3464
rect 22923 3415 22965 3424
rect 23107 3464 23165 3465
rect 23107 3424 23116 3464
rect 23156 3424 23165 3464
rect 23107 3423 23165 3424
rect 23595 3464 23637 3473
rect 23595 3424 23596 3464
rect 23636 3424 23637 3464
rect 23595 3415 23637 3424
rect 23779 3464 23837 3465
rect 23779 3424 23788 3464
rect 23828 3424 23837 3464
rect 23779 3423 23837 3424
rect 23979 3464 24021 3473
rect 23979 3424 23980 3464
rect 24020 3424 24021 3464
rect 23979 3415 24021 3424
rect 24163 3464 24221 3465
rect 24163 3424 24172 3464
rect 24212 3424 24221 3464
rect 24163 3423 24221 3424
rect 24363 3464 24405 3473
rect 24363 3424 24364 3464
rect 24404 3424 24405 3464
rect 24363 3415 24405 3424
rect 24547 3464 24605 3465
rect 24547 3424 24556 3464
rect 24596 3424 24605 3464
rect 24547 3423 24605 3424
rect 25315 3464 25373 3465
rect 25315 3424 25324 3464
rect 25364 3424 25373 3464
rect 25315 3423 25373 3424
rect 25515 3464 25557 3473
rect 25515 3424 25516 3464
rect 25556 3424 25557 3464
rect 25515 3415 25557 3424
rect 25699 3464 25757 3465
rect 25699 3424 25708 3464
rect 25748 3424 25757 3464
rect 25699 3423 25757 3424
rect 25899 3464 25941 3473
rect 25899 3424 25900 3464
rect 25940 3424 25941 3464
rect 25899 3415 25941 3424
rect 26083 3464 26141 3465
rect 26083 3424 26092 3464
rect 26132 3424 26141 3464
rect 26083 3423 26141 3424
rect 26283 3464 26325 3473
rect 26283 3424 26284 3464
rect 26324 3424 26325 3464
rect 26283 3415 26325 3424
rect 26763 3464 26805 3473
rect 26763 3424 26764 3464
rect 26804 3424 26805 3464
rect 26763 3415 26805 3424
rect 26947 3464 27005 3465
rect 26947 3424 26956 3464
rect 26996 3424 27005 3464
rect 26947 3423 27005 3424
rect 27147 3464 27189 3473
rect 27147 3424 27148 3464
rect 27188 3424 27189 3464
rect 27147 3415 27189 3424
rect 27331 3464 27389 3465
rect 27331 3424 27340 3464
rect 27380 3424 27389 3464
rect 27331 3423 27389 3424
rect 27619 3464 27677 3465
rect 27619 3424 27628 3464
rect 27668 3424 27677 3464
rect 27619 3423 27677 3424
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 28387 3464 28445 3465
rect 28387 3424 28396 3464
rect 28436 3424 28445 3464
rect 28387 3423 28445 3424
rect 28587 3464 28629 3473
rect 28587 3424 28588 3464
rect 28628 3424 28629 3464
rect 28587 3415 28629 3424
rect 28771 3464 28829 3465
rect 28771 3424 28780 3464
rect 28820 3424 28829 3464
rect 28771 3423 28829 3424
rect 28971 3464 29013 3473
rect 28971 3424 28972 3464
rect 29012 3424 29013 3464
rect 28971 3415 29013 3424
rect 29155 3464 29213 3465
rect 29155 3424 29164 3464
rect 29204 3424 29213 3464
rect 29155 3423 29213 3424
rect 29355 3464 29397 3473
rect 29355 3424 29356 3464
rect 29396 3424 29397 3464
rect 29355 3415 29397 3424
rect 29643 3464 29685 3473
rect 29643 3424 29644 3464
rect 29684 3424 29685 3464
rect 29643 3415 29685 3424
rect 29827 3464 29885 3465
rect 29827 3424 29836 3464
rect 29876 3424 29885 3464
rect 29827 3423 29885 3424
rect 30027 3464 30069 3473
rect 30027 3424 30028 3464
rect 30068 3424 30069 3464
rect 30027 3415 30069 3424
rect 30211 3464 30269 3465
rect 30211 3424 30220 3464
rect 30260 3424 30269 3464
rect 30211 3423 30269 3424
rect 30411 3464 30453 3473
rect 30411 3424 30412 3464
rect 30452 3424 30453 3464
rect 30411 3415 30453 3424
rect 30595 3464 30653 3465
rect 30595 3424 30604 3464
rect 30644 3424 30653 3464
rect 30595 3423 30653 3424
rect 31267 3464 31325 3465
rect 31267 3424 31276 3464
rect 31316 3424 31325 3464
rect 31267 3423 31325 3424
rect 31467 3464 31509 3473
rect 31467 3424 31468 3464
rect 31508 3424 31509 3464
rect 31467 3415 31509 3424
rect 31659 3464 31701 3473
rect 31659 3424 31660 3464
rect 31700 3424 31701 3464
rect 31659 3415 31701 3424
rect 31843 3464 31901 3465
rect 31843 3424 31852 3464
rect 31892 3424 31901 3464
rect 31843 3423 31901 3424
rect 32043 3464 32085 3473
rect 32043 3424 32044 3464
rect 32084 3424 32085 3464
rect 32043 3415 32085 3424
rect 32227 3464 32285 3465
rect 32227 3424 32236 3464
rect 32276 3424 32285 3464
rect 32227 3423 32285 3424
rect 32427 3464 32469 3473
rect 32427 3424 32428 3464
rect 32468 3424 32469 3464
rect 32427 3415 32469 3424
rect 32611 3464 32669 3465
rect 32611 3424 32620 3464
rect 32660 3424 32669 3464
rect 32611 3423 32669 3424
rect 32811 3464 32853 3473
rect 32811 3424 32812 3464
rect 32852 3424 32853 3464
rect 32811 3415 32853 3424
rect 32995 3464 33053 3465
rect 32995 3424 33004 3464
rect 33044 3424 33053 3464
rect 32995 3423 33053 3424
rect 33195 3464 33237 3473
rect 33195 3424 33196 3464
rect 33236 3424 33237 3464
rect 33195 3415 33237 3424
rect 33379 3464 33437 3465
rect 33379 3424 33388 3464
rect 33428 3424 33437 3464
rect 33379 3423 33437 3424
rect 33579 3464 33621 3473
rect 33579 3424 33580 3464
rect 33620 3424 33621 3464
rect 33579 3415 33621 3424
rect 33763 3464 33821 3465
rect 33763 3424 33772 3464
rect 33812 3424 33821 3464
rect 33763 3423 33821 3424
rect 33963 3464 34005 3473
rect 33963 3424 33964 3464
rect 34004 3424 34005 3464
rect 33963 3415 34005 3424
rect 34147 3464 34205 3465
rect 34147 3424 34156 3464
rect 34196 3424 34205 3464
rect 34147 3423 34205 3424
rect 34347 3464 34389 3473
rect 34347 3424 34348 3464
rect 34388 3424 34389 3464
rect 34347 3415 34389 3424
rect 34531 3464 34589 3465
rect 34531 3424 34540 3464
rect 34580 3424 34589 3464
rect 34531 3423 34589 3424
rect 34731 3464 34773 3473
rect 34731 3424 34732 3464
rect 34772 3424 34773 3464
rect 34731 3415 34773 3424
rect 34915 3464 34973 3465
rect 34915 3424 34924 3464
rect 34964 3424 34973 3464
rect 34915 3423 34973 3424
rect 35115 3464 35157 3473
rect 35115 3424 35116 3464
rect 35156 3424 35157 3464
rect 35115 3415 35157 3424
rect 35299 3464 35357 3465
rect 35299 3424 35308 3464
rect 35348 3424 35357 3464
rect 35299 3423 35357 3424
rect 35499 3464 35541 3473
rect 35499 3424 35500 3464
rect 35540 3424 35541 3464
rect 35499 3415 35541 3424
rect 35683 3464 35741 3465
rect 35683 3424 35692 3464
rect 35732 3424 35741 3464
rect 35683 3423 35741 3424
rect 35883 3464 35925 3473
rect 35883 3424 35884 3464
rect 35924 3424 35925 3464
rect 35883 3415 35925 3424
rect 36067 3464 36125 3465
rect 36067 3424 36076 3464
rect 36116 3424 36125 3464
rect 36067 3423 36125 3424
rect 36267 3464 36309 3473
rect 36267 3424 36268 3464
rect 36308 3424 36309 3464
rect 36267 3415 36309 3424
rect 36451 3464 36509 3465
rect 36451 3424 36460 3464
rect 36500 3424 36509 3464
rect 36451 3423 36509 3424
rect 36651 3464 36693 3473
rect 36651 3424 36652 3464
rect 36692 3424 36693 3464
rect 36651 3415 36693 3424
rect 36835 3464 36893 3465
rect 36835 3424 36844 3464
rect 36884 3424 36893 3464
rect 36835 3423 36893 3424
rect 37795 3464 37853 3465
rect 37795 3424 37804 3464
rect 37844 3424 37853 3464
rect 37795 3423 37853 3424
rect 37995 3464 38037 3473
rect 37995 3424 37996 3464
rect 38036 3424 38037 3464
rect 37995 3415 38037 3424
rect 38083 3464 38141 3465
rect 38083 3424 38092 3464
rect 38132 3424 38141 3464
rect 38083 3423 38141 3424
rect 38275 3464 38333 3465
rect 38275 3424 38284 3464
rect 38324 3424 38333 3464
rect 38275 3423 38333 3424
rect 38475 3464 38517 3473
rect 38475 3424 38476 3464
rect 38516 3424 38517 3464
rect 38475 3415 38517 3424
rect 38859 3464 38901 3473
rect 38859 3424 38860 3464
rect 38900 3424 38901 3464
rect 38859 3415 38901 3424
rect 39043 3464 39101 3465
rect 39043 3424 39052 3464
rect 39092 3424 39101 3464
rect 39043 3423 39101 3424
rect 39243 3464 39285 3473
rect 39243 3424 39244 3464
rect 39284 3424 39285 3464
rect 39243 3415 39285 3424
rect 39427 3464 39485 3465
rect 39427 3424 39436 3464
rect 39476 3424 39485 3464
rect 39427 3423 39485 3424
rect 39627 3464 39669 3473
rect 39627 3424 39628 3464
rect 39668 3424 39669 3464
rect 39627 3415 39669 3424
rect 39811 3464 39869 3465
rect 39811 3424 39820 3464
rect 39860 3424 39869 3464
rect 39811 3423 39869 3424
rect 40299 3464 40341 3473
rect 40299 3424 40300 3464
rect 40340 3424 40341 3464
rect 40299 3415 40341 3424
rect 40483 3464 40541 3465
rect 40483 3424 40492 3464
rect 40532 3424 40541 3464
rect 40483 3423 40541 3424
rect 40779 3464 40821 3473
rect 40779 3424 40780 3464
rect 40820 3424 40821 3464
rect 40779 3415 40821 3424
rect 40963 3464 41021 3465
rect 40963 3424 40972 3464
rect 41012 3424 41021 3464
rect 40963 3423 41021 3424
rect 41163 3464 41205 3473
rect 41163 3424 41164 3464
rect 41204 3424 41205 3464
rect 41163 3415 41205 3424
rect 41347 3464 41405 3465
rect 41347 3424 41356 3464
rect 41396 3424 41405 3464
rect 41347 3423 41405 3424
rect 41931 3464 41973 3473
rect 41931 3424 41932 3464
rect 41972 3424 41973 3464
rect 41931 3415 41973 3424
rect 42115 3464 42173 3465
rect 42115 3424 42124 3464
rect 42164 3424 42173 3464
rect 42115 3423 42173 3424
rect 42307 3464 42365 3465
rect 42307 3424 42316 3464
rect 42356 3424 42365 3464
rect 42307 3423 42365 3424
rect 42507 3464 42549 3473
rect 42507 3424 42508 3464
rect 42548 3424 42549 3464
rect 42507 3415 42549 3424
rect 42595 3464 42653 3465
rect 42595 3424 42604 3464
rect 42644 3424 42653 3464
rect 42595 3423 42653 3424
rect 42795 3464 42837 3473
rect 42795 3424 42796 3464
rect 42836 3424 42837 3464
rect 42795 3415 42837 3424
rect 42979 3464 43037 3465
rect 42979 3424 42988 3464
rect 43028 3424 43037 3464
rect 42979 3423 43037 3424
rect 44427 3464 44469 3473
rect 44427 3424 44428 3464
rect 44468 3424 44469 3464
rect 44427 3415 44469 3424
rect 44611 3464 44669 3465
rect 44611 3424 44620 3464
rect 44660 3424 44669 3464
rect 44611 3423 44669 3424
rect 45195 3464 45237 3473
rect 45195 3424 45196 3464
rect 45236 3424 45237 3464
rect 45195 3415 45237 3424
rect 45379 3464 45437 3465
rect 45379 3424 45388 3464
rect 45428 3424 45437 3464
rect 45379 3423 45437 3424
rect 45579 3464 45621 3473
rect 45579 3424 45580 3464
rect 45620 3424 45621 3464
rect 45579 3415 45621 3424
rect 45763 3464 45821 3465
rect 45763 3424 45772 3464
rect 45812 3424 45821 3464
rect 45763 3423 45821 3424
rect 45963 3464 46005 3473
rect 45963 3424 45964 3464
rect 46004 3424 46005 3464
rect 45963 3415 46005 3424
rect 46147 3464 46205 3465
rect 46147 3424 46156 3464
rect 46196 3424 46205 3464
rect 46147 3423 46205 3424
rect 46819 3464 46877 3465
rect 46819 3424 46828 3464
rect 46868 3424 46877 3464
rect 46819 3423 46877 3424
rect 47019 3464 47061 3473
rect 47019 3424 47020 3464
rect 47060 3424 47061 3464
rect 47019 3415 47061 3424
rect 47203 3464 47261 3465
rect 47203 3424 47212 3464
rect 47252 3424 47261 3464
rect 47203 3423 47261 3424
rect 47403 3464 47445 3473
rect 47403 3424 47404 3464
rect 47444 3424 47445 3464
rect 47403 3415 47445 3424
rect 47587 3464 47645 3465
rect 47587 3424 47596 3464
rect 47636 3424 47645 3464
rect 47587 3423 47645 3424
rect 47787 3464 47829 3473
rect 47787 3424 47788 3464
rect 47828 3424 47829 3464
rect 47787 3415 47829 3424
rect 48939 3464 48981 3473
rect 48939 3424 48940 3464
rect 48980 3424 48981 3464
rect 48939 3415 48981 3424
rect 49123 3464 49181 3465
rect 49123 3424 49132 3464
rect 49172 3424 49181 3464
rect 49123 3423 49181 3424
rect 50091 3464 50133 3473
rect 50091 3424 50092 3464
rect 50132 3424 50133 3464
rect 50091 3415 50133 3424
rect 50283 3464 50325 3473
rect 50283 3424 50284 3464
rect 50324 3424 50325 3464
rect 50283 3415 50325 3424
rect 50667 3464 50709 3473
rect 50667 3424 50668 3464
rect 50708 3424 50709 3464
rect 50667 3415 50709 3424
rect 50955 3464 50997 3473
rect 50955 3424 50956 3464
rect 50996 3424 50997 3464
rect 50955 3415 50997 3424
rect 51139 3464 51197 3465
rect 51139 3424 51148 3464
rect 51188 3424 51197 3464
rect 51139 3423 51197 3424
rect 52587 3464 52629 3473
rect 52587 3424 52588 3464
rect 52628 3424 52629 3464
rect 52587 3415 52629 3424
rect 52771 3464 52829 3465
rect 52771 3424 52780 3464
rect 52820 3424 52829 3464
rect 52771 3423 52829 3424
rect 53251 3464 53309 3465
rect 53251 3424 53260 3464
rect 53300 3424 53309 3464
rect 53251 3423 53309 3424
rect 53451 3464 53493 3473
rect 53451 3424 53452 3464
rect 53492 3424 53493 3464
rect 53451 3415 53493 3424
rect 54883 3464 54941 3465
rect 54883 3424 54892 3464
rect 54932 3424 54941 3464
rect 54883 3423 54941 3424
rect 55083 3464 55125 3473
rect 55083 3424 55084 3464
rect 55124 3424 55125 3464
rect 55083 3415 55125 3424
rect 55267 3464 55325 3465
rect 55267 3424 55276 3464
rect 55316 3424 55325 3464
rect 55267 3423 55325 3424
rect 55467 3464 55509 3473
rect 55467 3424 55468 3464
rect 55508 3424 55509 3464
rect 55467 3415 55509 3424
rect 56619 3464 56661 3473
rect 56619 3424 56620 3464
rect 56660 3424 56661 3464
rect 56619 3415 56661 3424
rect 56907 3464 56949 3473
rect 56907 3424 56908 3464
rect 56948 3424 56949 3464
rect 56907 3415 56949 3424
rect 57099 3464 57141 3473
rect 57099 3424 57100 3464
rect 57140 3424 57141 3464
rect 57099 3415 57141 3424
rect 58147 3464 58205 3465
rect 58147 3424 58156 3464
rect 58196 3424 58205 3464
rect 58147 3423 58205 3424
rect 58347 3464 58389 3473
rect 58347 3424 58348 3464
rect 58388 3424 58389 3464
rect 58635 3464 58677 3473
rect 58347 3415 58389 3424
rect 58531 3451 58589 3452
rect 58531 3411 58540 3451
rect 58580 3411 58589 3451
rect 58635 3424 58636 3464
rect 58676 3424 58677 3464
rect 58635 3415 58677 3424
rect 58819 3464 58877 3465
rect 58819 3424 58828 3464
rect 58868 3424 58877 3464
rect 58819 3423 58877 3424
rect 59011 3464 59069 3465
rect 59011 3424 59020 3464
rect 59060 3424 59069 3464
rect 59011 3423 59069 3424
rect 59115 3464 59157 3473
rect 59115 3424 59116 3464
rect 59156 3424 59157 3464
rect 59115 3415 59157 3424
rect 59299 3464 59357 3465
rect 59299 3424 59308 3464
rect 59348 3424 59357 3464
rect 59299 3423 59357 3424
rect 61603 3464 61661 3465
rect 61603 3424 61612 3464
rect 61652 3424 61661 3464
rect 61603 3423 61661 3424
rect 61803 3464 61845 3473
rect 61803 3424 61804 3464
rect 61844 3424 61845 3464
rect 61803 3415 61845 3424
rect 63139 3464 63197 3465
rect 63139 3424 63148 3464
rect 63188 3424 63197 3464
rect 63139 3423 63197 3424
rect 63339 3464 63381 3473
rect 63339 3424 63340 3464
rect 63380 3424 63381 3464
rect 63339 3415 63381 3424
rect 63811 3464 63869 3465
rect 63811 3424 63820 3464
rect 63860 3424 63869 3464
rect 63811 3423 63869 3424
rect 64011 3464 64053 3473
rect 64011 3424 64012 3464
rect 64052 3424 64053 3464
rect 64011 3415 64053 3424
rect 64195 3464 64253 3465
rect 64195 3424 64204 3464
rect 64244 3424 64253 3464
rect 64195 3423 64253 3424
rect 64395 3464 64437 3473
rect 64395 3424 64396 3464
rect 64436 3424 64437 3464
rect 64395 3415 64437 3424
rect 64579 3464 64637 3465
rect 64579 3424 64588 3464
rect 64628 3424 64637 3464
rect 64579 3423 64637 3424
rect 64779 3464 64821 3473
rect 64779 3424 64780 3464
rect 64820 3424 64821 3464
rect 64779 3415 64821 3424
rect 65251 3464 65309 3465
rect 65251 3424 65260 3464
rect 65300 3424 65309 3464
rect 65251 3423 65309 3424
rect 65451 3464 65493 3473
rect 65451 3424 65452 3464
rect 65492 3424 65493 3464
rect 65451 3415 65493 3424
rect 65635 3464 65693 3465
rect 65635 3424 65644 3464
rect 65684 3424 65693 3464
rect 65635 3423 65693 3424
rect 65835 3464 65877 3473
rect 65835 3424 65836 3464
rect 65876 3424 65877 3464
rect 65835 3415 65877 3424
rect 66019 3464 66077 3465
rect 66019 3424 66028 3464
rect 66068 3424 66077 3464
rect 66019 3423 66077 3424
rect 66219 3464 66261 3473
rect 66219 3424 66220 3464
rect 66260 3424 66261 3464
rect 66219 3415 66261 3424
rect 66787 3464 66845 3465
rect 66787 3424 66796 3464
rect 66836 3424 66845 3464
rect 66787 3423 66845 3424
rect 66987 3464 67029 3473
rect 66987 3424 66988 3464
rect 67028 3424 67029 3464
rect 66987 3415 67029 3424
rect 67171 3464 67229 3465
rect 67171 3424 67180 3464
rect 67220 3424 67229 3464
rect 67171 3423 67229 3424
rect 67371 3464 67413 3473
rect 67371 3424 67372 3464
rect 67412 3424 67413 3464
rect 67371 3415 67413 3424
rect 68611 3464 68669 3465
rect 68611 3424 68620 3464
rect 68660 3424 68669 3464
rect 68611 3423 68669 3424
rect 68811 3464 68853 3473
rect 68811 3424 68812 3464
rect 68852 3424 68853 3464
rect 68811 3415 68853 3424
rect 68995 3464 69053 3465
rect 68995 3424 69004 3464
rect 69044 3424 69053 3464
rect 68995 3423 69053 3424
rect 69195 3464 69237 3473
rect 69195 3424 69196 3464
rect 69236 3424 69237 3464
rect 69195 3415 69237 3424
rect 69379 3464 69437 3465
rect 69379 3424 69388 3464
rect 69428 3424 69437 3464
rect 69379 3423 69437 3424
rect 69579 3464 69621 3473
rect 69579 3424 69580 3464
rect 69620 3424 69621 3464
rect 69579 3415 69621 3424
rect 69763 3464 69821 3465
rect 69763 3424 69772 3464
rect 69812 3424 69821 3464
rect 69763 3423 69821 3424
rect 69963 3464 70005 3473
rect 69963 3424 69964 3464
rect 70004 3424 70005 3464
rect 69963 3415 70005 3424
rect 70147 3464 70205 3465
rect 70147 3424 70156 3464
rect 70196 3424 70205 3464
rect 70147 3423 70205 3424
rect 70347 3464 70389 3473
rect 70347 3424 70348 3464
rect 70388 3424 70389 3464
rect 70347 3415 70389 3424
rect 70531 3464 70589 3465
rect 70531 3424 70540 3464
rect 70580 3424 70589 3464
rect 70531 3423 70589 3424
rect 70731 3464 70773 3473
rect 70731 3424 70732 3464
rect 70772 3424 70773 3464
rect 70731 3415 70773 3424
rect 70915 3464 70973 3465
rect 70915 3424 70924 3464
rect 70964 3424 70973 3464
rect 70915 3423 70973 3424
rect 71115 3464 71157 3473
rect 71115 3424 71116 3464
rect 71156 3424 71157 3464
rect 71115 3415 71157 3424
rect 71299 3464 71357 3465
rect 71299 3424 71308 3464
rect 71348 3424 71357 3464
rect 71299 3423 71357 3424
rect 71499 3464 71541 3473
rect 71499 3424 71500 3464
rect 71540 3424 71541 3464
rect 71499 3415 71541 3424
rect 71683 3464 71741 3465
rect 71683 3424 71692 3464
rect 71732 3424 71741 3464
rect 71683 3423 71741 3424
rect 71883 3464 71925 3473
rect 71883 3424 71884 3464
rect 71924 3424 71925 3464
rect 71883 3415 71925 3424
rect 72067 3464 72125 3465
rect 72067 3424 72076 3464
rect 72116 3424 72125 3464
rect 72067 3423 72125 3424
rect 72267 3464 72309 3473
rect 72267 3424 72268 3464
rect 72308 3424 72309 3464
rect 72267 3415 72309 3424
rect 72451 3464 72509 3465
rect 72451 3424 72460 3464
rect 72500 3424 72509 3464
rect 72451 3423 72509 3424
rect 72651 3464 72693 3473
rect 72651 3424 72652 3464
rect 72692 3424 72693 3464
rect 72651 3415 72693 3424
rect 72835 3464 72893 3465
rect 72835 3424 72844 3464
rect 72884 3424 72893 3464
rect 72835 3423 72893 3424
rect 73035 3464 73077 3473
rect 73035 3424 73036 3464
rect 73076 3424 73077 3464
rect 73035 3415 73077 3424
rect 74947 3464 75005 3465
rect 74947 3424 74956 3464
rect 74996 3424 75005 3464
rect 74947 3423 75005 3424
rect 75147 3464 75189 3473
rect 75147 3424 75148 3464
rect 75188 3424 75189 3464
rect 75147 3415 75189 3424
rect 75331 3464 75389 3465
rect 75331 3424 75340 3464
rect 75380 3424 75389 3464
rect 75331 3423 75389 3424
rect 75531 3464 75573 3473
rect 75531 3424 75532 3464
rect 75572 3424 75573 3464
rect 75531 3415 75573 3424
rect 76003 3464 76061 3465
rect 76003 3424 76012 3464
rect 76052 3424 76061 3464
rect 76003 3423 76061 3424
rect 76203 3464 76245 3473
rect 76203 3424 76204 3464
rect 76244 3424 76245 3464
rect 76203 3415 76245 3424
rect 76387 3464 76445 3465
rect 76387 3424 76396 3464
rect 76436 3424 76445 3464
rect 76387 3423 76445 3424
rect 76587 3464 76629 3473
rect 76587 3424 76588 3464
rect 76628 3424 76629 3464
rect 76587 3415 76629 3424
rect 76771 3464 76829 3465
rect 76771 3424 76780 3464
rect 76820 3424 76829 3464
rect 76771 3423 76829 3424
rect 76971 3464 77013 3473
rect 76971 3424 76972 3464
rect 77012 3424 77013 3464
rect 76971 3415 77013 3424
rect 77451 3464 77493 3473
rect 77451 3424 77452 3464
rect 77492 3424 77493 3464
rect 77451 3415 77493 3424
rect 77635 3464 77693 3465
rect 77635 3424 77644 3464
rect 77684 3424 77693 3464
rect 77635 3423 77693 3424
rect 77923 3464 77981 3465
rect 77923 3424 77932 3464
rect 77972 3424 77981 3464
rect 77923 3423 77981 3424
rect 78123 3464 78165 3473
rect 78123 3424 78124 3464
rect 78164 3424 78165 3464
rect 78123 3415 78165 3424
rect 78307 3464 78365 3465
rect 78307 3424 78316 3464
rect 78356 3424 78365 3464
rect 78307 3423 78365 3424
rect 78507 3464 78549 3473
rect 78507 3424 78508 3464
rect 78548 3424 78549 3464
rect 78507 3415 78549 3424
rect 78987 3464 79029 3473
rect 78987 3424 78988 3464
rect 79028 3424 79029 3464
rect 78987 3415 79029 3424
rect 79171 3464 79229 3465
rect 79171 3424 79180 3464
rect 79220 3424 79229 3464
rect 79171 3423 79229 3424
rect 79371 3464 79413 3473
rect 79371 3424 79372 3464
rect 79412 3424 79413 3464
rect 79371 3415 79413 3424
rect 79555 3464 79613 3465
rect 79555 3424 79564 3464
rect 79604 3424 79613 3464
rect 79555 3423 79613 3424
rect 79755 3464 79797 3473
rect 79755 3424 79756 3464
rect 79796 3424 79797 3464
rect 79755 3415 79797 3424
rect 79939 3464 79997 3465
rect 79939 3424 79948 3464
rect 79988 3424 79997 3464
rect 79939 3423 79997 3424
rect 80139 3464 80181 3473
rect 80139 3424 80140 3464
rect 80180 3424 80181 3464
rect 80139 3415 80181 3424
rect 80323 3464 80381 3465
rect 80323 3424 80332 3464
rect 80372 3424 80381 3464
rect 80323 3423 80381 3424
rect 81091 3464 81149 3465
rect 81091 3424 81100 3464
rect 81140 3424 81149 3464
rect 81091 3423 81149 3424
rect 81291 3464 81333 3473
rect 81291 3424 81292 3464
rect 81332 3424 81333 3464
rect 81291 3415 81333 3424
rect 81475 3464 81533 3465
rect 81475 3424 81484 3464
rect 81524 3424 81533 3464
rect 81475 3423 81533 3424
rect 81675 3464 81717 3473
rect 81675 3424 81676 3464
rect 81716 3424 81717 3464
rect 81675 3415 81717 3424
rect 82147 3464 82205 3465
rect 82147 3424 82156 3464
rect 82196 3424 82205 3464
rect 82147 3423 82205 3424
rect 82347 3464 82389 3473
rect 82347 3424 82348 3464
rect 82388 3424 82389 3464
rect 82347 3415 82389 3424
rect 82531 3464 82589 3465
rect 82531 3424 82540 3464
rect 82580 3424 82589 3464
rect 82531 3423 82589 3424
rect 82731 3464 82773 3473
rect 82731 3424 82732 3464
rect 82772 3424 82773 3464
rect 82731 3415 82773 3424
rect 82915 3464 82973 3465
rect 82915 3424 82924 3464
rect 82964 3424 82973 3464
rect 82915 3423 82973 3424
rect 83115 3464 83157 3473
rect 83115 3424 83116 3464
rect 83156 3424 83157 3464
rect 83115 3415 83157 3424
rect 83595 3464 83637 3473
rect 83595 3424 83596 3464
rect 83636 3424 83637 3464
rect 83595 3415 83637 3424
rect 83779 3464 83837 3465
rect 83779 3424 83788 3464
rect 83828 3424 83837 3464
rect 83779 3423 83837 3424
rect 83979 3464 84021 3473
rect 83979 3424 83980 3464
rect 84020 3424 84021 3464
rect 83979 3415 84021 3424
rect 84163 3464 84221 3465
rect 84163 3424 84172 3464
rect 84212 3424 84221 3464
rect 84163 3423 84221 3424
rect 84363 3464 84405 3473
rect 84363 3424 84364 3464
rect 84404 3424 84405 3464
rect 84363 3415 84405 3424
rect 84547 3464 84605 3465
rect 84547 3424 84556 3464
rect 84596 3424 84605 3464
rect 84547 3423 84605 3424
rect 86851 3464 86909 3465
rect 86851 3424 86860 3464
rect 86900 3424 86909 3464
rect 86851 3423 86909 3424
rect 87051 3464 87093 3473
rect 87051 3424 87052 3464
rect 87092 3424 87093 3464
rect 87051 3415 87093 3424
rect 87235 3464 87293 3465
rect 87235 3424 87244 3464
rect 87284 3424 87293 3464
rect 87235 3423 87293 3424
rect 87435 3464 87477 3473
rect 87435 3424 87436 3464
rect 87476 3424 87477 3464
rect 87435 3415 87477 3424
rect 87619 3464 87677 3465
rect 87619 3424 87628 3464
rect 87668 3424 87677 3464
rect 87619 3423 87677 3424
rect 87819 3464 87861 3473
rect 87819 3424 87820 3464
rect 87860 3424 87861 3464
rect 87819 3415 87861 3424
rect 88003 3464 88061 3465
rect 88003 3424 88012 3464
rect 88052 3424 88061 3464
rect 88003 3423 88061 3424
rect 88203 3464 88245 3473
rect 88203 3424 88204 3464
rect 88244 3424 88245 3464
rect 88203 3415 88245 3424
rect 88387 3464 88445 3465
rect 88387 3424 88396 3464
rect 88436 3424 88445 3464
rect 88387 3423 88445 3424
rect 88587 3464 88629 3473
rect 88587 3424 88588 3464
rect 88628 3424 88629 3464
rect 88587 3415 88629 3424
rect 88771 3464 88829 3465
rect 88771 3424 88780 3464
rect 88820 3424 88829 3464
rect 88771 3423 88829 3424
rect 88971 3464 89013 3473
rect 88971 3424 88972 3464
rect 89012 3424 89013 3464
rect 88971 3415 89013 3424
rect 89155 3464 89213 3465
rect 89155 3424 89164 3464
rect 89204 3424 89213 3464
rect 89155 3423 89213 3424
rect 89355 3464 89397 3473
rect 89355 3424 89356 3464
rect 89396 3424 89397 3464
rect 89355 3415 89397 3424
rect 89539 3464 89597 3465
rect 89539 3424 89548 3464
rect 89588 3424 89597 3464
rect 89539 3423 89597 3424
rect 89739 3464 89781 3473
rect 89739 3424 89740 3464
rect 89780 3424 89781 3464
rect 89739 3415 89781 3424
rect 89923 3464 89981 3465
rect 89923 3424 89932 3464
rect 89972 3424 89981 3464
rect 89923 3423 89981 3424
rect 90123 3464 90165 3473
rect 90123 3424 90124 3464
rect 90164 3424 90165 3464
rect 90123 3415 90165 3424
rect 90307 3464 90365 3465
rect 90307 3424 90316 3464
rect 90356 3424 90365 3464
rect 90307 3423 90365 3424
rect 90507 3464 90549 3473
rect 90507 3424 90508 3464
rect 90548 3424 90549 3464
rect 90507 3415 90549 3424
rect 90691 3464 90749 3465
rect 90691 3424 90700 3464
rect 90740 3424 90749 3464
rect 90691 3423 90749 3424
rect 90891 3464 90933 3473
rect 90891 3424 90892 3464
rect 90932 3424 90933 3464
rect 90891 3415 90933 3424
rect 91075 3464 91133 3465
rect 91075 3424 91084 3464
rect 91124 3424 91133 3464
rect 91075 3423 91133 3424
rect 91275 3464 91317 3473
rect 91275 3424 91276 3464
rect 91316 3424 91317 3464
rect 91275 3415 91317 3424
rect 91459 3464 91517 3465
rect 91459 3424 91468 3464
rect 91508 3424 91517 3464
rect 91459 3423 91517 3424
rect 91659 3464 91701 3473
rect 91659 3424 91660 3464
rect 91700 3424 91701 3464
rect 91659 3415 91701 3424
rect 91843 3464 91901 3465
rect 91843 3424 91852 3464
rect 91892 3424 91901 3464
rect 91843 3423 91901 3424
rect 92043 3464 92085 3473
rect 92043 3424 92044 3464
rect 92084 3424 92085 3464
rect 92043 3415 92085 3424
rect 92227 3464 92285 3465
rect 92227 3424 92236 3464
rect 92276 3424 92285 3464
rect 92227 3423 92285 3424
rect 92427 3464 92469 3473
rect 92427 3424 92428 3464
rect 92468 3424 92469 3464
rect 92427 3415 92469 3424
rect 92619 3464 92661 3473
rect 92619 3424 92620 3464
rect 92660 3424 92661 3464
rect 92619 3415 92661 3424
rect 92803 3464 92861 3465
rect 92803 3424 92812 3464
rect 92852 3424 92861 3464
rect 92803 3423 92861 3424
rect 93283 3464 93341 3465
rect 93283 3424 93292 3464
rect 93332 3424 93341 3464
rect 93283 3423 93341 3424
rect 93483 3464 93525 3473
rect 93483 3424 93484 3464
rect 93524 3424 93525 3464
rect 93483 3415 93525 3424
rect 94051 3464 94109 3465
rect 94051 3424 94060 3464
rect 94100 3424 94109 3464
rect 94051 3423 94109 3424
rect 94251 3464 94293 3473
rect 94251 3424 94252 3464
rect 94292 3424 94293 3464
rect 94251 3415 94293 3424
rect 94435 3464 94493 3465
rect 94435 3424 94444 3464
rect 94484 3424 94493 3464
rect 94435 3423 94493 3424
rect 94635 3464 94677 3473
rect 94635 3424 94636 3464
rect 94676 3424 94677 3464
rect 94635 3415 94677 3424
rect 94819 3464 94877 3465
rect 94819 3424 94828 3464
rect 94868 3424 94877 3464
rect 94819 3423 94877 3424
rect 95019 3464 95061 3473
rect 95019 3424 95020 3464
rect 95060 3424 95061 3464
rect 95019 3415 95061 3424
rect 95491 3464 95549 3465
rect 95491 3424 95500 3464
rect 95540 3424 95549 3464
rect 95491 3423 95549 3424
rect 95691 3464 95733 3473
rect 95691 3424 95692 3464
rect 95732 3424 95733 3464
rect 95691 3415 95733 3424
rect 95971 3464 96029 3465
rect 95971 3424 95980 3464
rect 96020 3424 96029 3464
rect 95971 3423 96029 3424
rect 96171 3464 96213 3473
rect 96171 3424 96172 3464
rect 96212 3424 96213 3464
rect 96171 3415 96213 3424
rect 58531 3410 58589 3411
rect 20148 3400 20190 3409
rect 50667 3296 50709 3305
rect 50667 3256 50668 3296
rect 50708 3256 50709 3296
rect 50667 3247 50709 3256
rect 52683 3296 52725 3305
rect 52683 3256 52684 3296
rect 52724 3256 52725 3296
rect 52683 3247 52725 3256
rect 56619 3296 56661 3305
rect 56619 3256 56620 3296
rect 56660 3256 56661 3296
rect 56619 3247 56661 3256
rect 1995 3212 2037 3221
rect 1995 3172 1996 3212
rect 2036 3172 2037 3212
rect 1995 3163 2037 3172
rect 4299 3212 4341 3221
rect 4299 3172 4300 3212
rect 4340 3172 4341 3212
rect 4299 3163 4341 3172
rect 4683 3212 4725 3221
rect 4683 3172 4684 3212
rect 4724 3172 4725 3212
rect 4683 3163 4725 3172
rect 5067 3212 5109 3221
rect 5067 3172 5068 3212
rect 5108 3172 5109 3212
rect 5067 3163 5109 3172
rect 5835 3212 5877 3221
rect 5835 3172 5836 3212
rect 5876 3172 5877 3212
rect 5835 3163 5877 3172
rect 6987 3212 7029 3221
rect 6987 3172 6988 3212
rect 7028 3172 7029 3212
rect 6987 3163 7029 3172
rect 7371 3212 7413 3221
rect 7371 3172 7372 3212
rect 7412 3172 7413 3212
rect 7371 3163 7413 3172
rect 7755 3212 7797 3221
rect 7755 3172 7756 3212
rect 7796 3172 7797 3212
rect 7755 3163 7797 3172
rect 8523 3212 8565 3221
rect 8523 3172 8524 3212
rect 8564 3172 8565 3212
rect 8523 3163 8565 3172
rect 8907 3212 8949 3221
rect 8907 3172 8908 3212
rect 8948 3172 8949 3212
rect 8907 3163 8949 3172
rect 9291 3212 9333 3221
rect 9291 3172 9292 3212
rect 9332 3172 9333 3212
rect 9291 3163 9333 3172
rect 9675 3212 9717 3221
rect 9675 3172 9676 3212
rect 9716 3172 9717 3212
rect 9675 3163 9717 3172
rect 10059 3212 10101 3221
rect 10059 3172 10060 3212
rect 10100 3172 10101 3212
rect 10059 3163 10101 3172
rect 10443 3212 10485 3221
rect 10443 3172 10444 3212
rect 10484 3172 10485 3212
rect 10443 3163 10485 3172
rect 10827 3212 10869 3221
rect 10827 3172 10828 3212
rect 10868 3172 10869 3212
rect 10827 3163 10869 3172
rect 11211 3212 11253 3221
rect 11211 3172 11212 3212
rect 11252 3172 11253 3212
rect 11211 3163 11253 3172
rect 11595 3212 11637 3221
rect 11595 3172 11596 3212
rect 11636 3172 11637 3212
rect 11595 3163 11637 3172
rect 11979 3212 12021 3221
rect 11979 3172 11980 3212
rect 12020 3172 12021 3212
rect 11979 3163 12021 3172
rect 12363 3212 12405 3221
rect 12363 3172 12364 3212
rect 12404 3172 12405 3212
rect 12363 3163 12405 3172
rect 13131 3212 13173 3221
rect 13131 3172 13132 3212
rect 13172 3172 13173 3212
rect 13131 3163 13173 3172
rect 13515 3212 13557 3221
rect 13515 3172 13516 3212
rect 13556 3172 13557 3212
rect 13515 3163 13557 3172
rect 13899 3212 13941 3221
rect 13899 3172 13900 3212
rect 13940 3172 13941 3212
rect 13899 3163 13941 3172
rect 14379 3212 14421 3221
rect 14379 3172 14380 3212
rect 14420 3172 14421 3212
rect 14379 3163 14421 3172
rect 14763 3212 14805 3221
rect 14763 3172 14764 3212
rect 14804 3172 14805 3212
rect 14763 3163 14805 3172
rect 15147 3212 15189 3221
rect 15147 3172 15148 3212
rect 15188 3172 15189 3212
rect 15147 3163 15189 3172
rect 15531 3212 15573 3221
rect 15531 3172 15532 3212
rect 15572 3172 15573 3212
rect 15531 3163 15573 3172
rect 15915 3212 15957 3221
rect 15915 3172 15916 3212
rect 15956 3172 15957 3212
rect 15915 3163 15957 3172
rect 16299 3212 16341 3221
rect 16299 3172 16300 3212
rect 16340 3172 16341 3212
rect 16299 3163 16341 3172
rect 16683 3212 16725 3221
rect 16683 3172 16684 3212
rect 16724 3172 16725 3212
rect 16683 3163 16725 3172
rect 17067 3212 17109 3221
rect 17067 3172 17068 3212
rect 17108 3172 17109 3212
rect 17067 3163 17109 3172
rect 17451 3212 17493 3221
rect 17451 3172 17452 3212
rect 17492 3172 17493 3212
rect 17451 3163 17493 3172
rect 17835 3212 17877 3221
rect 17835 3172 17836 3212
rect 17876 3172 17877 3212
rect 17835 3163 17877 3172
rect 18219 3212 18261 3221
rect 18219 3172 18220 3212
rect 18260 3172 18261 3212
rect 18219 3163 18261 3172
rect 18603 3212 18645 3221
rect 18603 3172 18604 3212
rect 18644 3172 18645 3212
rect 18603 3163 18645 3172
rect 18891 3212 18933 3221
rect 18891 3172 18892 3212
rect 18932 3172 18933 3212
rect 18891 3163 18933 3172
rect 20043 3212 20085 3221
rect 20043 3172 20044 3212
rect 20084 3172 20085 3212
rect 20043 3163 20085 3172
rect 20811 3212 20853 3221
rect 20811 3172 20812 3212
rect 20852 3172 20853 3212
rect 20811 3163 20853 3172
rect 21195 3212 21237 3221
rect 21195 3172 21196 3212
rect 21236 3172 21237 3212
rect 21195 3163 21237 3172
rect 21579 3212 21621 3221
rect 21579 3172 21580 3212
rect 21620 3172 21621 3212
rect 21579 3163 21621 3172
rect 22251 3212 22293 3221
rect 22251 3172 22252 3212
rect 22292 3172 22293 3212
rect 22251 3163 22293 3172
rect 22635 3212 22677 3221
rect 22635 3172 22636 3212
rect 22676 3172 22677 3212
rect 22635 3163 22677 3172
rect 23019 3212 23061 3221
rect 23019 3172 23020 3212
rect 23060 3172 23061 3212
rect 23019 3163 23061 3172
rect 23691 3212 23733 3221
rect 23691 3172 23692 3212
rect 23732 3172 23733 3212
rect 23691 3163 23733 3172
rect 24075 3212 24117 3221
rect 24075 3172 24076 3212
rect 24116 3172 24117 3212
rect 24075 3163 24117 3172
rect 24459 3212 24501 3221
rect 24459 3172 24460 3212
rect 24500 3172 24501 3212
rect 24459 3163 24501 3172
rect 25419 3212 25461 3221
rect 25419 3172 25420 3212
rect 25460 3172 25461 3212
rect 25419 3163 25461 3172
rect 25803 3212 25845 3221
rect 25803 3172 25804 3212
rect 25844 3172 25845 3212
rect 25803 3163 25845 3172
rect 26187 3212 26229 3221
rect 26187 3172 26188 3212
rect 26228 3172 26229 3212
rect 26187 3163 26229 3172
rect 26859 3212 26901 3221
rect 26859 3172 26860 3212
rect 26900 3172 26901 3212
rect 26859 3163 26901 3172
rect 27243 3212 27285 3221
rect 27243 3172 27244 3212
rect 27284 3172 27285 3212
rect 27243 3163 27285 3172
rect 27723 3212 27765 3221
rect 27723 3172 27724 3212
rect 27764 3172 27765 3212
rect 27723 3163 27765 3172
rect 28491 3212 28533 3221
rect 28491 3172 28492 3212
rect 28532 3172 28533 3212
rect 28491 3163 28533 3172
rect 28875 3212 28917 3221
rect 28875 3172 28876 3212
rect 28916 3172 28917 3212
rect 28875 3163 28917 3172
rect 29259 3212 29301 3221
rect 29259 3172 29260 3212
rect 29300 3172 29301 3212
rect 29259 3163 29301 3172
rect 29739 3212 29781 3221
rect 29739 3172 29740 3212
rect 29780 3172 29781 3212
rect 29739 3163 29781 3172
rect 30123 3212 30165 3221
rect 30123 3172 30124 3212
rect 30164 3172 30165 3212
rect 30123 3163 30165 3172
rect 30507 3212 30549 3221
rect 30507 3172 30508 3212
rect 30548 3172 30549 3212
rect 30507 3163 30549 3172
rect 31371 3212 31413 3221
rect 31371 3172 31372 3212
rect 31412 3172 31413 3212
rect 31371 3163 31413 3172
rect 31755 3212 31797 3221
rect 31755 3172 31756 3212
rect 31796 3172 31797 3212
rect 31755 3163 31797 3172
rect 32139 3212 32181 3221
rect 32139 3172 32140 3212
rect 32180 3172 32181 3212
rect 32139 3163 32181 3172
rect 32523 3212 32565 3221
rect 32523 3172 32524 3212
rect 32564 3172 32565 3212
rect 32523 3163 32565 3172
rect 32907 3212 32949 3221
rect 32907 3172 32908 3212
rect 32948 3172 32949 3212
rect 32907 3163 32949 3172
rect 33291 3212 33333 3221
rect 33291 3172 33292 3212
rect 33332 3172 33333 3212
rect 33291 3163 33333 3172
rect 34059 3212 34101 3221
rect 34059 3172 34060 3212
rect 34100 3172 34101 3212
rect 34059 3163 34101 3172
rect 34443 3212 34485 3221
rect 34443 3172 34444 3212
rect 34484 3172 34485 3212
rect 34443 3163 34485 3172
rect 34827 3212 34869 3221
rect 34827 3172 34828 3212
rect 34868 3172 34869 3212
rect 34827 3163 34869 3172
rect 35211 3212 35253 3221
rect 35211 3172 35212 3212
rect 35252 3172 35253 3212
rect 35211 3163 35253 3172
rect 35595 3212 35637 3221
rect 35595 3172 35596 3212
rect 35636 3172 35637 3212
rect 35595 3163 35637 3172
rect 35979 3212 36021 3221
rect 35979 3172 35980 3212
rect 36020 3172 36021 3212
rect 35979 3163 36021 3172
rect 36363 3212 36405 3221
rect 36363 3172 36364 3212
rect 36404 3172 36405 3212
rect 36363 3163 36405 3172
rect 36747 3212 36789 3221
rect 36747 3172 36748 3212
rect 36788 3172 36789 3212
rect 36747 3163 36789 3172
rect 37803 3212 37845 3221
rect 37803 3172 37804 3212
rect 37844 3172 37845 3212
rect 37803 3163 37845 3172
rect 38379 3212 38421 3221
rect 38379 3172 38380 3212
rect 38420 3172 38421 3212
rect 38379 3163 38421 3172
rect 38955 3212 38997 3221
rect 38955 3172 38956 3212
rect 38996 3172 38997 3212
rect 38955 3163 38997 3172
rect 39339 3212 39381 3221
rect 39339 3172 39340 3212
rect 39380 3172 39381 3212
rect 39339 3163 39381 3172
rect 39723 3212 39765 3221
rect 39723 3172 39724 3212
rect 39764 3172 39765 3212
rect 39723 3163 39765 3172
rect 40395 3212 40437 3221
rect 40395 3172 40396 3212
rect 40436 3172 40437 3212
rect 40395 3163 40437 3172
rect 40875 3212 40917 3221
rect 40875 3172 40876 3212
rect 40916 3172 40917 3212
rect 40875 3163 40917 3172
rect 41259 3212 41301 3221
rect 41259 3172 41260 3212
rect 41300 3172 41301 3212
rect 41259 3163 41301 3172
rect 42027 3212 42069 3221
rect 42027 3172 42028 3212
rect 42068 3172 42069 3212
rect 42027 3163 42069 3172
rect 42315 3212 42357 3221
rect 42315 3172 42316 3212
rect 42356 3172 42357 3212
rect 42315 3163 42357 3172
rect 42891 3212 42933 3221
rect 42891 3172 42892 3212
rect 42932 3172 42933 3212
rect 42891 3163 42933 3172
rect 44523 3212 44565 3221
rect 44523 3172 44524 3212
rect 44564 3172 44565 3212
rect 44523 3163 44565 3172
rect 45291 3212 45333 3221
rect 45291 3172 45292 3212
rect 45332 3172 45333 3212
rect 45291 3163 45333 3172
rect 45675 3212 45717 3221
rect 45675 3172 45676 3212
rect 45716 3172 45717 3212
rect 45675 3163 45717 3172
rect 46059 3212 46101 3221
rect 46059 3172 46060 3212
rect 46100 3172 46101 3212
rect 46059 3163 46101 3172
rect 46923 3212 46965 3221
rect 46923 3172 46924 3212
rect 46964 3172 46965 3212
rect 46923 3163 46965 3172
rect 47307 3212 47349 3221
rect 47307 3172 47308 3212
rect 47348 3172 47349 3212
rect 47307 3163 47349 3172
rect 47691 3212 47733 3221
rect 47691 3172 47692 3212
rect 47732 3172 47733 3212
rect 47691 3163 47733 3172
rect 49035 3212 49077 3221
rect 49035 3172 49036 3212
rect 49076 3172 49077 3212
rect 49035 3163 49077 3172
rect 50283 3212 50325 3221
rect 50283 3172 50284 3212
rect 50324 3172 50325 3212
rect 50283 3163 50325 3172
rect 50475 3212 50517 3221
rect 50475 3172 50476 3212
rect 50516 3172 50517 3212
rect 50475 3163 50517 3172
rect 51051 3212 51093 3221
rect 51051 3172 51052 3212
rect 51092 3172 51093 3212
rect 51051 3163 51093 3172
rect 53355 3212 53397 3221
rect 53355 3172 53356 3212
rect 53396 3172 53397 3212
rect 53355 3163 53397 3172
rect 54987 3212 55029 3221
rect 54987 3172 54988 3212
rect 55028 3172 55029 3212
rect 54987 3163 55029 3172
rect 55371 3212 55413 3221
rect 55371 3172 55372 3212
rect 55412 3172 55413 3212
rect 55371 3163 55413 3172
rect 56427 3212 56469 3221
rect 56427 3172 56428 3212
rect 56468 3172 56469 3212
rect 56427 3163 56469 3172
rect 56907 3212 56949 3221
rect 56907 3172 56908 3212
rect 56948 3172 56949 3212
rect 56907 3163 56949 3172
rect 58251 3212 58293 3221
rect 58251 3172 58252 3212
rect 58292 3172 58293 3212
rect 58251 3163 58293 3172
rect 58827 3212 58869 3221
rect 58827 3172 58828 3212
rect 58868 3172 58869 3212
rect 58827 3163 58869 3172
rect 59307 3212 59349 3221
rect 59307 3172 59308 3212
rect 59348 3172 59349 3212
rect 59307 3163 59349 3172
rect 61707 3212 61749 3221
rect 61707 3172 61708 3212
rect 61748 3172 61749 3212
rect 61707 3163 61749 3172
rect 63243 3212 63285 3221
rect 63243 3172 63244 3212
rect 63284 3172 63285 3212
rect 63243 3163 63285 3172
rect 63915 3212 63957 3221
rect 63915 3172 63916 3212
rect 63956 3172 63957 3212
rect 63915 3163 63957 3172
rect 64299 3212 64341 3221
rect 64299 3172 64300 3212
rect 64340 3172 64341 3212
rect 64299 3163 64341 3172
rect 64683 3212 64725 3221
rect 64683 3172 64684 3212
rect 64724 3172 64725 3212
rect 64683 3163 64725 3172
rect 65355 3212 65397 3221
rect 65355 3172 65356 3212
rect 65396 3172 65397 3212
rect 65355 3163 65397 3172
rect 65739 3212 65781 3221
rect 65739 3172 65740 3212
rect 65780 3172 65781 3212
rect 65739 3163 65781 3172
rect 66123 3212 66165 3221
rect 66123 3172 66124 3212
rect 66164 3172 66165 3212
rect 66123 3163 66165 3172
rect 66891 3212 66933 3221
rect 66891 3172 66892 3212
rect 66932 3172 66933 3212
rect 66891 3163 66933 3172
rect 67275 3212 67317 3221
rect 67275 3172 67276 3212
rect 67316 3172 67317 3212
rect 67275 3163 67317 3172
rect 68715 3212 68757 3221
rect 68715 3172 68716 3212
rect 68756 3172 68757 3212
rect 68715 3163 68757 3172
rect 69099 3212 69141 3221
rect 69099 3172 69100 3212
rect 69140 3172 69141 3212
rect 69099 3163 69141 3172
rect 69483 3212 69525 3221
rect 69483 3172 69484 3212
rect 69524 3172 69525 3212
rect 69483 3163 69525 3172
rect 69867 3212 69909 3221
rect 69867 3172 69868 3212
rect 69908 3172 69909 3212
rect 69867 3163 69909 3172
rect 70251 3212 70293 3221
rect 70251 3172 70252 3212
rect 70292 3172 70293 3212
rect 70251 3163 70293 3172
rect 70635 3212 70677 3221
rect 70635 3172 70636 3212
rect 70676 3172 70677 3212
rect 70635 3163 70677 3172
rect 71019 3212 71061 3221
rect 71019 3172 71020 3212
rect 71060 3172 71061 3212
rect 71019 3163 71061 3172
rect 71403 3212 71445 3221
rect 71403 3172 71404 3212
rect 71444 3172 71445 3212
rect 71403 3163 71445 3172
rect 71787 3212 71829 3221
rect 71787 3172 71788 3212
rect 71828 3172 71829 3212
rect 71787 3163 71829 3172
rect 72171 3212 72213 3221
rect 72171 3172 72172 3212
rect 72212 3172 72213 3212
rect 72171 3163 72213 3172
rect 72555 3212 72597 3221
rect 72555 3172 72556 3212
rect 72596 3172 72597 3212
rect 72555 3163 72597 3172
rect 72939 3212 72981 3221
rect 72939 3172 72940 3212
rect 72980 3172 72981 3212
rect 72939 3163 72981 3172
rect 75051 3212 75093 3221
rect 75051 3172 75052 3212
rect 75092 3172 75093 3212
rect 75051 3163 75093 3172
rect 75435 3212 75477 3221
rect 75435 3172 75436 3212
rect 75476 3172 75477 3212
rect 75435 3163 75477 3172
rect 76107 3212 76149 3221
rect 76107 3172 76108 3212
rect 76148 3172 76149 3212
rect 76107 3163 76149 3172
rect 76491 3212 76533 3221
rect 76491 3172 76492 3212
rect 76532 3172 76533 3212
rect 76491 3163 76533 3172
rect 76875 3212 76917 3221
rect 76875 3172 76876 3212
rect 76916 3172 76917 3212
rect 76875 3163 76917 3172
rect 77547 3212 77589 3221
rect 77547 3172 77548 3212
rect 77588 3172 77589 3212
rect 77547 3163 77589 3172
rect 78027 3212 78069 3221
rect 78027 3172 78028 3212
rect 78068 3172 78069 3212
rect 78027 3163 78069 3172
rect 78411 3212 78453 3221
rect 78411 3172 78412 3212
rect 78452 3172 78453 3212
rect 78411 3163 78453 3172
rect 79083 3212 79125 3221
rect 79083 3172 79084 3212
rect 79124 3172 79125 3212
rect 79083 3163 79125 3172
rect 79467 3212 79509 3221
rect 79467 3172 79468 3212
rect 79508 3172 79509 3212
rect 79467 3163 79509 3172
rect 79851 3212 79893 3221
rect 79851 3172 79852 3212
rect 79892 3172 79893 3212
rect 79851 3163 79893 3172
rect 80235 3212 80277 3221
rect 80235 3172 80236 3212
rect 80276 3172 80277 3212
rect 80235 3163 80277 3172
rect 81195 3212 81237 3221
rect 81195 3172 81196 3212
rect 81236 3172 81237 3212
rect 81195 3163 81237 3172
rect 81579 3212 81621 3221
rect 81579 3172 81580 3212
rect 81620 3172 81621 3212
rect 81579 3163 81621 3172
rect 82251 3212 82293 3221
rect 82251 3172 82252 3212
rect 82292 3172 82293 3212
rect 82251 3163 82293 3172
rect 82635 3212 82677 3221
rect 82635 3172 82636 3212
rect 82676 3172 82677 3212
rect 82635 3163 82677 3172
rect 83019 3212 83061 3221
rect 83019 3172 83020 3212
rect 83060 3172 83061 3212
rect 83019 3163 83061 3172
rect 83691 3212 83733 3221
rect 83691 3172 83692 3212
rect 83732 3172 83733 3212
rect 83691 3163 83733 3172
rect 84075 3212 84117 3221
rect 84075 3172 84076 3212
rect 84116 3172 84117 3212
rect 84075 3163 84117 3172
rect 84459 3212 84501 3221
rect 84459 3172 84460 3212
rect 84500 3172 84501 3212
rect 84459 3163 84501 3172
rect 86955 3212 86997 3221
rect 86955 3172 86956 3212
rect 86996 3172 86997 3212
rect 86955 3163 86997 3172
rect 87339 3212 87381 3221
rect 87339 3172 87340 3212
rect 87380 3172 87381 3212
rect 87339 3163 87381 3172
rect 87723 3212 87765 3221
rect 87723 3172 87724 3212
rect 87764 3172 87765 3212
rect 87723 3163 87765 3172
rect 88107 3212 88149 3221
rect 88107 3172 88108 3212
rect 88148 3172 88149 3212
rect 88107 3163 88149 3172
rect 88491 3212 88533 3221
rect 88491 3172 88492 3212
rect 88532 3172 88533 3212
rect 88491 3163 88533 3172
rect 88875 3212 88917 3221
rect 88875 3172 88876 3212
rect 88916 3172 88917 3212
rect 88875 3163 88917 3172
rect 89259 3212 89301 3221
rect 89259 3172 89260 3212
rect 89300 3172 89301 3212
rect 89259 3163 89301 3172
rect 89643 3212 89685 3221
rect 89643 3172 89644 3212
rect 89684 3172 89685 3212
rect 89643 3163 89685 3172
rect 90027 3212 90069 3221
rect 90027 3172 90028 3212
rect 90068 3172 90069 3212
rect 90027 3163 90069 3172
rect 90411 3212 90453 3221
rect 90411 3172 90412 3212
rect 90452 3172 90453 3212
rect 90411 3163 90453 3172
rect 90795 3212 90837 3221
rect 90795 3172 90796 3212
rect 90836 3172 90837 3212
rect 90795 3163 90837 3172
rect 91179 3212 91221 3221
rect 91179 3172 91180 3212
rect 91220 3172 91221 3212
rect 91179 3163 91221 3172
rect 91563 3212 91605 3221
rect 91563 3172 91564 3212
rect 91604 3172 91605 3212
rect 91563 3163 91605 3172
rect 91947 3212 91989 3221
rect 91947 3172 91948 3212
rect 91988 3172 91989 3212
rect 91947 3163 91989 3172
rect 92331 3212 92373 3221
rect 92331 3172 92332 3212
rect 92372 3172 92373 3212
rect 92331 3163 92373 3172
rect 92715 3212 92757 3221
rect 92715 3172 92716 3212
rect 92756 3172 92757 3212
rect 92715 3163 92757 3172
rect 93387 3212 93429 3221
rect 93387 3172 93388 3212
rect 93428 3172 93429 3212
rect 93387 3163 93429 3172
rect 94155 3212 94197 3221
rect 94155 3172 94156 3212
rect 94196 3172 94197 3212
rect 94155 3163 94197 3172
rect 94539 3212 94581 3221
rect 94539 3172 94540 3212
rect 94580 3172 94581 3212
rect 94539 3163 94581 3172
rect 94923 3212 94965 3221
rect 94923 3172 94924 3212
rect 94964 3172 94965 3212
rect 94923 3163 94965 3172
rect 95595 3212 95637 3221
rect 95595 3172 95596 3212
rect 95636 3172 95637 3212
rect 95595 3163 95637 3172
rect 96075 3212 96117 3221
rect 96075 3172 96076 3212
rect 96116 3172 96117 3212
rect 96075 3163 96117 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 54891 2792 54933 2801
rect 54891 2752 54892 2792
rect 54932 2752 54933 2792
rect 55755 2792 55797 2801
rect 54891 2743 54933 2752
rect 55275 2766 55317 2775
rect 55275 2726 55276 2766
rect 55316 2726 55317 2766
rect 55755 2752 55756 2792
rect 55796 2752 55797 2792
rect 55755 2743 55797 2752
rect 58635 2792 58677 2801
rect 58635 2752 58636 2792
rect 58676 2752 58677 2792
rect 58635 2743 58677 2752
rect 60939 2792 60981 2801
rect 60939 2752 60940 2792
rect 60980 2752 60981 2792
rect 60939 2743 60981 2752
rect 61419 2792 61461 2801
rect 61419 2752 61420 2792
rect 61460 2752 61461 2792
rect 61419 2743 61461 2752
rect 55275 2717 55317 2726
rect 73892 2647 73950 2648
rect 1603 2624 1661 2625
rect 1603 2584 1612 2624
rect 1652 2584 1661 2624
rect 1603 2583 1661 2584
rect 1803 2624 1845 2633
rect 1803 2584 1804 2624
rect 1844 2584 1845 2624
rect 1803 2575 1845 2584
rect 2091 2624 2133 2633
rect 2091 2584 2092 2624
rect 2132 2584 2133 2624
rect 2091 2575 2133 2584
rect 2275 2624 2333 2625
rect 2275 2584 2284 2624
rect 2324 2584 2333 2624
rect 2275 2583 2333 2584
rect 2475 2624 2517 2633
rect 2475 2584 2476 2624
rect 2516 2584 2517 2624
rect 2475 2575 2517 2584
rect 2659 2624 2717 2625
rect 2659 2584 2668 2624
rect 2708 2584 2717 2624
rect 2659 2583 2717 2584
rect 2955 2624 2997 2633
rect 2955 2584 2956 2624
rect 2996 2584 2997 2624
rect 2955 2575 2997 2584
rect 3139 2624 3197 2625
rect 3139 2584 3148 2624
rect 3188 2584 3197 2624
rect 3139 2583 3197 2584
rect 3339 2624 3381 2633
rect 3339 2584 3340 2624
rect 3380 2584 3381 2624
rect 3339 2575 3381 2584
rect 3523 2624 3581 2625
rect 3523 2584 3532 2624
rect 3572 2584 3581 2624
rect 3523 2583 3581 2584
rect 3723 2624 3765 2633
rect 3723 2584 3724 2624
rect 3764 2584 3765 2624
rect 3723 2575 3765 2584
rect 3907 2624 3965 2625
rect 3907 2584 3916 2624
rect 3956 2584 3965 2624
rect 3907 2583 3965 2584
rect 6123 2624 6165 2633
rect 6123 2584 6124 2624
rect 6164 2584 6165 2624
rect 6123 2575 6165 2584
rect 6307 2624 6365 2625
rect 6307 2584 6316 2624
rect 6356 2584 6365 2624
rect 6307 2583 6365 2584
rect 6603 2624 6645 2633
rect 6603 2584 6604 2624
rect 6644 2584 6645 2624
rect 6603 2575 6645 2584
rect 6787 2624 6845 2625
rect 6787 2584 6796 2624
rect 6836 2584 6845 2624
rect 6787 2583 6845 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7171 2624 7229 2625
rect 7171 2584 7180 2624
rect 7220 2584 7229 2624
rect 7171 2583 7229 2584
rect 8035 2624 8093 2625
rect 8035 2584 8044 2624
rect 8084 2584 8093 2624
rect 8035 2583 8093 2584
rect 8235 2624 8277 2633
rect 8235 2584 8236 2624
rect 8276 2584 8277 2624
rect 8235 2575 8277 2584
rect 12555 2624 12597 2633
rect 12555 2584 12556 2624
rect 12596 2584 12597 2624
rect 12555 2575 12597 2584
rect 12739 2624 12797 2625
rect 12739 2584 12748 2624
rect 12788 2584 12797 2624
rect 12739 2583 12797 2584
rect 14091 2624 14133 2633
rect 14091 2584 14092 2624
rect 14132 2584 14133 2624
rect 14091 2575 14133 2584
rect 14275 2624 14333 2625
rect 14275 2584 14284 2624
rect 14324 2584 14333 2624
rect 14275 2583 14333 2584
rect 19651 2624 19709 2625
rect 19651 2584 19660 2624
rect 19700 2584 19709 2624
rect 19651 2583 19709 2584
rect 19851 2624 19893 2633
rect 19851 2584 19852 2624
rect 19892 2584 19893 2624
rect 19851 2575 19893 2584
rect 20235 2624 20277 2633
rect 20235 2584 20236 2624
rect 20276 2584 20277 2624
rect 20235 2575 20277 2584
rect 20419 2624 20477 2625
rect 20419 2584 20428 2624
rect 20468 2584 20477 2624
rect 20419 2583 20477 2584
rect 21859 2624 21917 2625
rect 21859 2584 21868 2624
rect 21908 2584 21917 2624
rect 21859 2583 21917 2584
rect 22059 2624 22101 2633
rect 22059 2584 22060 2624
rect 22100 2584 22101 2624
rect 22059 2575 22101 2584
rect 23395 2624 23453 2625
rect 23395 2584 23404 2624
rect 23444 2584 23453 2624
rect 23395 2583 23453 2584
rect 23595 2624 23637 2633
rect 23595 2584 23596 2624
rect 23636 2584 23637 2624
rect 23595 2575 23637 2584
rect 26379 2624 26421 2633
rect 26379 2584 26380 2624
rect 26420 2584 26421 2624
rect 26379 2575 26421 2584
rect 26563 2624 26621 2625
rect 26563 2584 26572 2624
rect 26612 2584 26621 2624
rect 26563 2583 26621 2584
rect 27915 2624 27957 2633
rect 27915 2584 27916 2624
rect 27956 2584 27957 2624
rect 27915 2575 27957 2584
rect 28099 2624 28157 2625
rect 28099 2584 28108 2624
rect 28148 2584 28157 2624
rect 28099 2583 28157 2584
rect 29539 2624 29597 2625
rect 29539 2584 29548 2624
rect 29588 2584 29597 2624
rect 29539 2583 29597 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 30699 2624 30741 2633
rect 30699 2584 30700 2624
rect 30740 2584 30741 2624
rect 30699 2575 30741 2584
rect 30883 2624 30941 2625
rect 30883 2584 30892 2624
rect 30932 2584 30941 2624
rect 30883 2583 30941 2584
rect 31651 2624 31709 2625
rect 31651 2584 31660 2624
rect 31700 2584 31709 2624
rect 31651 2583 31709 2584
rect 31851 2624 31893 2633
rect 31851 2584 31852 2624
rect 31892 2584 31893 2624
rect 31851 2575 31893 2584
rect 37603 2624 37661 2625
rect 37603 2584 37612 2624
rect 37652 2584 37661 2624
rect 37603 2583 37661 2584
rect 37803 2624 37845 2633
rect 37803 2584 37804 2624
rect 37844 2584 37845 2624
rect 38371 2624 38429 2625
rect 37803 2575 37845 2584
rect 38187 2611 38229 2620
rect 38187 2571 38188 2611
rect 38228 2571 38229 2611
rect 38371 2584 38380 2624
rect 38420 2584 38429 2624
rect 38371 2583 38429 2584
rect 38571 2624 38613 2633
rect 38571 2584 38572 2624
rect 38612 2584 38613 2624
rect 38571 2575 38613 2584
rect 38755 2624 38813 2625
rect 38755 2584 38764 2624
rect 38804 2584 38813 2624
rect 38755 2583 38813 2584
rect 40011 2624 40053 2633
rect 40011 2584 40012 2624
rect 40052 2584 40053 2624
rect 40011 2575 40053 2584
rect 40195 2624 40253 2625
rect 40195 2584 40204 2624
rect 40244 2584 40253 2624
rect 40195 2583 40253 2584
rect 41643 2624 41685 2633
rect 41643 2584 41644 2624
rect 41684 2584 41685 2624
rect 41643 2575 41685 2584
rect 41827 2624 41885 2625
rect 41827 2584 41836 2624
rect 41876 2584 41885 2624
rect 41827 2583 41885 2584
rect 42027 2624 42069 2633
rect 42027 2584 42028 2624
rect 42068 2584 42069 2624
rect 42027 2575 42069 2584
rect 42211 2624 42269 2625
rect 42211 2584 42220 2624
rect 42260 2584 42269 2624
rect 42211 2583 42269 2584
rect 42795 2624 42837 2633
rect 42795 2584 42796 2624
rect 42836 2584 42837 2624
rect 42795 2575 42837 2584
rect 42979 2624 43037 2625
rect 42979 2584 42988 2624
rect 43028 2584 43037 2624
rect 42979 2583 43037 2584
rect 44043 2624 44085 2633
rect 44043 2584 44044 2624
rect 44084 2584 44085 2624
rect 44043 2575 44085 2584
rect 44227 2624 44285 2625
rect 44227 2584 44236 2624
rect 44276 2584 44285 2624
rect 44227 2583 44285 2584
rect 44811 2624 44853 2633
rect 44811 2584 44812 2624
rect 44852 2584 44853 2624
rect 44811 2575 44853 2584
rect 44995 2624 45053 2625
rect 44995 2584 45004 2624
rect 45044 2584 45053 2624
rect 44995 2583 45053 2584
rect 46347 2624 46389 2633
rect 46347 2584 46348 2624
rect 46388 2584 46389 2624
rect 46347 2575 46389 2584
rect 46531 2624 46589 2625
rect 46531 2584 46540 2624
rect 46580 2584 46589 2624
rect 46531 2583 46589 2584
rect 47883 2624 47925 2633
rect 47883 2584 47884 2624
rect 47924 2584 47925 2624
rect 47883 2575 47925 2584
rect 48067 2624 48125 2625
rect 48067 2584 48076 2624
rect 48116 2584 48125 2624
rect 48067 2583 48125 2584
rect 48267 2624 48309 2633
rect 48267 2584 48268 2624
rect 48308 2584 48309 2624
rect 48267 2575 48309 2584
rect 48451 2624 48509 2625
rect 48451 2584 48460 2624
rect 48500 2584 48509 2624
rect 48451 2583 48509 2584
rect 48651 2624 48693 2633
rect 48651 2584 48652 2624
rect 48692 2584 48693 2624
rect 48651 2575 48693 2584
rect 48835 2624 48893 2625
rect 48835 2584 48844 2624
rect 48884 2584 48893 2624
rect 48835 2583 48893 2584
rect 49131 2624 49173 2633
rect 49131 2584 49132 2624
rect 49172 2584 49173 2624
rect 49131 2575 49173 2584
rect 49315 2624 49373 2625
rect 49315 2584 49324 2624
rect 49364 2584 49373 2624
rect 49315 2583 49373 2584
rect 54699 2624 54741 2633
rect 54699 2584 54700 2624
rect 54740 2584 54741 2624
rect 54699 2575 54741 2584
rect 54891 2613 54933 2622
rect 38187 2562 38229 2571
rect 54891 2573 54892 2613
rect 54932 2573 54933 2613
rect 54891 2564 54933 2573
rect 55275 2616 55317 2625
rect 55275 2576 55276 2616
rect 55316 2576 55317 2616
rect 55275 2567 55317 2576
rect 55755 2624 55797 2633
rect 55755 2584 55756 2624
rect 55796 2584 55797 2624
rect 55755 2575 55797 2584
rect 56043 2624 56085 2633
rect 56043 2584 56044 2624
rect 56084 2584 56085 2624
rect 56043 2575 56085 2584
rect 56235 2624 56277 2633
rect 56235 2584 56236 2624
rect 56276 2584 56277 2624
rect 56235 2575 56277 2584
rect 58635 2624 58677 2633
rect 58635 2584 58636 2624
rect 58676 2584 58677 2624
rect 58635 2575 58677 2584
rect 60459 2624 60501 2633
rect 60459 2584 60460 2624
rect 60500 2584 60501 2624
rect 60459 2575 60501 2584
rect 60651 2624 60693 2633
rect 60651 2584 60652 2624
rect 60692 2584 60693 2624
rect 60651 2575 60693 2584
rect 60939 2624 60981 2633
rect 60939 2584 60940 2624
rect 60980 2584 60981 2624
rect 60939 2575 60981 2584
rect 61419 2624 61461 2633
rect 61419 2584 61420 2624
rect 61460 2584 61461 2624
rect 61419 2575 61461 2584
rect 61803 2624 61845 2633
rect 61803 2584 61804 2624
rect 61844 2584 61845 2624
rect 61803 2575 61845 2584
rect 61995 2624 62037 2633
rect 61995 2584 61996 2624
rect 62036 2584 62037 2624
rect 61995 2575 62037 2584
rect 62851 2624 62909 2625
rect 62851 2584 62860 2624
rect 62900 2584 62909 2624
rect 62851 2583 62909 2584
rect 63051 2624 63093 2633
rect 63051 2584 63052 2624
rect 63092 2584 63093 2624
rect 63051 2575 63093 2584
rect 63331 2624 63389 2625
rect 63331 2584 63340 2624
rect 63380 2584 63389 2624
rect 63331 2583 63389 2584
rect 63531 2624 63573 2633
rect 63531 2584 63532 2624
rect 63572 2584 63573 2624
rect 63531 2575 63573 2584
rect 67371 2624 67413 2633
rect 67371 2584 67372 2624
rect 67412 2584 67413 2624
rect 67371 2575 67413 2584
rect 67555 2624 67613 2625
rect 67555 2584 67564 2624
rect 67604 2584 67613 2624
rect 67555 2583 67613 2584
rect 72931 2624 72989 2625
rect 72931 2584 72940 2624
rect 72980 2584 72989 2624
rect 72931 2583 72989 2584
rect 73131 2624 73173 2633
rect 73131 2584 73132 2624
rect 73172 2584 73173 2624
rect 73131 2575 73173 2584
rect 73315 2624 73373 2625
rect 73315 2584 73324 2624
rect 73364 2584 73373 2624
rect 73315 2583 73373 2584
rect 73515 2624 73557 2633
rect 73515 2584 73516 2624
rect 73556 2584 73557 2624
rect 73515 2575 73557 2584
rect 73699 2624 73757 2625
rect 73699 2584 73708 2624
rect 73748 2584 73757 2624
rect 73892 2607 73901 2647
rect 73941 2607 73950 2647
rect 97700 2647 97758 2648
rect 73892 2606 73950 2607
rect 74091 2624 74133 2633
rect 73699 2583 73757 2584
rect 74091 2584 74092 2624
rect 74132 2584 74133 2624
rect 74755 2624 74813 2625
rect 74091 2575 74133 2584
rect 74275 2603 74333 2604
rect 74275 2563 74284 2603
rect 74324 2563 74333 2603
rect 74755 2584 74764 2624
rect 74804 2584 74813 2624
rect 74755 2583 74813 2584
rect 74955 2624 74997 2633
rect 74955 2584 74956 2624
rect 74996 2584 74997 2624
rect 74955 2575 74997 2584
rect 75619 2624 75677 2625
rect 75619 2584 75628 2624
rect 75668 2584 75677 2624
rect 75619 2583 75677 2584
rect 75819 2624 75861 2633
rect 75819 2584 75820 2624
rect 75860 2584 75861 2624
rect 75819 2575 75861 2584
rect 77067 2624 77109 2633
rect 77067 2584 77068 2624
rect 77108 2584 77109 2624
rect 77067 2575 77109 2584
rect 77251 2624 77309 2625
rect 77251 2584 77260 2624
rect 77300 2584 77309 2624
rect 77251 2583 77309 2584
rect 78603 2624 78645 2633
rect 78603 2584 78604 2624
rect 78644 2584 78645 2624
rect 78603 2575 78645 2584
rect 78787 2624 78845 2625
rect 78787 2584 78796 2624
rect 78836 2584 78845 2624
rect 78787 2583 78845 2584
rect 81675 2624 81717 2633
rect 81675 2584 81676 2624
rect 81716 2584 81717 2624
rect 81675 2575 81717 2584
rect 81859 2624 81917 2625
rect 81859 2584 81868 2624
rect 81908 2584 81917 2624
rect 81859 2583 81917 2584
rect 83211 2624 83253 2633
rect 83211 2584 83212 2624
rect 83252 2584 83253 2624
rect 83211 2575 83253 2584
rect 83395 2624 83453 2625
rect 83395 2584 83404 2624
rect 83444 2584 83453 2624
rect 83395 2583 83453 2584
rect 84747 2624 84789 2633
rect 84747 2584 84748 2624
rect 84788 2584 84789 2624
rect 84747 2575 84789 2584
rect 84931 2624 84989 2625
rect 84931 2584 84940 2624
rect 84980 2584 84989 2624
rect 84931 2583 84989 2584
rect 85131 2624 85173 2633
rect 85131 2584 85132 2624
rect 85172 2584 85173 2624
rect 85131 2575 85173 2584
rect 85315 2624 85373 2625
rect 85315 2584 85324 2624
rect 85364 2584 85373 2624
rect 85315 2583 85373 2584
rect 85515 2624 85557 2633
rect 85515 2584 85516 2624
rect 85556 2584 85557 2624
rect 85515 2575 85557 2584
rect 85699 2624 85757 2625
rect 85699 2584 85708 2624
rect 85748 2584 85757 2624
rect 85699 2583 85757 2584
rect 85899 2624 85941 2633
rect 85899 2584 85900 2624
rect 85940 2584 85941 2624
rect 85899 2575 85941 2584
rect 86083 2624 86141 2625
rect 86083 2584 86092 2624
rect 86132 2584 86141 2624
rect 86083 2583 86141 2584
rect 86283 2624 86325 2633
rect 86283 2584 86284 2624
rect 86324 2584 86325 2624
rect 86283 2575 86325 2584
rect 86467 2624 86525 2625
rect 86467 2584 86476 2624
rect 86516 2584 86525 2624
rect 86467 2583 86525 2584
rect 92899 2624 92957 2625
rect 92899 2584 92908 2624
rect 92948 2584 92957 2624
rect 92899 2583 92957 2584
rect 93099 2624 93141 2633
rect 93099 2584 93100 2624
rect 93140 2584 93141 2624
rect 93099 2575 93141 2584
rect 93571 2624 93629 2625
rect 93571 2584 93580 2624
rect 93620 2584 93629 2624
rect 93571 2583 93629 2584
rect 93771 2624 93813 2633
rect 93771 2584 93772 2624
rect 93812 2584 93813 2624
rect 93771 2575 93813 2584
rect 95107 2624 95165 2625
rect 95107 2584 95116 2624
rect 95156 2584 95165 2624
rect 95107 2583 95165 2584
rect 95307 2624 95349 2633
rect 95307 2584 95308 2624
rect 95348 2584 95349 2624
rect 95307 2575 95349 2584
rect 96355 2624 96413 2625
rect 96355 2584 96364 2624
rect 96404 2584 96413 2624
rect 96355 2583 96413 2584
rect 96555 2624 96597 2633
rect 96555 2584 96556 2624
rect 96596 2584 96597 2624
rect 96555 2575 96597 2584
rect 96739 2624 96797 2625
rect 96739 2584 96748 2624
rect 96788 2584 96797 2624
rect 96739 2583 96797 2584
rect 96939 2624 96981 2633
rect 96939 2584 96940 2624
rect 96980 2584 96981 2624
rect 96939 2575 96981 2584
rect 97123 2624 97181 2625
rect 97123 2584 97132 2624
rect 97172 2584 97181 2624
rect 97123 2583 97181 2584
rect 97323 2624 97365 2633
rect 97323 2584 97324 2624
rect 97364 2584 97365 2624
rect 97323 2575 97365 2584
rect 97507 2624 97565 2625
rect 97507 2584 97516 2624
rect 97556 2584 97565 2624
rect 97700 2607 97709 2647
rect 97749 2607 97758 2647
rect 97700 2606 97758 2607
rect 97899 2624 97941 2633
rect 97507 2583 97565 2584
rect 97899 2584 97900 2624
rect 97940 2584 97941 2624
rect 97899 2575 97941 2584
rect 98083 2624 98141 2625
rect 98083 2584 98092 2624
rect 98132 2584 98141 2624
rect 98083 2583 98141 2584
rect 74275 2562 74333 2563
rect 1707 2540 1749 2549
rect 1707 2500 1708 2540
rect 1748 2500 1749 2540
rect 1707 2491 1749 2500
rect 2187 2540 2229 2549
rect 2187 2500 2188 2540
rect 2228 2500 2229 2540
rect 2187 2491 2229 2500
rect 2571 2540 2613 2549
rect 2571 2500 2572 2540
rect 2612 2500 2613 2540
rect 2571 2491 2613 2500
rect 3051 2540 3093 2549
rect 3051 2500 3052 2540
rect 3092 2500 3093 2540
rect 3051 2491 3093 2500
rect 3435 2540 3477 2549
rect 3435 2500 3436 2540
rect 3476 2500 3477 2540
rect 3435 2491 3477 2500
rect 3819 2540 3861 2549
rect 3819 2500 3820 2540
rect 3860 2500 3861 2540
rect 3819 2491 3861 2500
rect 6219 2540 6261 2549
rect 6219 2500 6220 2540
rect 6260 2500 6261 2540
rect 6219 2491 6261 2500
rect 6699 2540 6741 2549
rect 6699 2500 6700 2540
rect 6740 2500 6741 2540
rect 6699 2491 6741 2500
rect 7083 2540 7125 2549
rect 7083 2500 7084 2540
rect 7124 2500 7125 2540
rect 7083 2491 7125 2500
rect 8139 2540 8181 2549
rect 8139 2500 8140 2540
rect 8180 2500 8181 2540
rect 8139 2491 8181 2500
rect 12651 2540 12693 2549
rect 12651 2500 12652 2540
rect 12692 2500 12693 2540
rect 12651 2491 12693 2500
rect 14187 2540 14229 2549
rect 14187 2500 14188 2540
rect 14228 2500 14229 2540
rect 14187 2491 14229 2500
rect 19755 2540 19797 2549
rect 19755 2500 19756 2540
rect 19796 2500 19797 2540
rect 19755 2491 19797 2500
rect 20331 2540 20373 2549
rect 20331 2500 20332 2540
rect 20372 2500 20373 2540
rect 20331 2491 20373 2500
rect 21963 2540 22005 2549
rect 21963 2500 21964 2540
rect 22004 2500 22005 2540
rect 21963 2491 22005 2500
rect 23499 2540 23541 2549
rect 23499 2500 23500 2540
rect 23540 2500 23541 2540
rect 23499 2491 23541 2500
rect 26475 2540 26517 2549
rect 26475 2500 26476 2540
rect 26516 2500 26517 2540
rect 26475 2491 26517 2500
rect 28011 2540 28053 2549
rect 28011 2500 28012 2540
rect 28052 2500 28053 2540
rect 28011 2491 28053 2500
rect 29643 2540 29685 2549
rect 29643 2500 29644 2540
rect 29684 2500 29685 2540
rect 29643 2491 29685 2500
rect 30795 2540 30837 2549
rect 30795 2500 30796 2540
rect 30836 2500 30837 2540
rect 30795 2491 30837 2500
rect 31755 2540 31797 2549
rect 31755 2500 31756 2540
rect 31796 2500 31797 2540
rect 31755 2491 31797 2500
rect 37707 2540 37749 2549
rect 37707 2500 37708 2540
rect 37748 2500 37749 2540
rect 37707 2491 37749 2500
rect 38283 2540 38325 2549
rect 38283 2500 38284 2540
rect 38324 2500 38325 2540
rect 38283 2491 38325 2500
rect 38667 2540 38709 2549
rect 38667 2500 38668 2540
rect 38708 2500 38709 2540
rect 38667 2491 38709 2500
rect 40107 2540 40149 2549
rect 40107 2500 40108 2540
rect 40148 2500 40149 2540
rect 40107 2491 40149 2500
rect 41739 2540 41781 2549
rect 41739 2500 41740 2540
rect 41780 2500 41781 2540
rect 41739 2491 41781 2500
rect 42123 2540 42165 2549
rect 42123 2500 42124 2540
rect 42164 2500 42165 2540
rect 42123 2491 42165 2500
rect 42891 2540 42933 2549
rect 42891 2500 42892 2540
rect 42932 2500 42933 2540
rect 42891 2491 42933 2500
rect 44139 2540 44181 2549
rect 44139 2500 44140 2540
rect 44180 2500 44181 2540
rect 44139 2491 44181 2500
rect 44907 2540 44949 2549
rect 44907 2500 44908 2540
rect 44948 2500 44949 2540
rect 44907 2491 44949 2500
rect 46443 2540 46485 2549
rect 46443 2500 46444 2540
rect 46484 2500 46485 2540
rect 46443 2491 46485 2500
rect 47979 2540 48021 2549
rect 47979 2500 47980 2540
rect 48020 2500 48021 2540
rect 47979 2491 48021 2500
rect 48363 2540 48405 2549
rect 48363 2500 48364 2540
rect 48404 2500 48405 2540
rect 48363 2491 48405 2500
rect 48747 2540 48789 2549
rect 48747 2500 48748 2540
rect 48788 2500 48789 2540
rect 48747 2491 48789 2500
rect 49227 2540 49269 2549
rect 49227 2500 49228 2540
rect 49268 2500 49269 2540
rect 49227 2491 49269 2500
rect 62955 2540 62997 2549
rect 62955 2500 62956 2540
rect 62996 2500 62997 2540
rect 62955 2491 62997 2500
rect 63435 2540 63477 2549
rect 63435 2500 63436 2540
rect 63476 2500 63477 2540
rect 63435 2491 63477 2500
rect 67467 2540 67509 2549
rect 67467 2500 67468 2540
rect 67508 2500 67509 2540
rect 67467 2491 67509 2500
rect 73035 2540 73077 2549
rect 73035 2500 73036 2540
rect 73076 2500 73077 2540
rect 73035 2491 73077 2500
rect 73419 2540 73461 2549
rect 73419 2500 73420 2540
rect 73460 2500 73461 2540
rect 73419 2491 73461 2500
rect 73803 2540 73845 2549
rect 73803 2500 73804 2540
rect 73844 2500 73845 2540
rect 73803 2491 73845 2500
rect 74187 2540 74229 2549
rect 74187 2500 74188 2540
rect 74228 2500 74229 2540
rect 74187 2491 74229 2500
rect 74859 2540 74901 2549
rect 74859 2500 74860 2540
rect 74900 2500 74901 2540
rect 74859 2491 74901 2500
rect 75723 2540 75765 2549
rect 75723 2500 75724 2540
rect 75764 2500 75765 2540
rect 75723 2491 75765 2500
rect 77163 2540 77205 2549
rect 77163 2500 77164 2540
rect 77204 2500 77205 2540
rect 77163 2491 77205 2500
rect 78699 2540 78741 2549
rect 78699 2500 78700 2540
rect 78740 2500 78741 2540
rect 78699 2491 78741 2500
rect 81771 2540 81813 2549
rect 81771 2500 81772 2540
rect 81812 2500 81813 2540
rect 81771 2491 81813 2500
rect 83307 2540 83349 2549
rect 83307 2500 83308 2540
rect 83348 2500 83349 2540
rect 83307 2491 83349 2500
rect 84843 2540 84885 2549
rect 84843 2500 84844 2540
rect 84884 2500 84885 2540
rect 84843 2491 84885 2500
rect 85227 2540 85269 2549
rect 85227 2500 85228 2540
rect 85268 2500 85269 2540
rect 85227 2491 85269 2500
rect 85611 2540 85653 2549
rect 85611 2500 85612 2540
rect 85652 2500 85653 2540
rect 85611 2491 85653 2500
rect 85995 2540 86037 2549
rect 85995 2500 85996 2540
rect 86036 2500 86037 2540
rect 85995 2491 86037 2500
rect 86379 2540 86421 2549
rect 86379 2500 86380 2540
rect 86420 2500 86421 2540
rect 86379 2491 86421 2500
rect 93003 2540 93045 2549
rect 93003 2500 93004 2540
rect 93044 2500 93045 2540
rect 93003 2491 93045 2500
rect 93675 2540 93717 2549
rect 93675 2500 93676 2540
rect 93716 2500 93717 2540
rect 93675 2491 93717 2500
rect 95211 2540 95253 2549
rect 95211 2500 95212 2540
rect 95252 2500 95253 2540
rect 95211 2491 95253 2500
rect 96459 2540 96501 2549
rect 96459 2500 96460 2540
rect 96500 2500 96501 2540
rect 96459 2491 96501 2500
rect 96843 2540 96885 2549
rect 96843 2500 96844 2540
rect 96884 2500 96885 2540
rect 96843 2491 96885 2500
rect 97227 2540 97269 2549
rect 97227 2500 97228 2540
rect 97268 2500 97269 2540
rect 97227 2491 97269 2500
rect 97611 2540 97653 2549
rect 97611 2500 97612 2540
rect 97652 2500 97653 2540
rect 97611 2491 97653 2500
rect 97995 2540 98037 2549
rect 97995 2500 97996 2540
rect 98036 2500 98037 2540
rect 97995 2491 98037 2500
rect 55083 2456 55125 2465
rect 55083 2416 55084 2456
rect 55124 2416 55125 2456
rect 55083 2407 55125 2416
rect 55563 2456 55605 2465
rect 55563 2416 55564 2456
rect 55604 2416 55605 2456
rect 55563 2407 55605 2416
rect 56139 2456 56181 2465
rect 56139 2416 56140 2456
rect 56180 2416 56181 2456
rect 56139 2407 56181 2416
rect 58827 2456 58869 2465
rect 58827 2416 58828 2456
rect 58868 2416 58869 2456
rect 58827 2407 58869 2416
rect 60555 2456 60597 2465
rect 60555 2416 60556 2456
rect 60596 2416 60597 2456
rect 60555 2407 60597 2416
rect 61131 2456 61173 2465
rect 61131 2416 61132 2456
rect 61172 2416 61173 2456
rect 61131 2407 61173 2416
rect 61611 2456 61653 2465
rect 61611 2416 61612 2456
rect 61652 2416 61653 2456
rect 61611 2407 61653 2416
rect 61899 2456 61941 2465
rect 61899 2416 61900 2456
rect 61940 2416 61941 2456
rect 61899 2407 61941 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 98083 1973 98141 1974
rect 1507 1952 1565 1953
rect 1507 1912 1516 1952
rect 1556 1912 1565 1952
rect 1507 1911 1565 1912
rect 1707 1952 1749 1961
rect 1707 1912 1708 1952
rect 1748 1912 1749 1952
rect 1707 1903 1749 1912
rect 5355 1952 5397 1961
rect 5355 1912 5356 1952
rect 5396 1912 5397 1952
rect 5355 1903 5397 1912
rect 5539 1952 5597 1953
rect 5539 1912 5548 1952
rect 5588 1912 5597 1952
rect 5539 1911 5597 1912
rect 6795 1952 6837 1961
rect 6795 1912 6796 1952
rect 6836 1912 6837 1952
rect 6795 1903 6837 1912
rect 6987 1952 7029 1961
rect 6987 1912 6988 1952
rect 7028 1912 7029 1952
rect 6987 1903 7029 1912
rect 19363 1952 19421 1953
rect 19363 1912 19372 1952
rect 19412 1912 19421 1952
rect 19363 1911 19421 1912
rect 19563 1952 19605 1961
rect 19563 1912 19564 1952
rect 19604 1912 19605 1952
rect 19563 1903 19605 1912
rect 24651 1952 24693 1961
rect 24651 1912 24652 1952
rect 24692 1912 24693 1952
rect 24651 1903 24693 1912
rect 24835 1952 24893 1953
rect 24835 1912 24844 1952
rect 24884 1912 24893 1952
rect 24835 1911 24893 1912
rect 25899 1952 25941 1961
rect 25899 1912 25900 1952
rect 25940 1912 25941 1952
rect 25899 1903 25941 1912
rect 26091 1952 26133 1961
rect 26091 1912 26092 1952
rect 26132 1912 26133 1952
rect 26091 1903 26133 1912
rect 31947 1952 31989 1961
rect 31947 1912 31948 1952
rect 31988 1912 31989 1952
rect 31947 1903 31989 1912
rect 32139 1952 32181 1961
rect 32139 1912 32140 1952
rect 32180 1912 32181 1952
rect 32139 1903 32181 1912
rect 43659 1952 43701 1961
rect 43659 1912 43660 1952
rect 43700 1912 43701 1952
rect 43659 1903 43701 1912
rect 43843 1952 43901 1953
rect 43843 1912 43852 1952
rect 43892 1912 43901 1952
rect 43843 1911 43901 1912
rect 51243 1952 51285 1961
rect 51243 1912 51244 1952
rect 51284 1912 51285 1952
rect 51243 1903 51285 1912
rect 51435 1952 51477 1961
rect 51435 1912 51436 1952
rect 51476 1912 51477 1952
rect 51435 1903 51477 1912
rect 51819 1952 51861 1961
rect 51819 1912 51820 1952
rect 51860 1912 51861 1952
rect 51819 1903 51861 1912
rect 52107 1952 52149 1961
rect 52107 1912 52108 1952
rect 52148 1912 52149 1952
rect 52107 1903 52149 1912
rect 52299 1952 52341 1961
rect 52299 1912 52300 1952
rect 52340 1912 52341 1952
rect 52299 1903 52341 1912
rect 52875 1952 52917 1961
rect 52875 1912 52876 1952
rect 52916 1912 52917 1952
rect 52875 1903 52917 1912
rect 53163 1952 53205 1961
rect 53163 1912 53164 1952
rect 53204 1912 53205 1952
rect 53163 1903 53205 1912
rect 53355 1952 53397 1961
rect 53355 1912 53356 1952
rect 53396 1912 53397 1952
rect 53355 1903 53397 1912
rect 54315 1952 54357 1961
rect 54315 1912 54316 1952
rect 54356 1912 54357 1952
rect 54315 1903 54357 1912
rect 54507 1952 54549 1961
rect 54507 1912 54508 1952
rect 54548 1912 54549 1952
rect 54507 1903 54549 1912
rect 57003 1952 57045 1961
rect 57003 1912 57004 1952
rect 57044 1912 57045 1952
rect 57003 1903 57045 1912
rect 57195 1952 57237 1961
rect 57195 1912 57196 1952
rect 57236 1912 57237 1952
rect 57195 1903 57237 1912
rect 57483 1952 57525 1961
rect 57483 1912 57484 1952
rect 57524 1912 57525 1952
rect 57483 1903 57525 1912
rect 57867 1952 57909 1961
rect 57867 1912 57868 1952
rect 57908 1912 57909 1952
rect 57867 1903 57909 1912
rect 58059 1952 58101 1961
rect 58059 1912 58060 1952
rect 58100 1912 58101 1952
rect 58059 1903 58101 1912
rect 58731 1952 58773 1961
rect 58731 1912 58732 1952
rect 58772 1912 58773 1952
rect 58731 1903 58773 1912
rect 58923 1952 58965 1961
rect 58923 1912 58924 1952
rect 58964 1912 58965 1952
rect 58923 1903 58965 1912
rect 59979 1952 60021 1961
rect 59979 1912 59980 1952
rect 60020 1912 60021 1952
rect 59979 1903 60021 1912
rect 60171 1952 60213 1961
rect 60171 1912 60172 1952
rect 60212 1912 60213 1952
rect 60171 1903 60213 1912
rect 62571 1952 62613 1961
rect 62571 1912 62572 1952
rect 62612 1912 62613 1952
rect 62571 1903 62613 1912
rect 62755 1952 62813 1953
rect 62755 1912 62764 1952
rect 62804 1912 62813 1952
rect 62755 1911 62813 1912
rect 64867 1952 64925 1953
rect 64867 1912 64876 1952
rect 64916 1912 64925 1952
rect 64867 1911 64925 1912
rect 65067 1952 65109 1961
rect 65067 1912 65068 1952
rect 65108 1912 65109 1952
rect 65067 1903 65109 1912
rect 66403 1952 66461 1953
rect 66403 1912 66412 1952
rect 66452 1912 66461 1952
rect 66403 1911 66461 1912
rect 66603 1952 66645 1961
rect 66603 1912 66604 1952
rect 66644 1912 66645 1952
rect 66603 1903 66645 1912
rect 67651 1952 67709 1953
rect 67651 1912 67660 1952
rect 67700 1912 67709 1952
rect 67651 1911 67709 1912
rect 67851 1952 67893 1961
rect 67851 1912 67852 1952
rect 67892 1912 67893 1952
rect 67851 1903 67893 1912
rect 79947 1952 79989 1961
rect 79947 1912 79948 1952
rect 79988 1912 79989 1952
rect 79947 1903 79989 1912
rect 80139 1952 80181 1961
rect 80139 1912 80140 1952
rect 80180 1912 80181 1952
rect 80139 1903 80181 1912
rect 80803 1952 80861 1953
rect 80803 1912 80812 1952
rect 80852 1912 80861 1952
rect 80803 1911 80861 1912
rect 81003 1952 81045 1961
rect 81003 1912 81004 1952
rect 81044 1912 81045 1952
rect 81003 1903 81045 1912
rect 92515 1952 92573 1953
rect 92515 1912 92524 1952
rect 92564 1912 92573 1952
rect 92515 1911 92573 1912
rect 92715 1952 92757 1961
rect 92715 1912 92716 1952
rect 92756 1912 92757 1952
rect 92715 1903 92757 1912
rect 97899 1952 97941 1961
rect 97899 1912 97900 1952
rect 97940 1912 97941 1952
rect 98083 1933 98092 1973
rect 98132 1933 98141 1973
rect 98083 1932 98141 1933
rect 97899 1903 97941 1912
rect 25995 1868 26037 1877
rect 25995 1828 25996 1868
rect 26036 1828 26037 1868
rect 25995 1819 26037 1828
rect 51339 1868 51381 1877
rect 51339 1828 51340 1868
rect 51380 1828 51381 1868
rect 51339 1819 51381 1828
rect 60075 1868 60117 1877
rect 60075 1828 60076 1868
rect 60116 1828 60117 1868
rect 60075 1819 60117 1828
rect 51819 1784 51861 1793
rect 51819 1744 51820 1784
rect 51860 1744 51861 1784
rect 51819 1735 51861 1744
rect 52875 1784 52917 1793
rect 52875 1744 52876 1784
rect 52916 1744 52917 1784
rect 52875 1735 52917 1744
rect 57483 1784 57525 1793
rect 57483 1744 57484 1784
rect 57524 1744 57525 1784
rect 57483 1735 57525 1744
rect 1611 1700 1653 1709
rect 1611 1660 1612 1700
rect 1652 1660 1653 1700
rect 1611 1651 1653 1660
rect 5451 1700 5493 1709
rect 5451 1660 5452 1700
rect 5492 1660 5493 1700
rect 5451 1651 5493 1660
rect 6795 1700 6837 1709
rect 6795 1660 6796 1700
rect 6836 1660 6837 1700
rect 6795 1651 6837 1660
rect 19467 1700 19509 1709
rect 19467 1660 19468 1700
rect 19508 1660 19509 1700
rect 19467 1651 19509 1660
rect 24747 1700 24789 1709
rect 24747 1660 24748 1700
rect 24788 1660 24789 1700
rect 24747 1651 24789 1660
rect 31947 1700 31989 1709
rect 31947 1660 31948 1700
rect 31988 1660 31989 1700
rect 31947 1651 31989 1660
rect 43755 1700 43797 1709
rect 43755 1660 43756 1700
rect 43796 1660 43797 1700
rect 43755 1651 43797 1660
rect 51627 1700 51669 1709
rect 51627 1660 51628 1700
rect 51668 1660 51669 1700
rect 51627 1651 51669 1660
rect 52107 1700 52149 1709
rect 52107 1660 52108 1700
rect 52148 1660 52149 1700
rect 52107 1651 52149 1660
rect 52683 1700 52725 1709
rect 52683 1660 52684 1700
rect 52724 1660 52725 1700
rect 52683 1651 52725 1660
rect 53163 1700 53205 1709
rect 53163 1660 53164 1700
rect 53204 1660 53205 1700
rect 53163 1651 53205 1660
rect 54507 1700 54549 1709
rect 54507 1660 54508 1700
rect 54548 1660 54549 1700
rect 54507 1651 54549 1660
rect 57195 1700 57237 1709
rect 57195 1660 57196 1700
rect 57236 1660 57237 1700
rect 57195 1651 57237 1660
rect 57675 1700 57717 1709
rect 57675 1660 57676 1700
rect 57716 1660 57717 1700
rect 57675 1651 57717 1660
rect 57867 1700 57909 1709
rect 57867 1660 57868 1700
rect 57908 1660 57909 1700
rect 57867 1651 57909 1660
rect 58731 1700 58773 1709
rect 58731 1660 58732 1700
rect 58772 1660 58773 1700
rect 58731 1651 58773 1660
rect 62667 1700 62709 1709
rect 62667 1660 62668 1700
rect 62708 1660 62709 1700
rect 62667 1651 62709 1660
rect 64971 1700 65013 1709
rect 64971 1660 64972 1700
rect 65012 1660 65013 1700
rect 64971 1651 65013 1660
rect 66507 1700 66549 1709
rect 66507 1660 66508 1700
rect 66548 1660 66549 1700
rect 66507 1651 66549 1660
rect 67755 1700 67797 1709
rect 67755 1660 67756 1700
rect 67796 1660 67797 1700
rect 67755 1651 67797 1660
rect 80139 1700 80181 1709
rect 80139 1660 80140 1700
rect 80180 1660 80181 1700
rect 80139 1651 80181 1660
rect 80907 1700 80949 1709
rect 80907 1660 80908 1700
rect 80948 1660 80949 1700
rect 80907 1651 80949 1660
rect 92619 1700 92661 1709
rect 92619 1660 92620 1700
rect 92660 1660 92661 1700
rect 92619 1651 92661 1660
rect 97995 1700 98037 1709
rect 97995 1660 97996 1700
rect 98036 1660 98037 1700
rect 97995 1651 98037 1660
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 6987 1364 7029 1373
rect 6987 1324 6988 1364
rect 7028 1324 7029 1364
rect 6987 1315 7029 1324
rect 14283 1364 14325 1373
rect 14283 1324 14284 1364
rect 14324 1324 14325 1364
rect 14283 1315 14325 1324
rect 16587 1364 16629 1373
rect 16587 1324 16588 1364
rect 16628 1324 16629 1364
rect 16587 1315 16629 1324
rect 20427 1364 20469 1373
rect 20427 1324 20428 1364
rect 20468 1324 20469 1364
rect 20427 1315 20469 1324
rect 24651 1364 24693 1373
rect 24651 1324 24652 1364
rect 24692 1324 24693 1364
rect 24651 1315 24693 1324
rect 30699 1364 30741 1373
rect 30699 1324 30700 1364
rect 30740 1324 30741 1364
rect 30699 1315 30741 1324
rect 63051 1364 63093 1373
rect 63051 1324 63052 1364
rect 63092 1324 63093 1364
rect 63051 1315 63093 1324
rect 66891 1364 66933 1373
rect 66891 1324 66892 1364
rect 66932 1324 66933 1364
rect 66891 1315 66933 1324
rect 70731 1364 70773 1373
rect 70731 1324 70732 1364
rect 70772 1324 70773 1364
rect 70731 1315 70773 1324
rect 72267 1364 72309 1373
rect 72267 1324 72268 1364
rect 72308 1324 72309 1364
rect 72267 1315 72309 1324
rect 82827 1364 82869 1373
rect 82827 1324 82828 1364
rect 82868 1324 82869 1364
rect 82827 1315 82869 1324
rect 85515 1364 85557 1373
rect 85515 1324 85516 1364
rect 85556 1324 85557 1364
rect 85515 1315 85557 1324
rect 85899 1364 85941 1373
rect 85899 1324 85900 1364
rect 85940 1324 85941 1364
rect 85899 1315 85941 1324
rect 98379 1364 98421 1373
rect 98379 1324 98380 1364
rect 98420 1324 98421 1364
rect 98379 1315 98421 1324
rect 31659 1280 31701 1289
rect 31659 1240 31660 1280
rect 31700 1240 31701 1280
rect 31659 1231 31701 1240
rect 50955 1280 50997 1289
rect 50955 1240 50956 1280
rect 50996 1240 50997 1280
rect 52203 1280 52245 1289
rect 50955 1231 50997 1240
rect 51435 1254 51477 1263
rect 51435 1214 51436 1254
rect 51476 1214 51477 1254
rect 52203 1240 52204 1280
rect 52244 1240 52245 1280
rect 52203 1231 52245 1240
rect 54123 1280 54165 1289
rect 54123 1240 54124 1280
rect 54164 1240 54165 1280
rect 54123 1231 54165 1240
rect 54603 1280 54645 1289
rect 54603 1240 54604 1280
rect 54644 1240 54645 1280
rect 54603 1231 54645 1240
rect 55083 1280 55125 1289
rect 55083 1240 55084 1280
rect 55124 1240 55125 1280
rect 55083 1231 55125 1240
rect 56715 1280 56757 1289
rect 56715 1240 56716 1280
rect 56756 1240 56757 1280
rect 56715 1231 56757 1240
rect 57195 1280 57237 1289
rect 57195 1240 57196 1280
rect 57236 1240 57237 1280
rect 57195 1231 57237 1240
rect 57771 1280 57813 1289
rect 57771 1240 57772 1280
rect 57812 1240 57813 1280
rect 57771 1231 57813 1240
rect 59307 1280 59349 1289
rect 59307 1240 59308 1280
rect 59348 1240 59349 1280
rect 59307 1231 59349 1240
rect 59595 1280 59637 1289
rect 59595 1240 59596 1280
rect 59636 1240 59637 1280
rect 59595 1231 59637 1240
rect 60171 1280 60213 1289
rect 60171 1240 60172 1280
rect 60212 1240 60213 1280
rect 60171 1231 60213 1240
rect 60651 1280 60693 1289
rect 60651 1240 60652 1280
rect 60692 1240 60693 1280
rect 60651 1231 60693 1240
rect 51435 1205 51477 1214
rect 66603 1196 66645 1205
rect 66603 1156 66604 1196
rect 66644 1156 66645 1196
rect 66603 1147 66645 1156
rect 4107 1125 4149 1134
rect 1035 1112 1077 1121
rect 1035 1072 1036 1112
rect 1076 1072 1077 1112
rect 1035 1063 1077 1072
rect 1227 1112 1269 1121
rect 1227 1072 1228 1112
rect 1268 1072 1269 1112
rect 1227 1063 1269 1072
rect 1419 1112 1461 1121
rect 1419 1072 1420 1112
rect 1460 1072 1461 1112
rect 1419 1063 1461 1072
rect 1611 1112 1653 1121
rect 1611 1072 1612 1112
rect 1652 1072 1653 1112
rect 1611 1063 1653 1072
rect 1803 1112 1845 1121
rect 1803 1072 1804 1112
rect 1844 1072 1845 1112
rect 1803 1063 1845 1072
rect 1995 1112 2037 1121
rect 1995 1072 1996 1112
rect 2036 1072 2037 1112
rect 1995 1063 2037 1072
rect 2187 1112 2229 1121
rect 2187 1072 2188 1112
rect 2228 1072 2229 1112
rect 2187 1063 2229 1072
rect 2379 1112 2421 1121
rect 2379 1072 2380 1112
rect 2420 1072 2421 1112
rect 2379 1063 2421 1072
rect 2571 1112 2613 1121
rect 2571 1072 2572 1112
rect 2612 1072 2613 1112
rect 2571 1063 2613 1072
rect 2763 1112 2805 1121
rect 2763 1072 2764 1112
rect 2804 1072 2805 1112
rect 2763 1063 2805 1072
rect 2955 1112 2997 1121
rect 2955 1072 2956 1112
rect 2996 1072 2997 1112
rect 2955 1063 2997 1072
rect 3147 1112 3189 1121
rect 3147 1072 3148 1112
rect 3188 1072 3189 1112
rect 3147 1063 3189 1072
rect 3339 1112 3381 1121
rect 3339 1072 3340 1112
rect 3380 1072 3381 1112
rect 3339 1063 3381 1072
rect 3531 1112 3573 1121
rect 3531 1072 3532 1112
rect 3572 1072 3573 1112
rect 3531 1063 3573 1072
rect 3723 1112 3765 1121
rect 3723 1072 3724 1112
rect 3764 1072 3765 1112
rect 3723 1063 3765 1072
rect 3915 1112 3957 1121
rect 3915 1072 3916 1112
rect 3956 1072 3957 1112
rect 4107 1085 4108 1125
rect 4148 1085 4149 1125
rect 4484 1125 4542 1126
rect 4107 1076 4149 1085
rect 4299 1112 4341 1121
rect 3915 1063 3957 1072
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4484 1085 4493 1125
rect 4533 1085 4542 1125
rect 6994 1125 7036 1134
rect 4484 1084 4542 1085
rect 4683 1112 4725 1121
rect 4299 1063 4341 1072
rect 4683 1072 4684 1112
rect 4724 1072 4725 1112
rect 4683 1063 4725 1072
rect 4875 1112 4917 1121
rect 4875 1072 4876 1112
rect 4916 1072 4917 1112
rect 4875 1063 4917 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5259 1112 5301 1121
rect 5259 1072 5260 1112
rect 5300 1072 5301 1112
rect 5259 1063 5301 1072
rect 5451 1112 5493 1121
rect 5451 1072 5452 1112
rect 5492 1072 5493 1112
rect 5451 1063 5493 1072
rect 5643 1112 5685 1121
rect 5643 1072 5644 1112
rect 5684 1072 5685 1112
rect 5643 1063 5685 1072
rect 5835 1112 5877 1121
rect 5835 1072 5836 1112
rect 5876 1072 5877 1112
rect 6411 1112 6453 1121
rect 5835 1063 5877 1072
rect 6029 1101 6087 1102
rect 6029 1061 6038 1101
rect 6078 1061 6087 1101
rect 6029 1060 6087 1061
rect 6208 1101 6266 1102
rect 6208 1061 6217 1101
rect 6257 1061 6266 1101
rect 6411 1072 6412 1112
rect 6452 1072 6453 1112
rect 6411 1063 6453 1072
rect 6603 1112 6645 1121
rect 6603 1072 6604 1112
rect 6644 1072 6645 1112
rect 6603 1063 6645 1072
rect 6798 1101 6856 1102
rect 6208 1060 6266 1061
rect 6798 1061 6807 1101
rect 6847 1061 6856 1101
rect 6994 1085 6995 1125
rect 7035 1085 7036 1125
rect 11595 1125 11637 1134
rect 6994 1076 7036 1085
rect 7179 1112 7221 1121
rect 7179 1072 7180 1112
rect 7220 1072 7221 1112
rect 7179 1063 7221 1072
rect 7371 1112 7413 1121
rect 7371 1072 7372 1112
rect 7412 1072 7413 1112
rect 7371 1063 7413 1072
rect 7563 1112 7605 1121
rect 7563 1072 7564 1112
rect 7604 1072 7605 1112
rect 7563 1063 7605 1072
rect 7755 1112 7797 1121
rect 7755 1072 7756 1112
rect 7796 1072 7797 1112
rect 7755 1063 7797 1072
rect 7947 1112 7989 1121
rect 7947 1072 7948 1112
rect 7988 1072 7989 1112
rect 7947 1063 7989 1072
rect 8139 1112 8181 1121
rect 8139 1072 8140 1112
rect 8180 1072 8181 1112
rect 8139 1063 8181 1072
rect 8331 1112 8373 1121
rect 8331 1072 8332 1112
rect 8372 1072 8373 1112
rect 8331 1063 8373 1072
rect 8523 1112 8565 1121
rect 8523 1072 8524 1112
rect 8564 1072 8565 1112
rect 8523 1063 8565 1072
rect 8715 1112 8757 1121
rect 8715 1072 8716 1112
rect 8756 1072 8757 1112
rect 8715 1063 8757 1072
rect 8907 1112 8949 1121
rect 8907 1072 8908 1112
rect 8948 1072 8949 1112
rect 8907 1063 8949 1072
rect 9099 1112 9141 1121
rect 9099 1072 9100 1112
rect 9140 1072 9141 1112
rect 9099 1063 9141 1072
rect 9291 1112 9333 1121
rect 9291 1072 9292 1112
rect 9332 1072 9333 1112
rect 9291 1063 9333 1072
rect 9483 1112 9525 1121
rect 9483 1072 9484 1112
rect 9524 1072 9525 1112
rect 9483 1063 9525 1072
rect 9675 1112 9717 1121
rect 9675 1072 9676 1112
rect 9716 1072 9717 1112
rect 9675 1063 9717 1072
rect 9867 1112 9909 1121
rect 9867 1072 9868 1112
rect 9908 1072 9909 1112
rect 9867 1063 9909 1072
rect 10059 1112 10101 1121
rect 10059 1072 10060 1112
rect 10100 1072 10101 1112
rect 10059 1063 10101 1072
rect 10251 1112 10293 1121
rect 10251 1072 10252 1112
rect 10292 1072 10293 1112
rect 10251 1063 10293 1072
rect 10443 1112 10485 1121
rect 10443 1072 10444 1112
rect 10484 1072 10485 1112
rect 10443 1063 10485 1072
rect 10635 1112 10677 1121
rect 10635 1072 10636 1112
rect 10676 1072 10677 1112
rect 10635 1063 10677 1072
rect 10827 1112 10869 1121
rect 10827 1072 10828 1112
rect 10868 1072 10869 1112
rect 10827 1063 10869 1072
rect 11019 1112 11061 1121
rect 11019 1072 11020 1112
rect 11060 1072 11061 1112
rect 11019 1063 11061 1072
rect 11211 1112 11253 1121
rect 11211 1072 11212 1112
rect 11252 1072 11253 1112
rect 11211 1063 11253 1072
rect 11403 1112 11445 1121
rect 11403 1072 11404 1112
rect 11444 1072 11445 1112
rect 11595 1085 11596 1125
rect 11636 1085 11637 1125
rect 16587 1125 16629 1134
rect 11595 1076 11637 1085
rect 11787 1112 11829 1121
rect 11403 1063 11445 1072
rect 11787 1072 11788 1112
rect 11828 1072 11829 1112
rect 11787 1063 11829 1072
rect 11979 1112 12021 1121
rect 11979 1072 11980 1112
rect 12020 1072 12021 1112
rect 11979 1063 12021 1072
rect 12171 1112 12213 1121
rect 12171 1072 12172 1112
rect 12212 1072 12213 1112
rect 12171 1063 12213 1072
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12747 1109 12789 1118
rect 12747 1069 12748 1109
rect 12788 1069 12789 1109
rect 6798 1060 6856 1061
rect 12747 1060 12789 1069
rect 12939 1112 12981 1121
rect 12939 1072 12940 1112
rect 12980 1072 12981 1112
rect 12939 1063 12981 1072
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 13131 1063 13173 1072
rect 13323 1112 13365 1121
rect 13323 1072 13324 1112
rect 13364 1072 13365 1112
rect 13323 1063 13365 1072
rect 13515 1112 13557 1121
rect 13515 1072 13516 1112
rect 13556 1072 13557 1112
rect 13515 1063 13557 1072
rect 13707 1112 13749 1121
rect 13707 1072 13708 1112
rect 13748 1072 13749 1112
rect 13707 1063 13749 1072
rect 13899 1112 13941 1121
rect 13899 1072 13900 1112
rect 13940 1072 13941 1112
rect 13899 1063 13941 1072
rect 14091 1112 14133 1121
rect 14091 1072 14092 1112
rect 14132 1072 14133 1112
rect 14091 1063 14133 1072
rect 14283 1112 14325 1121
rect 14283 1072 14284 1112
rect 14324 1072 14325 1112
rect 14283 1063 14325 1072
rect 14475 1112 14517 1121
rect 14475 1072 14476 1112
rect 14516 1072 14517 1112
rect 14475 1063 14517 1072
rect 14667 1112 14709 1121
rect 14667 1072 14668 1112
rect 14708 1072 14709 1112
rect 14667 1063 14709 1072
rect 14859 1112 14901 1121
rect 14859 1072 14860 1112
rect 14900 1072 14901 1112
rect 14859 1063 14901 1072
rect 15051 1112 15093 1121
rect 15051 1072 15052 1112
rect 15092 1072 15093 1112
rect 15051 1063 15093 1072
rect 15243 1112 15285 1121
rect 15243 1072 15244 1112
rect 15284 1072 15285 1112
rect 15243 1063 15285 1072
rect 15435 1112 15477 1121
rect 15435 1072 15436 1112
rect 15476 1072 15477 1112
rect 15435 1063 15477 1072
rect 15627 1112 15669 1121
rect 15627 1072 15628 1112
rect 15668 1072 15669 1112
rect 15627 1063 15669 1072
rect 15819 1112 15861 1121
rect 15819 1072 15820 1112
rect 15860 1072 15861 1112
rect 15819 1063 15861 1072
rect 16011 1112 16053 1121
rect 16011 1072 16012 1112
rect 16052 1072 16053 1112
rect 16011 1063 16053 1072
rect 16203 1112 16245 1121
rect 16203 1072 16204 1112
rect 16244 1072 16245 1112
rect 16203 1063 16245 1072
rect 16395 1112 16437 1121
rect 16395 1072 16396 1112
rect 16436 1072 16437 1112
rect 16587 1085 16588 1125
rect 16628 1085 16629 1125
rect 16587 1076 16629 1085
rect 16779 1125 16821 1134
rect 16779 1085 16780 1125
rect 16820 1085 16821 1125
rect 19275 1125 19317 1134
rect 16779 1076 16821 1085
rect 16971 1112 17013 1121
rect 16395 1063 16437 1072
rect 16971 1072 16972 1112
rect 17012 1072 17013 1112
rect 16971 1063 17013 1072
rect 17163 1112 17205 1121
rect 17163 1072 17164 1112
rect 17204 1072 17205 1112
rect 17163 1063 17205 1072
rect 17355 1112 17397 1121
rect 17355 1072 17356 1112
rect 17396 1072 17397 1112
rect 17355 1063 17397 1072
rect 17547 1112 17589 1121
rect 17547 1072 17548 1112
rect 17588 1072 17589 1112
rect 17547 1063 17589 1072
rect 17739 1112 17781 1121
rect 17739 1072 17740 1112
rect 17780 1072 17781 1112
rect 17739 1063 17781 1072
rect 17931 1112 17973 1121
rect 17931 1072 17932 1112
rect 17972 1072 17973 1112
rect 18315 1112 18357 1121
rect 17931 1063 17973 1072
rect 18105 1109 18163 1110
rect 18105 1069 18114 1109
rect 18154 1069 18163 1109
rect 18105 1068 18163 1069
rect 18315 1072 18316 1112
rect 18356 1072 18357 1112
rect 18315 1063 18357 1072
rect 18507 1112 18549 1121
rect 18507 1072 18508 1112
rect 18548 1072 18549 1112
rect 18507 1063 18549 1072
rect 18699 1112 18741 1121
rect 18699 1072 18700 1112
rect 18740 1072 18741 1112
rect 18699 1063 18741 1072
rect 18891 1112 18933 1121
rect 18891 1072 18892 1112
rect 18932 1072 18933 1112
rect 18891 1063 18933 1072
rect 19083 1112 19125 1121
rect 19083 1072 19084 1112
rect 19124 1072 19125 1112
rect 19275 1085 19276 1125
rect 19316 1085 19317 1125
rect 21579 1125 21621 1134
rect 19275 1076 19317 1085
rect 19467 1112 19509 1121
rect 19083 1063 19125 1072
rect 19467 1072 19468 1112
rect 19508 1072 19509 1112
rect 19467 1063 19509 1072
rect 19659 1112 19701 1121
rect 19659 1072 19660 1112
rect 19700 1072 19701 1112
rect 19659 1063 19701 1072
rect 19851 1112 19893 1121
rect 19851 1072 19852 1112
rect 19892 1072 19893 1112
rect 19851 1063 19893 1072
rect 20043 1112 20085 1121
rect 20043 1072 20044 1112
rect 20084 1072 20085 1112
rect 20043 1063 20085 1072
rect 20235 1112 20277 1121
rect 20235 1072 20236 1112
rect 20276 1072 20277 1112
rect 20235 1063 20277 1072
rect 20427 1112 20469 1121
rect 20427 1072 20428 1112
rect 20468 1072 20469 1112
rect 20811 1112 20853 1121
rect 20427 1063 20469 1072
rect 20619 1101 20661 1110
rect 20619 1061 20620 1101
rect 20660 1061 20661 1101
rect 20811 1072 20812 1112
rect 20852 1072 20853 1112
rect 20811 1063 20853 1072
rect 21003 1112 21045 1121
rect 21003 1072 21004 1112
rect 21044 1072 21045 1112
rect 21003 1063 21045 1072
rect 21195 1112 21237 1121
rect 21195 1072 21196 1112
rect 21236 1072 21237 1112
rect 21195 1063 21237 1072
rect 21387 1112 21429 1121
rect 21387 1072 21388 1112
rect 21428 1072 21429 1112
rect 21579 1085 21580 1125
rect 21620 1085 21621 1125
rect 32235 1125 32277 1134
rect 21579 1076 21621 1085
rect 21771 1112 21813 1121
rect 21387 1063 21429 1072
rect 21771 1072 21772 1112
rect 21812 1072 21813 1112
rect 21771 1063 21813 1072
rect 21963 1112 22005 1121
rect 21963 1072 21964 1112
rect 22004 1072 22005 1112
rect 21963 1063 22005 1072
rect 22155 1112 22197 1121
rect 22155 1072 22156 1112
rect 22196 1072 22197 1112
rect 22155 1063 22197 1072
rect 22347 1112 22389 1121
rect 22347 1072 22348 1112
rect 22388 1072 22389 1112
rect 22347 1063 22389 1072
rect 22539 1112 22581 1121
rect 22539 1072 22540 1112
rect 22580 1072 22581 1112
rect 22539 1063 22581 1072
rect 22731 1112 22773 1121
rect 22731 1072 22732 1112
rect 22772 1072 22773 1112
rect 22731 1063 22773 1072
rect 22923 1112 22965 1121
rect 22923 1072 22924 1112
rect 22964 1072 22965 1112
rect 22923 1063 22965 1072
rect 23115 1112 23157 1121
rect 23115 1072 23116 1112
rect 23156 1072 23157 1112
rect 23115 1063 23157 1072
rect 23307 1112 23349 1121
rect 23307 1072 23308 1112
rect 23348 1072 23349 1112
rect 23307 1063 23349 1072
rect 23499 1112 23541 1121
rect 23499 1072 23500 1112
rect 23540 1072 23541 1112
rect 23499 1063 23541 1072
rect 23691 1112 23733 1121
rect 23691 1072 23692 1112
rect 23732 1072 23733 1112
rect 23691 1063 23733 1072
rect 23883 1112 23925 1121
rect 23883 1072 23884 1112
rect 23924 1072 23925 1112
rect 23883 1063 23925 1072
rect 24075 1112 24117 1121
rect 24075 1072 24076 1112
rect 24116 1072 24117 1112
rect 24075 1063 24117 1072
rect 24267 1112 24309 1121
rect 24267 1072 24268 1112
rect 24308 1072 24309 1112
rect 24267 1063 24309 1072
rect 24459 1112 24501 1121
rect 24459 1072 24460 1112
rect 24500 1072 24501 1112
rect 24459 1063 24501 1072
rect 24651 1112 24693 1121
rect 24651 1072 24652 1112
rect 24692 1072 24693 1112
rect 24651 1063 24693 1072
rect 24843 1112 24885 1121
rect 24843 1072 24844 1112
rect 24884 1072 24885 1112
rect 24843 1063 24885 1072
rect 25035 1112 25077 1121
rect 25035 1072 25036 1112
rect 25076 1072 25077 1112
rect 25035 1063 25077 1072
rect 25515 1112 25557 1121
rect 25515 1072 25516 1112
rect 25556 1072 25557 1112
rect 25515 1063 25557 1072
rect 25707 1112 25749 1121
rect 25707 1072 25708 1112
rect 25748 1072 25749 1112
rect 25707 1063 25749 1072
rect 25899 1112 25941 1121
rect 25899 1072 25900 1112
rect 25940 1072 25941 1112
rect 25899 1063 25941 1072
rect 26091 1112 26133 1121
rect 26091 1072 26092 1112
rect 26132 1072 26133 1112
rect 26091 1063 26133 1072
rect 26283 1112 26325 1121
rect 26283 1072 26284 1112
rect 26324 1072 26325 1112
rect 26283 1063 26325 1072
rect 26475 1112 26517 1121
rect 26475 1072 26476 1112
rect 26516 1072 26517 1112
rect 26475 1063 26517 1072
rect 26667 1112 26709 1121
rect 26667 1072 26668 1112
rect 26708 1072 26709 1112
rect 26667 1063 26709 1072
rect 26859 1112 26901 1121
rect 26859 1072 26860 1112
rect 26900 1072 26901 1112
rect 26859 1063 26901 1072
rect 27051 1112 27093 1121
rect 27051 1072 27052 1112
rect 27092 1072 27093 1112
rect 27051 1063 27093 1072
rect 27243 1112 27285 1121
rect 27243 1072 27244 1112
rect 27284 1072 27285 1112
rect 27243 1063 27285 1072
rect 27435 1112 27477 1121
rect 27435 1072 27436 1112
rect 27476 1072 27477 1112
rect 27435 1063 27477 1072
rect 27627 1112 27669 1121
rect 27627 1072 27628 1112
rect 27668 1072 27669 1112
rect 27627 1063 27669 1072
rect 27819 1112 27861 1121
rect 27819 1072 27820 1112
rect 27860 1072 27861 1112
rect 27819 1063 27861 1072
rect 28011 1112 28053 1121
rect 28011 1072 28012 1112
rect 28052 1072 28053 1112
rect 28011 1063 28053 1072
rect 28203 1112 28245 1121
rect 28203 1072 28204 1112
rect 28244 1072 28245 1112
rect 28203 1063 28245 1072
rect 28395 1112 28437 1121
rect 28395 1072 28396 1112
rect 28436 1072 28437 1112
rect 28395 1063 28437 1072
rect 28587 1112 28629 1121
rect 28587 1072 28588 1112
rect 28628 1072 28629 1112
rect 28587 1063 28629 1072
rect 28779 1112 28821 1121
rect 28779 1072 28780 1112
rect 28820 1072 28821 1112
rect 28779 1063 28821 1072
rect 28971 1112 29013 1121
rect 28971 1072 28972 1112
rect 29012 1072 29013 1112
rect 28971 1063 29013 1072
rect 29163 1112 29205 1121
rect 29163 1072 29164 1112
rect 29204 1072 29205 1112
rect 29163 1063 29205 1072
rect 29355 1112 29397 1121
rect 29355 1072 29356 1112
rect 29396 1072 29397 1112
rect 29355 1063 29397 1072
rect 29547 1112 29589 1121
rect 29547 1072 29548 1112
rect 29588 1072 29589 1112
rect 29547 1063 29589 1072
rect 29739 1112 29781 1121
rect 29739 1072 29740 1112
rect 29780 1072 29781 1112
rect 29739 1063 29781 1072
rect 29931 1112 29973 1121
rect 29931 1072 29932 1112
rect 29972 1072 29973 1112
rect 29931 1063 29973 1072
rect 30123 1112 30165 1121
rect 30123 1072 30124 1112
rect 30164 1072 30165 1112
rect 30123 1063 30165 1072
rect 30315 1112 30357 1121
rect 30315 1072 30316 1112
rect 30356 1072 30357 1112
rect 30315 1063 30357 1072
rect 30507 1112 30549 1121
rect 30507 1072 30508 1112
rect 30548 1072 30549 1112
rect 30507 1063 30549 1072
rect 30699 1112 30741 1121
rect 30699 1072 30700 1112
rect 30740 1072 30741 1112
rect 30699 1063 30741 1072
rect 30891 1112 30933 1121
rect 30891 1072 30892 1112
rect 30932 1072 30933 1112
rect 30891 1063 30933 1072
rect 31083 1112 31125 1121
rect 31083 1072 31084 1112
rect 31124 1072 31125 1112
rect 31083 1063 31125 1072
rect 31467 1112 31509 1121
rect 31467 1072 31468 1112
rect 31508 1072 31509 1112
rect 31467 1063 31509 1072
rect 31659 1112 31701 1121
rect 31659 1072 31660 1112
rect 31700 1072 31701 1112
rect 31659 1063 31701 1072
rect 31851 1112 31893 1121
rect 31851 1072 31852 1112
rect 31892 1072 31893 1112
rect 31851 1063 31893 1072
rect 32043 1112 32085 1121
rect 32043 1072 32044 1112
rect 32084 1072 32085 1112
rect 32235 1085 32236 1125
rect 32276 1085 32277 1125
rect 34155 1125 34197 1134
rect 32235 1076 32277 1085
rect 32427 1112 32469 1121
rect 32043 1063 32085 1072
rect 32427 1072 32428 1112
rect 32468 1072 32469 1112
rect 32427 1063 32469 1072
rect 32619 1112 32661 1121
rect 32619 1072 32620 1112
rect 32660 1072 32661 1112
rect 32619 1063 32661 1072
rect 32811 1112 32853 1121
rect 32811 1072 32812 1112
rect 32852 1072 32853 1112
rect 33195 1112 33237 1121
rect 32811 1063 32853 1072
rect 33003 1101 33045 1110
rect 20619 1052 20661 1061
rect 33003 1061 33004 1101
rect 33044 1061 33045 1101
rect 33195 1072 33196 1112
rect 33236 1072 33237 1112
rect 33195 1063 33237 1072
rect 33387 1112 33429 1121
rect 33387 1072 33388 1112
rect 33428 1072 33429 1112
rect 33387 1063 33429 1072
rect 33579 1112 33621 1121
rect 33579 1072 33580 1112
rect 33620 1072 33621 1112
rect 33579 1063 33621 1072
rect 33771 1112 33813 1121
rect 33771 1072 33772 1112
rect 33812 1072 33813 1112
rect 33771 1063 33813 1072
rect 33963 1112 34005 1121
rect 33963 1072 33964 1112
rect 34004 1072 34005 1112
rect 34155 1085 34156 1125
rect 34196 1085 34197 1125
rect 35115 1125 35157 1134
rect 34155 1076 34197 1085
rect 34347 1112 34389 1121
rect 33963 1063 34005 1072
rect 34347 1072 34348 1112
rect 34388 1072 34389 1112
rect 34347 1063 34389 1072
rect 34539 1112 34581 1121
rect 34539 1072 34540 1112
rect 34580 1072 34581 1112
rect 34539 1063 34581 1072
rect 34731 1112 34773 1121
rect 34731 1072 34732 1112
rect 34772 1072 34773 1112
rect 34731 1063 34773 1072
rect 34923 1112 34965 1121
rect 34923 1072 34924 1112
rect 34964 1072 34965 1112
rect 35115 1085 35116 1125
rect 35156 1085 35157 1125
rect 44334 1125 44392 1126
rect 35115 1076 35157 1085
rect 35307 1112 35349 1121
rect 34923 1063 34965 1072
rect 35307 1072 35308 1112
rect 35348 1072 35349 1112
rect 35307 1063 35349 1072
rect 35499 1112 35541 1121
rect 35499 1072 35500 1112
rect 35540 1072 35541 1112
rect 35499 1063 35541 1072
rect 35691 1112 35733 1121
rect 35691 1072 35692 1112
rect 35732 1072 35733 1112
rect 35691 1063 35733 1072
rect 35883 1112 35925 1121
rect 35883 1072 35884 1112
rect 35924 1072 35925 1112
rect 35883 1063 35925 1072
rect 36075 1112 36117 1121
rect 36075 1072 36076 1112
rect 36116 1072 36117 1112
rect 36075 1063 36117 1072
rect 36267 1112 36309 1121
rect 36267 1072 36268 1112
rect 36308 1072 36309 1112
rect 36267 1063 36309 1072
rect 36459 1112 36501 1121
rect 36459 1072 36460 1112
rect 36500 1072 36501 1112
rect 36459 1063 36501 1072
rect 36651 1112 36693 1121
rect 36651 1072 36652 1112
rect 36692 1072 36693 1112
rect 36651 1063 36693 1072
rect 36843 1112 36885 1121
rect 36843 1072 36844 1112
rect 36884 1072 36885 1112
rect 36843 1063 36885 1072
rect 37035 1112 37077 1121
rect 37035 1072 37036 1112
rect 37076 1072 37077 1112
rect 37035 1063 37077 1072
rect 37323 1112 37365 1121
rect 37323 1072 37324 1112
rect 37364 1072 37365 1112
rect 37323 1063 37365 1072
rect 37515 1112 37557 1121
rect 37515 1072 37516 1112
rect 37556 1072 37557 1112
rect 37515 1063 37557 1072
rect 37707 1112 37749 1121
rect 37707 1072 37708 1112
rect 37748 1072 37749 1112
rect 37707 1063 37749 1072
rect 37899 1112 37941 1121
rect 37899 1072 37900 1112
rect 37940 1072 37941 1112
rect 37899 1063 37941 1072
rect 38091 1112 38133 1121
rect 38091 1072 38092 1112
rect 38132 1072 38133 1112
rect 38091 1063 38133 1072
rect 38283 1112 38325 1121
rect 38283 1072 38284 1112
rect 38324 1072 38325 1112
rect 38283 1063 38325 1072
rect 38475 1112 38517 1121
rect 38475 1072 38476 1112
rect 38516 1072 38517 1112
rect 38475 1063 38517 1072
rect 38667 1112 38709 1121
rect 38667 1072 38668 1112
rect 38708 1072 38709 1112
rect 38667 1063 38709 1072
rect 38859 1112 38901 1121
rect 38859 1072 38860 1112
rect 38900 1072 38901 1112
rect 38859 1063 38901 1072
rect 39051 1112 39093 1121
rect 39051 1072 39052 1112
rect 39092 1072 39093 1112
rect 39051 1063 39093 1072
rect 39243 1112 39285 1121
rect 39243 1072 39244 1112
rect 39284 1072 39285 1112
rect 39243 1063 39285 1072
rect 39435 1112 39477 1121
rect 39435 1072 39436 1112
rect 39476 1072 39477 1112
rect 39435 1063 39477 1072
rect 39627 1112 39669 1121
rect 39627 1072 39628 1112
rect 39668 1072 39669 1112
rect 39627 1063 39669 1072
rect 39819 1112 39861 1121
rect 39819 1072 39820 1112
rect 39860 1072 39861 1112
rect 39819 1063 39861 1072
rect 40011 1112 40053 1121
rect 40011 1072 40012 1112
rect 40052 1072 40053 1112
rect 40011 1063 40053 1072
rect 40203 1112 40245 1121
rect 40203 1072 40204 1112
rect 40244 1072 40245 1112
rect 40203 1063 40245 1072
rect 40395 1112 40437 1121
rect 40395 1072 40396 1112
rect 40436 1072 40437 1112
rect 40395 1063 40437 1072
rect 40587 1112 40629 1121
rect 40587 1072 40588 1112
rect 40628 1072 40629 1112
rect 40587 1063 40629 1072
rect 40779 1112 40821 1121
rect 40779 1072 40780 1112
rect 40820 1072 40821 1112
rect 40779 1063 40821 1072
rect 40971 1112 41013 1121
rect 40971 1072 40972 1112
rect 41012 1072 41013 1112
rect 40971 1063 41013 1072
rect 41163 1112 41205 1121
rect 41163 1072 41164 1112
rect 41204 1072 41205 1112
rect 41163 1063 41205 1072
rect 41355 1112 41397 1121
rect 41355 1072 41356 1112
rect 41396 1072 41397 1112
rect 41355 1063 41397 1072
rect 41547 1112 41589 1121
rect 41547 1072 41548 1112
rect 41588 1072 41589 1112
rect 41547 1063 41589 1072
rect 41739 1112 41781 1121
rect 41739 1072 41740 1112
rect 41780 1072 41781 1112
rect 42123 1112 42165 1121
rect 41739 1063 41781 1072
rect 41934 1101 41992 1102
rect 33003 1052 33045 1061
rect 41934 1061 41943 1101
rect 41983 1061 41992 1101
rect 42123 1072 42124 1112
rect 42164 1072 42165 1112
rect 42123 1063 42165 1072
rect 42315 1112 42357 1121
rect 42315 1072 42316 1112
rect 42356 1072 42357 1112
rect 42315 1063 42357 1072
rect 42507 1112 42549 1121
rect 42507 1072 42508 1112
rect 42548 1072 42549 1112
rect 42507 1063 42549 1072
rect 42699 1112 42741 1121
rect 42699 1072 42700 1112
rect 42740 1072 42741 1112
rect 42699 1063 42741 1072
rect 42891 1112 42933 1121
rect 42891 1072 42892 1112
rect 42932 1072 42933 1112
rect 42891 1063 42933 1072
rect 43083 1112 43125 1121
rect 43083 1072 43084 1112
rect 43124 1072 43125 1112
rect 43083 1063 43125 1072
rect 43275 1112 43317 1121
rect 43275 1072 43276 1112
rect 43316 1072 43317 1112
rect 43275 1063 43317 1072
rect 43563 1112 43605 1121
rect 43563 1072 43564 1112
rect 43604 1072 43605 1112
rect 43563 1063 43605 1072
rect 43755 1112 43797 1121
rect 43755 1072 43756 1112
rect 43796 1072 43797 1112
rect 43755 1063 43797 1072
rect 43947 1112 43989 1121
rect 43947 1072 43948 1112
rect 43988 1072 43989 1112
rect 43947 1063 43989 1072
rect 44139 1112 44181 1121
rect 44139 1072 44140 1112
rect 44180 1072 44181 1112
rect 44334 1085 44343 1125
rect 44383 1085 44392 1125
rect 54603 1124 54645 1133
rect 63819 1125 63861 1134
rect 44334 1084 44392 1085
rect 44523 1112 44565 1121
rect 44139 1063 44181 1072
rect 44523 1072 44524 1112
rect 44564 1072 44565 1112
rect 44523 1063 44565 1072
rect 44715 1112 44757 1121
rect 44715 1072 44716 1112
rect 44756 1072 44757 1112
rect 44715 1063 44757 1072
rect 44907 1112 44949 1121
rect 44907 1072 44908 1112
rect 44948 1072 44949 1112
rect 44907 1063 44949 1072
rect 45099 1112 45141 1121
rect 45099 1072 45100 1112
rect 45140 1072 45141 1112
rect 45099 1063 45141 1072
rect 45291 1112 45333 1121
rect 45291 1072 45292 1112
rect 45332 1072 45333 1112
rect 45291 1063 45333 1072
rect 45483 1112 45525 1121
rect 45483 1072 45484 1112
rect 45524 1072 45525 1112
rect 45483 1063 45525 1072
rect 45675 1112 45717 1121
rect 45675 1072 45676 1112
rect 45716 1072 45717 1112
rect 45675 1063 45717 1072
rect 45867 1112 45909 1121
rect 45867 1072 45868 1112
rect 45908 1072 45909 1112
rect 45867 1063 45909 1072
rect 46059 1112 46101 1121
rect 46059 1072 46060 1112
rect 46100 1072 46101 1112
rect 46059 1063 46101 1072
rect 46251 1112 46293 1121
rect 46251 1072 46252 1112
rect 46292 1072 46293 1112
rect 46251 1063 46293 1072
rect 46443 1112 46485 1121
rect 46443 1072 46444 1112
rect 46484 1072 46485 1112
rect 46443 1063 46485 1072
rect 46635 1112 46677 1121
rect 46635 1072 46636 1112
rect 46676 1072 46677 1112
rect 46635 1063 46677 1072
rect 46827 1112 46869 1121
rect 46827 1072 46828 1112
rect 46868 1072 46869 1112
rect 46827 1063 46869 1072
rect 47019 1112 47061 1121
rect 47019 1072 47020 1112
rect 47060 1072 47061 1112
rect 47019 1063 47061 1072
rect 47211 1112 47253 1121
rect 47211 1072 47212 1112
rect 47252 1072 47253 1112
rect 47211 1063 47253 1072
rect 47403 1112 47445 1121
rect 47403 1072 47404 1112
rect 47444 1072 47445 1112
rect 47403 1063 47445 1072
rect 47595 1112 47637 1121
rect 47595 1072 47596 1112
rect 47636 1072 47637 1112
rect 47595 1063 47637 1072
rect 47787 1112 47829 1121
rect 47787 1072 47788 1112
rect 47828 1072 47829 1112
rect 47787 1063 47829 1072
rect 47979 1112 48021 1121
rect 47979 1072 47980 1112
rect 48020 1072 48021 1112
rect 47979 1063 48021 1072
rect 48171 1112 48213 1121
rect 48171 1072 48172 1112
rect 48212 1072 48213 1112
rect 48171 1063 48213 1072
rect 48363 1112 48405 1121
rect 48363 1072 48364 1112
rect 48404 1072 48405 1112
rect 48363 1063 48405 1072
rect 48555 1112 48597 1121
rect 48555 1072 48556 1112
rect 48596 1072 48597 1112
rect 48555 1063 48597 1072
rect 48747 1112 48789 1121
rect 48747 1072 48748 1112
rect 48788 1072 48789 1112
rect 48747 1063 48789 1072
rect 48939 1112 48981 1121
rect 48939 1072 48940 1112
rect 48980 1072 48981 1112
rect 48939 1063 48981 1072
rect 49131 1112 49173 1121
rect 49131 1072 49132 1112
rect 49172 1072 49173 1112
rect 49131 1063 49173 1072
rect 49323 1112 49365 1121
rect 49323 1072 49324 1112
rect 49364 1072 49365 1112
rect 49323 1063 49365 1072
rect 49515 1112 49557 1121
rect 49515 1072 49516 1112
rect 49556 1072 49557 1112
rect 49515 1063 49557 1072
rect 50379 1112 50421 1121
rect 50379 1072 50380 1112
rect 50420 1072 50421 1112
rect 50379 1063 50421 1072
rect 50571 1112 50613 1121
rect 50571 1072 50572 1112
rect 50612 1072 50613 1112
rect 50571 1063 50613 1072
rect 50955 1112 50997 1121
rect 50955 1072 50956 1112
rect 50996 1072 50997 1112
rect 50955 1063 50997 1072
rect 51435 1112 51477 1121
rect 51435 1072 51436 1112
rect 51476 1072 51477 1112
rect 51435 1063 51477 1072
rect 52203 1112 52245 1121
rect 52203 1072 52204 1112
rect 52244 1072 52245 1112
rect 52203 1063 52245 1072
rect 52491 1112 52533 1121
rect 52491 1072 52492 1112
rect 52532 1072 52533 1112
rect 52491 1063 52533 1072
rect 52683 1112 52725 1121
rect 52683 1072 52684 1112
rect 52724 1072 52725 1112
rect 52683 1063 52725 1072
rect 53547 1112 53589 1121
rect 53547 1072 53548 1112
rect 53588 1072 53589 1112
rect 53547 1063 53589 1072
rect 53739 1112 53781 1121
rect 53739 1072 53740 1112
rect 53780 1072 53781 1112
rect 53739 1063 53781 1072
rect 54123 1112 54165 1121
rect 54123 1072 54124 1112
rect 54164 1072 54165 1112
rect 54603 1084 54604 1124
rect 54644 1084 54645 1124
rect 54603 1075 54645 1084
rect 55083 1112 55125 1121
rect 54123 1063 54165 1072
rect 55083 1072 55084 1112
rect 55124 1072 55125 1112
rect 55083 1063 55125 1072
rect 55371 1112 55413 1121
rect 55371 1072 55372 1112
rect 55412 1072 55413 1112
rect 55371 1063 55413 1072
rect 55563 1112 55605 1121
rect 55563 1072 55564 1112
rect 55604 1072 55605 1112
rect 55563 1063 55605 1072
rect 56235 1112 56277 1121
rect 56235 1072 56236 1112
rect 56276 1072 56277 1112
rect 56235 1063 56277 1072
rect 56427 1112 56469 1121
rect 56427 1072 56428 1112
rect 56468 1072 56469 1112
rect 56427 1063 56469 1072
rect 56715 1115 56757 1124
rect 56715 1075 56716 1115
rect 56756 1075 56757 1115
rect 56715 1066 56757 1075
rect 57195 1112 57237 1121
rect 57195 1072 57196 1112
rect 57236 1072 57237 1112
rect 57195 1063 57237 1072
rect 57771 1112 57813 1121
rect 57771 1072 57772 1112
rect 57812 1072 57813 1112
rect 57771 1063 57813 1072
rect 58155 1112 58197 1121
rect 58155 1072 58156 1112
rect 58196 1072 58197 1112
rect 58155 1063 58197 1072
rect 58347 1112 58389 1121
rect 58347 1072 58348 1112
rect 58388 1072 58389 1112
rect 58347 1063 58389 1072
rect 59115 1112 59157 1121
rect 59115 1072 59116 1112
rect 59156 1072 59157 1112
rect 59115 1063 59157 1072
rect 59307 1112 59349 1121
rect 59307 1072 59308 1112
rect 59348 1072 59349 1112
rect 59307 1063 59349 1072
rect 59595 1112 59637 1121
rect 59595 1072 59596 1112
rect 59636 1072 59637 1112
rect 59595 1063 59637 1072
rect 60171 1112 60213 1121
rect 60171 1072 60172 1112
rect 60212 1072 60213 1112
rect 60171 1063 60213 1072
rect 60651 1112 60693 1121
rect 60651 1072 60652 1112
rect 60692 1072 60693 1112
rect 60651 1063 60693 1072
rect 60939 1112 60981 1121
rect 60939 1072 60940 1112
rect 60980 1072 60981 1112
rect 60939 1063 60981 1072
rect 61131 1112 61173 1121
rect 61131 1072 61132 1112
rect 61172 1072 61173 1112
rect 61131 1063 61173 1072
rect 62667 1112 62709 1121
rect 62667 1072 62668 1112
rect 62708 1072 62709 1112
rect 63051 1112 63093 1121
rect 62667 1063 62709 1072
rect 62859 1101 62901 1110
rect 41934 1060 41992 1061
rect 62859 1061 62860 1101
rect 62900 1061 62901 1101
rect 63051 1072 63052 1112
rect 63092 1072 63093 1112
rect 63051 1063 63093 1072
rect 63243 1112 63285 1121
rect 63243 1072 63244 1112
rect 63284 1072 63285 1112
rect 63243 1063 63285 1072
rect 63435 1112 63477 1121
rect 63435 1072 63436 1112
rect 63476 1072 63477 1112
rect 63435 1063 63477 1072
rect 63627 1112 63669 1121
rect 63627 1072 63628 1112
rect 63668 1072 63669 1112
rect 63819 1085 63820 1125
rect 63860 1085 63861 1125
rect 66884 1125 66926 1134
rect 63819 1076 63861 1085
rect 64011 1112 64053 1121
rect 63627 1063 63669 1072
rect 64011 1072 64012 1112
rect 64052 1072 64053 1112
rect 64011 1063 64053 1072
rect 64203 1112 64245 1121
rect 64203 1072 64204 1112
rect 64244 1072 64245 1112
rect 64203 1063 64245 1072
rect 64395 1112 64437 1121
rect 64395 1072 64396 1112
rect 64436 1072 64437 1112
rect 64395 1063 64437 1072
rect 64587 1112 64629 1121
rect 64587 1072 64588 1112
rect 64628 1072 64629 1112
rect 64587 1063 64629 1072
rect 64779 1112 64821 1121
rect 64779 1072 64780 1112
rect 64820 1072 64821 1112
rect 64779 1063 64821 1072
rect 64971 1112 65013 1121
rect 64971 1072 64972 1112
rect 65012 1072 65013 1112
rect 64971 1063 65013 1072
rect 65163 1112 65205 1121
rect 65163 1072 65164 1112
rect 65204 1072 65205 1112
rect 65163 1063 65205 1072
rect 65355 1112 65397 1121
rect 65355 1072 65356 1112
rect 65396 1072 65397 1112
rect 65355 1063 65397 1072
rect 65547 1112 65589 1121
rect 65547 1072 65548 1112
rect 65588 1072 65589 1112
rect 65547 1063 65589 1072
rect 65739 1112 65781 1121
rect 65739 1072 65740 1112
rect 65780 1072 65781 1112
rect 65739 1063 65781 1072
rect 65931 1112 65973 1121
rect 65931 1072 65932 1112
rect 65972 1072 65973 1112
rect 65931 1063 65973 1072
rect 66123 1112 66165 1121
rect 66123 1072 66124 1112
rect 66164 1072 66165 1112
rect 66123 1063 66165 1072
rect 66315 1112 66357 1121
rect 66315 1072 66316 1112
rect 66356 1072 66357 1112
rect 66315 1063 66357 1072
rect 66507 1112 66549 1121
rect 66507 1072 66508 1112
rect 66548 1072 66549 1112
rect 66507 1063 66549 1072
rect 66699 1112 66741 1121
rect 66699 1072 66700 1112
rect 66740 1072 66741 1112
rect 66884 1085 66885 1125
rect 66925 1085 66926 1125
rect 66884 1076 66926 1085
rect 67083 1112 67125 1121
rect 66699 1063 66741 1072
rect 67083 1072 67084 1112
rect 67124 1072 67125 1112
rect 67083 1063 67125 1072
rect 67275 1112 67317 1121
rect 67275 1072 67276 1112
rect 67316 1072 67317 1112
rect 67275 1063 67317 1072
rect 67467 1112 67509 1121
rect 67467 1072 67468 1112
rect 67508 1072 67509 1112
rect 67467 1063 67509 1072
rect 67659 1112 67701 1121
rect 67659 1072 67660 1112
rect 67700 1072 67701 1112
rect 67659 1063 67701 1072
rect 67851 1112 67893 1121
rect 67851 1072 67852 1112
rect 67892 1072 67893 1112
rect 67851 1063 67893 1072
rect 68043 1112 68085 1121
rect 68043 1072 68044 1112
rect 68084 1072 68085 1112
rect 68043 1063 68085 1072
rect 68235 1112 68277 1121
rect 68235 1072 68236 1112
rect 68276 1072 68277 1112
rect 68235 1063 68277 1072
rect 68427 1112 68469 1121
rect 68427 1072 68428 1112
rect 68468 1072 68469 1112
rect 68427 1063 68469 1072
rect 68619 1112 68661 1121
rect 68619 1072 68620 1112
rect 68660 1072 68661 1112
rect 68619 1063 68661 1072
rect 68811 1112 68853 1121
rect 68811 1072 68812 1112
rect 68852 1072 68853 1112
rect 68811 1063 68853 1072
rect 69003 1112 69045 1121
rect 69003 1072 69004 1112
rect 69044 1072 69045 1112
rect 69003 1063 69045 1072
rect 69195 1112 69237 1121
rect 69195 1072 69196 1112
rect 69236 1072 69237 1112
rect 69195 1063 69237 1072
rect 69387 1112 69429 1121
rect 69387 1072 69388 1112
rect 69428 1072 69429 1112
rect 69771 1112 69813 1121
rect 69387 1063 69429 1072
rect 69581 1109 69639 1110
rect 69581 1069 69590 1109
rect 69630 1069 69639 1109
rect 69581 1068 69639 1069
rect 69771 1072 69772 1112
rect 69812 1072 69813 1112
rect 69771 1063 69813 1072
rect 69963 1112 70005 1121
rect 69963 1072 69964 1112
rect 70004 1072 70005 1112
rect 69963 1063 70005 1072
rect 70155 1112 70197 1121
rect 70155 1072 70156 1112
rect 70196 1072 70197 1112
rect 70155 1063 70197 1072
rect 70347 1112 70389 1121
rect 70347 1072 70348 1112
rect 70388 1072 70389 1112
rect 70347 1063 70389 1072
rect 70520 1117 70562 1126
rect 85899 1125 85941 1134
rect 70520 1077 70521 1117
rect 70561 1077 70562 1117
rect 70520 1068 70562 1077
rect 70731 1112 70773 1121
rect 70731 1072 70732 1112
rect 70772 1072 70773 1112
rect 70731 1063 70773 1072
rect 70923 1112 70965 1121
rect 70923 1072 70924 1112
rect 70964 1072 70965 1112
rect 70923 1063 70965 1072
rect 71115 1112 71157 1121
rect 71115 1072 71116 1112
rect 71156 1072 71157 1112
rect 71115 1063 71157 1072
rect 71307 1112 71349 1121
rect 71307 1072 71308 1112
rect 71348 1072 71349 1112
rect 71307 1063 71349 1072
rect 71499 1112 71541 1121
rect 71499 1072 71500 1112
rect 71540 1072 71541 1112
rect 71499 1063 71541 1072
rect 71691 1112 71733 1121
rect 71691 1072 71692 1112
rect 71732 1072 71733 1112
rect 71691 1063 71733 1072
rect 71883 1112 71925 1121
rect 71883 1072 71884 1112
rect 71924 1072 71925 1112
rect 71883 1063 71925 1072
rect 72075 1112 72117 1121
rect 72075 1072 72076 1112
rect 72116 1072 72117 1112
rect 72075 1063 72117 1072
rect 72267 1112 72309 1121
rect 72267 1072 72268 1112
rect 72308 1072 72309 1112
rect 72267 1063 72309 1072
rect 72459 1112 72501 1121
rect 72459 1072 72460 1112
rect 72500 1072 72501 1112
rect 72459 1063 72501 1072
rect 72651 1112 72693 1121
rect 72651 1072 72652 1112
rect 72692 1072 72693 1112
rect 72651 1063 72693 1072
rect 72843 1112 72885 1121
rect 72843 1072 72844 1112
rect 72884 1072 72885 1112
rect 72843 1063 72885 1072
rect 73035 1112 73077 1121
rect 73035 1072 73036 1112
rect 73076 1072 73077 1112
rect 73035 1063 73077 1072
rect 73227 1112 73269 1121
rect 73227 1072 73228 1112
rect 73268 1072 73269 1112
rect 73227 1063 73269 1072
rect 73419 1112 73461 1121
rect 73419 1072 73420 1112
rect 73460 1072 73461 1112
rect 73419 1063 73461 1072
rect 73611 1112 73653 1121
rect 73611 1072 73612 1112
rect 73652 1072 73653 1112
rect 73611 1063 73653 1072
rect 73803 1112 73845 1121
rect 73803 1072 73804 1112
rect 73844 1072 73845 1112
rect 73803 1063 73845 1072
rect 73995 1112 74037 1121
rect 73995 1072 73996 1112
rect 74036 1072 74037 1112
rect 73995 1063 74037 1072
rect 74187 1112 74229 1121
rect 74187 1072 74188 1112
rect 74228 1072 74229 1112
rect 74187 1063 74229 1072
rect 74379 1112 74421 1121
rect 74379 1072 74380 1112
rect 74420 1072 74421 1112
rect 74379 1063 74421 1072
rect 74571 1112 74613 1121
rect 74571 1072 74572 1112
rect 74612 1072 74613 1112
rect 74571 1063 74613 1072
rect 74763 1112 74805 1121
rect 74763 1072 74764 1112
rect 74804 1072 74805 1112
rect 74763 1063 74805 1072
rect 74955 1112 74997 1121
rect 74955 1072 74956 1112
rect 74996 1072 74997 1112
rect 74955 1063 74997 1072
rect 75147 1112 75189 1121
rect 75147 1072 75148 1112
rect 75188 1072 75189 1112
rect 75147 1063 75189 1072
rect 75339 1113 75381 1122
rect 75339 1073 75340 1113
rect 75380 1073 75381 1113
rect 75339 1064 75381 1073
rect 75531 1112 75573 1121
rect 75531 1072 75532 1112
rect 75572 1072 75573 1112
rect 75531 1063 75573 1072
rect 75723 1112 75765 1121
rect 75723 1072 75724 1112
rect 75764 1072 75765 1112
rect 75723 1063 75765 1072
rect 75915 1112 75957 1121
rect 75915 1072 75916 1112
rect 75956 1072 75957 1112
rect 75915 1063 75957 1072
rect 76107 1112 76149 1121
rect 76107 1072 76108 1112
rect 76148 1072 76149 1112
rect 76107 1063 76149 1072
rect 76299 1112 76341 1121
rect 76299 1072 76300 1112
rect 76340 1072 76341 1112
rect 76683 1112 76725 1121
rect 76299 1063 76341 1072
rect 76491 1101 76533 1110
rect 62859 1052 62901 1061
rect 76491 1061 76492 1101
rect 76532 1061 76533 1101
rect 76683 1072 76684 1112
rect 76724 1072 76725 1112
rect 76683 1063 76725 1072
rect 76875 1112 76917 1121
rect 76875 1072 76876 1112
rect 76916 1072 76917 1112
rect 76875 1063 76917 1072
rect 77067 1112 77109 1121
rect 77067 1072 77068 1112
rect 77108 1072 77109 1112
rect 77067 1063 77109 1072
rect 77259 1112 77301 1121
rect 77259 1072 77260 1112
rect 77300 1072 77301 1112
rect 77259 1063 77301 1072
rect 77451 1112 77493 1121
rect 77451 1072 77452 1112
rect 77492 1072 77493 1112
rect 77451 1063 77493 1072
rect 77643 1112 77685 1121
rect 77643 1072 77644 1112
rect 77684 1072 77685 1112
rect 77643 1063 77685 1072
rect 77835 1112 77877 1121
rect 77835 1072 77836 1112
rect 77876 1072 77877 1112
rect 77835 1063 77877 1072
rect 78027 1112 78069 1121
rect 78027 1072 78028 1112
rect 78068 1072 78069 1112
rect 78027 1063 78069 1072
rect 78219 1112 78261 1121
rect 78219 1072 78220 1112
rect 78260 1072 78261 1112
rect 78219 1063 78261 1072
rect 78411 1112 78453 1121
rect 78411 1072 78412 1112
rect 78452 1072 78453 1112
rect 78411 1063 78453 1072
rect 78603 1112 78645 1121
rect 78603 1072 78604 1112
rect 78644 1072 78645 1112
rect 78603 1063 78645 1072
rect 78795 1112 78837 1121
rect 78795 1072 78796 1112
rect 78836 1072 78837 1112
rect 78795 1063 78837 1072
rect 78987 1112 79029 1121
rect 78987 1072 78988 1112
rect 79028 1072 79029 1112
rect 78987 1063 79029 1072
rect 79179 1112 79221 1121
rect 79179 1072 79180 1112
rect 79220 1072 79221 1112
rect 79179 1063 79221 1072
rect 79371 1112 79413 1121
rect 79371 1072 79372 1112
rect 79412 1072 79413 1112
rect 79371 1063 79413 1072
rect 79563 1112 79605 1121
rect 79563 1072 79564 1112
rect 79604 1072 79605 1112
rect 79563 1063 79605 1072
rect 79755 1112 79797 1121
rect 79755 1072 79756 1112
rect 79796 1072 79797 1112
rect 79755 1063 79797 1072
rect 79947 1112 79989 1121
rect 79947 1072 79948 1112
rect 79988 1072 79989 1112
rect 79947 1063 79989 1072
rect 80139 1112 80181 1121
rect 80139 1072 80140 1112
rect 80180 1072 80181 1112
rect 80139 1063 80181 1072
rect 80331 1112 80373 1121
rect 80331 1072 80332 1112
rect 80372 1072 80373 1112
rect 80331 1063 80373 1072
rect 80523 1112 80565 1121
rect 80523 1072 80524 1112
rect 80564 1072 80565 1112
rect 80523 1063 80565 1072
rect 80907 1112 80949 1121
rect 80907 1072 80908 1112
rect 80948 1072 80949 1112
rect 80907 1063 80949 1072
rect 81099 1112 81141 1121
rect 81099 1072 81100 1112
rect 81140 1072 81141 1112
rect 81099 1063 81141 1072
rect 81291 1112 81333 1121
rect 81291 1072 81292 1112
rect 81332 1072 81333 1112
rect 81291 1063 81333 1072
rect 81483 1112 81525 1121
rect 81483 1072 81484 1112
rect 81524 1072 81525 1112
rect 81483 1063 81525 1072
rect 81675 1112 81717 1121
rect 81675 1072 81676 1112
rect 81716 1072 81717 1112
rect 81675 1063 81717 1072
rect 81867 1112 81909 1121
rect 81867 1072 81868 1112
rect 81908 1072 81909 1112
rect 81867 1063 81909 1072
rect 82059 1112 82101 1121
rect 82059 1072 82060 1112
rect 82100 1072 82101 1112
rect 82059 1063 82101 1072
rect 82251 1112 82293 1121
rect 82251 1072 82252 1112
rect 82292 1072 82293 1112
rect 82251 1063 82293 1072
rect 82443 1112 82485 1121
rect 82443 1072 82444 1112
rect 82484 1072 82485 1112
rect 82443 1063 82485 1072
rect 82635 1112 82677 1121
rect 82635 1072 82636 1112
rect 82676 1072 82677 1112
rect 82635 1063 82677 1072
rect 82827 1112 82869 1121
rect 82827 1072 82828 1112
rect 82868 1072 82869 1112
rect 82827 1063 82869 1072
rect 83019 1112 83061 1121
rect 83019 1072 83020 1112
rect 83060 1072 83061 1112
rect 83019 1063 83061 1072
rect 83211 1112 83253 1121
rect 83211 1072 83212 1112
rect 83252 1072 83253 1112
rect 83595 1112 83637 1121
rect 83211 1063 83253 1072
rect 83384 1109 83442 1110
rect 83384 1069 83393 1109
rect 83433 1069 83442 1109
rect 83384 1068 83442 1069
rect 83595 1072 83596 1112
rect 83636 1072 83637 1112
rect 83595 1063 83637 1072
rect 83792 1109 83834 1118
rect 83792 1069 83793 1109
rect 83833 1069 83834 1109
rect 76491 1052 76533 1061
rect 83792 1060 83834 1069
rect 83979 1112 84021 1121
rect 83979 1072 83980 1112
rect 84020 1072 84021 1112
rect 83979 1063 84021 1072
rect 84171 1112 84213 1121
rect 84171 1072 84172 1112
rect 84212 1072 84213 1112
rect 84171 1063 84213 1072
rect 84363 1112 84405 1121
rect 84363 1072 84364 1112
rect 84404 1072 84405 1112
rect 84363 1063 84405 1072
rect 84555 1112 84597 1121
rect 84555 1072 84556 1112
rect 84596 1072 84597 1112
rect 84555 1063 84597 1072
rect 84747 1112 84789 1121
rect 84747 1072 84748 1112
rect 84788 1072 84789 1112
rect 84747 1063 84789 1072
rect 84939 1112 84981 1121
rect 84939 1072 84940 1112
rect 84980 1072 84981 1112
rect 84939 1063 84981 1072
rect 85131 1112 85173 1121
rect 85131 1072 85132 1112
rect 85172 1072 85173 1112
rect 85131 1063 85173 1072
rect 85323 1112 85365 1121
rect 85323 1072 85324 1112
rect 85364 1072 85365 1112
rect 85323 1063 85365 1072
rect 85515 1112 85557 1121
rect 85515 1072 85516 1112
rect 85556 1072 85557 1112
rect 85515 1063 85557 1072
rect 85707 1112 85749 1121
rect 85707 1072 85708 1112
rect 85748 1072 85749 1112
rect 85899 1085 85900 1125
rect 85940 1085 85941 1125
rect 88395 1125 88437 1134
rect 85899 1076 85941 1085
rect 86091 1112 86133 1121
rect 85707 1063 85749 1072
rect 86091 1072 86092 1112
rect 86132 1072 86133 1112
rect 86091 1063 86133 1072
rect 86283 1112 86325 1121
rect 86283 1072 86284 1112
rect 86324 1072 86325 1112
rect 86283 1063 86325 1072
rect 86475 1112 86517 1121
rect 86475 1072 86476 1112
rect 86516 1072 86517 1112
rect 86475 1063 86517 1072
rect 86667 1112 86709 1121
rect 86667 1072 86668 1112
rect 86708 1072 86709 1112
rect 86667 1063 86709 1072
rect 86859 1112 86901 1121
rect 86859 1072 86860 1112
rect 86900 1072 86901 1112
rect 86859 1063 86901 1072
rect 87051 1112 87093 1121
rect 87051 1072 87052 1112
rect 87092 1072 87093 1112
rect 87051 1063 87093 1072
rect 87243 1112 87285 1121
rect 87243 1072 87244 1112
rect 87284 1072 87285 1112
rect 87243 1063 87285 1072
rect 87435 1112 87477 1121
rect 87435 1072 87436 1112
rect 87476 1072 87477 1112
rect 87435 1063 87477 1072
rect 87627 1112 87669 1121
rect 87627 1072 87628 1112
rect 87668 1072 87669 1112
rect 87627 1063 87669 1072
rect 87819 1112 87861 1121
rect 87819 1072 87820 1112
rect 87860 1072 87861 1112
rect 87819 1063 87861 1072
rect 88011 1112 88053 1121
rect 88011 1072 88012 1112
rect 88052 1072 88053 1112
rect 88011 1063 88053 1072
rect 88203 1112 88245 1121
rect 88203 1072 88204 1112
rect 88244 1072 88245 1112
rect 88395 1085 88396 1125
rect 88436 1085 88437 1125
rect 97218 1125 97276 1126
rect 88395 1076 88437 1085
rect 88587 1112 88629 1121
rect 88203 1063 88245 1072
rect 88587 1072 88588 1112
rect 88628 1072 88629 1112
rect 88587 1063 88629 1072
rect 88779 1112 88821 1121
rect 88779 1072 88780 1112
rect 88820 1072 88821 1112
rect 88779 1063 88821 1072
rect 88971 1112 89013 1121
rect 88971 1072 88972 1112
rect 89012 1072 89013 1112
rect 88971 1063 89013 1072
rect 89163 1112 89205 1121
rect 89163 1072 89164 1112
rect 89204 1072 89205 1112
rect 89163 1063 89205 1072
rect 89355 1112 89397 1121
rect 89355 1072 89356 1112
rect 89396 1072 89397 1112
rect 89355 1063 89397 1072
rect 89547 1112 89589 1121
rect 89547 1072 89548 1112
rect 89588 1072 89589 1112
rect 89547 1063 89589 1072
rect 89739 1112 89781 1121
rect 89739 1072 89740 1112
rect 89780 1072 89781 1112
rect 89739 1063 89781 1072
rect 89931 1112 89973 1121
rect 89931 1072 89932 1112
rect 89972 1072 89973 1112
rect 89931 1063 89973 1072
rect 90123 1112 90165 1121
rect 90123 1072 90124 1112
rect 90164 1072 90165 1112
rect 90123 1063 90165 1072
rect 90315 1112 90357 1121
rect 90315 1072 90316 1112
rect 90356 1072 90357 1112
rect 90315 1063 90357 1072
rect 90507 1112 90549 1121
rect 90507 1072 90508 1112
rect 90548 1072 90549 1112
rect 90891 1112 90933 1121
rect 90507 1063 90549 1072
rect 90699 1101 90741 1110
rect 90699 1061 90700 1101
rect 90740 1061 90741 1101
rect 90891 1072 90892 1112
rect 90932 1072 90933 1112
rect 90891 1063 90933 1072
rect 91083 1112 91125 1121
rect 91083 1072 91084 1112
rect 91124 1072 91125 1112
rect 91083 1063 91125 1072
rect 91275 1112 91317 1121
rect 91275 1072 91276 1112
rect 91316 1072 91317 1112
rect 91275 1063 91317 1072
rect 91467 1112 91509 1121
rect 91467 1072 91468 1112
rect 91508 1072 91509 1112
rect 91467 1063 91509 1072
rect 91659 1112 91701 1121
rect 91659 1072 91660 1112
rect 91700 1072 91701 1112
rect 91659 1063 91701 1072
rect 91851 1112 91893 1121
rect 91851 1072 91852 1112
rect 91892 1072 91893 1112
rect 91851 1063 91893 1072
rect 92043 1112 92085 1121
rect 92043 1072 92044 1112
rect 92084 1072 92085 1112
rect 92043 1063 92085 1072
rect 92235 1112 92277 1121
rect 92235 1072 92236 1112
rect 92276 1072 92277 1112
rect 92235 1063 92277 1072
rect 92427 1112 92469 1121
rect 92427 1072 92428 1112
rect 92468 1072 92469 1112
rect 92427 1063 92469 1072
rect 92619 1112 92661 1121
rect 92619 1072 92620 1112
rect 92660 1072 92661 1112
rect 92619 1063 92661 1072
rect 92811 1112 92853 1121
rect 92811 1072 92812 1112
rect 92852 1072 92853 1112
rect 92811 1063 92853 1072
rect 93003 1112 93045 1121
rect 93003 1072 93004 1112
rect 93044 1072 93045 1112
rect 93003 1063 93045 1072
rect 93195 1112 93237 1121
rect 93195 1072 93196 1112
rect 93236 1072 93237 1112
rect 93195 1063 93237 1072
rect 93387 1112 93429 1121
rect 93387 1072 93388 1112
rect 93428 1072 93429 1112
rect 93387 1063 93429 1072
rect 93579 1112 93621 1121
rect 93579 1072 93580 1112
rect 93620 1072 93621 1112
rect 93579 1063 93621 1072
rect 93771 1112 93813 1121
rect 93771 1072 93772 1112
rect 93812 1072 93813 1112
rect 93771 1063 93813 1072
rect 93963 1112 94005 1121
rect 93963 1072 93964 1112
rect 94004 1072 94005 1112
rect 93963 1063 94005 1072
rect 94155 1112 94197 1121
rect 94155 1072 94156 1112
rect 94196 1072 94197 1112
rect 94155 1063 94197 1072
rect 94347 1112 94389 1121
rect 94347 1072 94348 1112
rect 94388 1072 94389 1112
rect 94347 1063 94389 1072
rect 94539 1101 94581 1110
rect 90699 1052 90741 1061
rect 94539 1061 94540 1101
rect 94580 1061 94581 1101
rect 94539 1052 94581 1061
rect 94731 1109 94773 1118
rect 95499 1112 95541 1121
rect 94731 1069 94732 1109
rect 94772 1069 94773 1109
rect 94731 1060 94773 1069
rect 94923 1101 94965 1110
rect 94923 1061 94924 1101
rect 94964 1061 94965 1101
rect 94923 1052 94965 1061
rect 95115 1101 95157 1110
rect 95115 1061 95116 1101
rect 95156 1061 95157 1101
rect 95115 1052 95157 1061
rect 95307 1101 95349 1110
rect 95307 1061 95308 1101
rect 95348 1061 95349 1101
rect 95499 1072 95500 1112
rect 95540 1072 95541 1112
rect 95499 1063 95541 1072
rect 95698 1109 95740 1118
rect 95698 1069 95699 1109
rect 95739 1069 95740 1109
rect 95307 1052 95349 1061
rect 95698 1060 95740 1069
rect 95883 1112 95925 1121
rect 95883 1072 95884 1112
rect 95924 1072 95925 1112
rect 95883 1063 95925 1072
rect 96075 1112 96117 1121
rect 96075 1072 96076 1112
rect 96116 1072 96117 1112
rect 96075 1063 96117 1072
rect 96267 1112 96309 1121
rect 96267 1072 96268 1112
rect 96308 1072 96309 1112
rect 96267 1063 96309 1072
rect 96459 1112 96501 1121
rect 96459 1072 96460 1112
rect 96500 1072 96501 1112
rect 96459 1063 96501 1072
rect 96651 1112 96693 1121
rect 96651 1072 96652 1112
rect 96692 1072 96693 1112
rect 96651 1063 96693 1072
rect 96843 1112 96885 1121
rect 96843 1072 96844 1112
rect 96884 1072 96885 1112
rect 96843 1063 96885 1072
rect 97035 1112 97077 1121
rect 97035 1072 97036 1112
rect 97076 1072 97077 1112
rect 97218 1085 97227 1125
rect 97267 1085 97276 1125
rect 97986 1125 98044 1126
rect 97218 1084 97276 1085
rect 97419 1112 97461 1121
rect 97035 1063 97077 1072
rect 97419 1072 97420 1112
rect 97460 1072 97461 1112
rect 97419 1063 97461 1072
rect 97611 1112 97653 1121
rect 97611 1072 97612 1112
rect 97652 1072 97653 1112
rect 97611 1063 97653 1072
rect 97803 1112 97845 1121
rect 97803 1072 97804 1112
rect 97844 1072 97845 1112
rect 97986 1085 97995 1125
rect 98035 1085 98044 1125
rect 97986 1084 98044 1085
rect 98187 1112 98229 1121
rect 97803 1063 97845 1072
rect 98187 1072 98188 1112
rect 98228 1072 98229 1112
rect 98187 1063 98229 1072
rect 98379 1112 98421 1121
rect 98379 1072 98380 1112
rect 98420 1072 98421 1112
rect 98379 1063 98421 1072
rect 98571 1112 98613 1121
rect 98571 1072 98572 1112
rect 98612 1072 98613 1112
rect 98571 1063 98613 1072
rect 98763 1112 98805 1121
rect 98763 1072 98764 1112
rect 98804 1072 98805 1112
rect 98763 1063 98805 1072
rect 98955 1112 98997 1121
rect 98955 1072 98956 1112
rect 98996 1072 98997 1112
rect 98955 1063 98997 1072
rect 99147 1112 99189 1121
rect 99147 1072 99148 1112
rect 99188 1072 99189 1112
rect 99147 1063 99189 1072
rect 5355 1028 5397 1037
rect 5355 988 5356 1028
rect 5396 988 5397 1028
rect 5355 979 5397 988
rect 35019 1028 35061 1037
rect 35019 988 35020 1028
rect 35060 988 35061 1028
rect 35019 979 35061 988
rect 67755 1028 67797 1037
rect 67755 988 67756 1028
rect 67796 988 67797 1028
rect 67755 979 67797 988
rect 89067 1028 89109 1037
rect 89067 988 89068 1028
rect 89108 988 89109 1028
rect 89067 979 89109 988
rect 91371 1028 91413 1037
rect 91371 988 91372 1028
rect 91412 988 91413 1028
rect 91371 979 91413 988
rect 92139 1028 92181 1037
rect 92139 988 92140 1028
rect 92180 988 92181 1028
rect 92139 979 92181 988
rect 97899 1028 97941 1037
rect 97899 988 97900 1028
rect 97940 988 97941 1028
rect 97899 979 97941 988
rect 1131 944 1173 953
rect 1131 904 1132 944
rect 1172 904 1173 944
rect 1131 895 1173 904
rect 1515 944 1557 953
rect 1515 904 1516 944
rect 1556 904 1557 944
rect 1515 895 1557 904
rect 1899 944 1941 953
rect 1899 904 1900 944
rect 1940 904 1941 944
rect 1899 895 1941 904
rect 2283 944 2325 953
rect 2283 904 2284 944
rect 2324 904 2325 944
rect 2283 895 2325 904
rect 2667 944 2709 953
rect 2667 904 2668 944
rect 2708 904 2709 944
rect 2667 895 2709 904
rect 3051 944 3093 953
rect 3051 904 3052 944
rect 3092 904 3093 944
rect 3051 895 3093 904
rect 3435 944 3477 953
rect 3435 904 3436 944
rect 3476 904 3477 944
rect 3435 895 3477 904
rect 3819 944 3861 953
rect 3819 904 3820 944
rect 3860 904 3861 944
rect 3819 895 3861 904
rect 4203 944 4245 953
rect 4203 904 4204 944
rect 4244 904 4245 944
rect 4203 895 4245 904
rect 4587 944 4629 953
rect 4587 904 4588 944
rect 4628 904 4629 944
rect 4587 895 4629 904
rect 4971 944 5013 953
rect 4971 904 4972 944
rect 5012 904 5013 944
rect 4971 895 5013 904
rect 5739 944 5781 953
rect 5739 904 5740 944
rect 5780 904 5781 944
rect 5739 895 5781 904
rect 6123 944 6165 953
rect 6123 904 6124 944
rect 6164 904 6165 944
rect 6123 895 6165 904
rect 6507 944 6549 953
rect 6507 904 6508 944
rect 6548 904 6549 944
rect 6507 895 6549 904
rect 7275 944 7317 953
rect 7275 904 7276 944
rect 7316 904 7317 944
rect 7275 895 7317 904
rect 7659 944 7701 953
rect 7659 904 7660 944
rect 7700 904 7701 944
rect 7659 895 7701 904
rect 8043 944 8085 953
rect 8043 904 8044 944
rect 8084 904 8085 944
rect 8043 895 8085 904
rect 8427 944 8469 953
rect 8427 904 8428 944
rect 8468 904 8469 944
rect 8427 895 8469 904
rect 8811 944 8853 953
rect 8811 904 8812 944
rect 8852 904 8853 944
rect 8811 895 8853 904
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 9579 944 9621 953
rect 9579 904 9580 944
rect 9620 904 9621 944
rect 9579 895 9621 904
rect 9963 944 10005 953
rect 9963 904 9964 944
rect 10004 904 10005 944
rect 9963 895 10005 904
rect 10347 944 10389 953
rect 10347 904 10348 944
rect 10388 904 10389 944
rect 10347 895 10389 904
rect 10731 944 10773 953
rect 10731 904 10732 944
rect 10772 904 10773 944
rect 10731 895 10773 904
rect 11115 944 11157 953
rect 11115 904 11116 944
rect 11156 904 11157 944
rect 11115 895 11157 904
rect 11499 944 11541 953
rect 11499 904 11500 944
rect 11540 904 11541 944
rect 11499 895 11541 904
rect 11883 944 11925 953
rect 11883 904 11884 944
rect 11924 904 11925 944
rect 11883 895 11925 904
rect 12267 944 12309 953
rect 12267 904 12268 944
rect 12308 904 12309 944
rect 12267 895 12309 904
rect 12651 944 12693 953
rect 12651 904 12652 944
rect 12692 904 12693 944
rect 12651 895 12693 904
rect 13035 944 13077 953
rect 13035 904 13036 944
rect 13076 904 13077 944
rect 13035 895 13077 904
rect 13419 944 13461 953
rect 13419 904 13420 944
rect 13460 904 13461 944
rect 13419 895 13461 904
rect 13803 944 13845 953
rect 13803 904 13804 944
rect 13844 904 13845 944
rect 13803 895 13845 904
rect 14571 944 14613 953
rect 14571 904 14572 944
rect 14612 904 14613 944
rect 14571 895 14613 904
rect 14955 944 14997 953
rect 14955 904 14956 944
rect 14996 904 14997 944
rect 14955 895 14997 904
rect 15339 944 15381 953
rect 15339 904 15340 944
rect 15380 904 15381 944
rect 15339 895 15381 904
rect 15723 944 15765 953
rect 15723 904 15724 944
rect 15764 904 15765 944
rect 15723 895 15765 904
rect 16107 944 16149 953
rect 16107 904 16108 944
rect 16148 904 16149 944
rect 16107 895 16149 904
rect 16875 944 16917 953
rect 16875 904 16876 944
rect 16916 904 16917 944
rect 16875 895 16917 904
rect 17259 944 17301 953
rect 17259 904 17260 944
rect 17300 904 17301 944
rect 17259 895 17301 904
rect 17643 944 17685 953
rect 17643 904 17644 944
rect 17684 904 17685 944
rect 17643 895 17685 904
rect 18027 944 18069 953
rect 18027 904 18028 944
rect 18068 904 18069 944
rect 18027 895 18069 904
rect 18411 944 18453 953
rect 18411 904 18412 944
rect 18452 904 18453 944
rect 18411 895 18453 904
rect 18795 944 18837 953
rect 18795 904 18796 944
rect 18836 904 18837 944
rect 18795 895 18837 904
rect 19179 944 19221 953
rect 19179 904 19180 944
rect 19220 904 19221 944
rect 19179 895 19221 904
rect 19563 944 19605 953
rect 19563 904 19564 944
rect 19604 904 19605 944
rect 19563 895 19605 904
rect 19947 944 19989 953
rect 19947 904 19948 944
rect 19988 904 19989 944
rect 19947 895 19989 904
rect 20715 944 20757 953
rect 20715 904 20716 944
rect 20756 904 20757 944
rect 20715 895 20757 904
rect 21099 944 21141 953
rect 21099 904 21100 944
rect 21140 904 21141 944
rect 21099 895 21141 904
rect 21483 944 21525 953
rect 21483 904 21484 944
rect 21524 904 21525 944
rect 21483 895 21525 904
rect 21867 944 21909 953
rect 21867 904 21868 944
rect 21908 904 21909 944
rect 21867 895 21909 904
rect 22251 944 22293 953
rect 22251 904 22252 944
rect 22292 904 22293 944
rect 22251 895 22293 904
rect 22635 944 22677 953
rect 22635 904 22636 944
rect 22676 904 22677 944
rect 22635 895 22677 904
rect 23019 944 23061 953
rect 23019 904 23020 944
rect 23060 904 23061 944
rect 23019 895 23061 904
rect 23403 944 23445 953
rect 23403 904 23404 944
rect 23444 904 23445 944
rect 23403 895 23445 904
rect 23787 944 23829 953
rect 23787 904 23788 944
rect 23828 904 23829 944
rect 23787 895 23829 904
rect 24171 944 24213 953
rect 24171 904 24172 944
rect 24212 904 24213 944
rect 24171 895 24213 904
rect 24939 944 24981 953
rect 24939 904 24940 944
rect 24980 904 24981 944
rect 24939 895 24981 904
rect 25611 944 25653 953
rect 25611 904 25612 944
rect 25652 904 25653 944
rect 25611 895 25653 904
rect 25995 944 26037 953
rect 25995 904 25996 944
rect 26036 904 26037 944
rect 25995 895 26037 904
rect 26379 944 26421 953
rect 26379 904 26380 944
rect 26420 904 26421 944
rect 26379 895 26421 904
rect 26763 944 26805 953
rect 26763 904 26764 944
rect 26804 904 26805 944
rect 26763 895 26805 904
rect 27147 944 27189 953
rect 27147 904 27148 944
rect 27188 904 27189 944
rect 27147 895 27189 904
rect 27531 944 27573 953
rect 27531 904 27532 944
rect 27572 904 27573 944
rect 27531 895 27573 904
rect 27915 944 27957 953
rect 27915 904 27916 944
rect 27956 904 27957 944
rect 27915 895 27957 904
rect 28299 944 28341 953
rect 28299 904 28300 944
rect 28340 904 28341 944
rect 28299 895 28341 904
rect 28683 944 28725 953
rect 28683 904 28684 944
rect 28724 904 28725 944
rect 28683 895 28725 904
rect 29067 944 29109 953
rect 29067 904 29068 944
rect 29108 904 29109 944
rect 29067 895 29109 904
rect 29451 944 29493 953
rect 29451 904 29452 944
rect 29492 904 29493 944
rect 29451 895 29493 904
rect 29835 944 29877 953
rect 29835 904 29836 944
rect 29876 904 29877 944
rect 29835 895 29877 904
rect 30219 944 30261 953
rect 30219 904 30220 944
rect 30260 904 30261 944
rect 30219 895 30261 904
rect 30987 944 31029 953
rect 30987 904 30988 944
rect 31028 904 31029 944
rect 30987 895 31029 904
rect 31947 944 31989 953
rect 31947 904 31948 944
rect 31988 904 31989 944
rect 31947 895 31989 904
rect 32331 944 32373 953
rect 32331 904 32332 944
rect 32372 904 32373 944
rect 32331 895 32373 904
rect 32715 944 32757 953
rect 32715 904 32716 944
rect 32756 904 32757 944
rect 32715 895 32757 904
rect 33099 944 33141 953
rect 33099 904 33100 944
rect 33140 904 33141 944
rect 33099 895 33141 904
rect 33483 944 33525 953
rect 33483 904 33484 944
rect 33524 904 33525 944
rect 33483 895 33525 904
rect 33867 944 33909 953
rect 33867 904 33868 944
rect 33908 904 33909 944
rect 33867 895 33909 904
rect 34251 944 34293 953
rect 34251 904 34252 944
rect 34292 904 34293 944
rect 34251 895 34293 904
rect 34635 944 34677 953
rect 34635 904 34636 944
rect 34676 904 34677 944
rect 34635 895 34677 904
rect 35403 944 35445 953
rect 35403 904 35404 944
rect 35444 904 35445 944
rect 35403 895 35445 904
rect 35787 944 35829 953
rect 35787 904 35788 944
rect 35828 904 35829 944
rect 35787 895 35829 904
rect 36171 944 36213 953
rect 36171 904 36172 944
rect 36212 904 36213 944
rect 36171 895 36213 904
rect 36555 944 36597 953
rect 36555 904 36556 944
rect 36596 904 36597 944
rect 36555 895 36597 904
rect 36939 944 36981 953
rect 36939 904 36940 944
rect 36980 904 36981 944
rect 36939 895 36981 904
rect 37419 944 37461 953
rect 37419 904 37420 944
rect 37460 904 37461 944
rect 37419 895 37461 904
rect 37803 944 37845 953
rect 37803 904 37804 944
rect 37844 904 37845 944
rect 37803 895 37845 904
rect 38187 944 38229 953
rect 38187 904 38188 944
rect 38228 904 38229 944
rect 38187 895 38229 904
rect 38571 944 38613 953
rect 38571 904 38572 944
rect 38612 904 38613 944
rect 38571 895 38613 904
rect 38955 944 38997 953
rect 38955 904 38956 944
rect 38996 904 38997 944
rect 38955 895 38997 904
rect 39339 944 39381 953
rect 39339 904 39340 944
rect 39380 904 39381 944
rect 39339 895 39381 904
rect 39723 944 39765 953
rect 39723 904 39724 944
rect 39764 904 39765 944
rect 39723 895 39765 904
rect 40107 944 40149 953
rect 40107 904 40108 944
rect 40148 904 40149 944
rect 40107 895 40149 904
rect 40491 944 40533 953
rect 40491 904 40492 944
rect 40532 904 40533 944
rect 40491 895 40533 904
rect 40875 944 40917 953
rect 40875 904 40876 944
rect 40916 904 40917 944
rect 40875 895 40917 904
rect 41259 944 41301 953
rect 41259 904 41260 944
rect 41300 904 41301 944
rect 41259 895 41301 904
rect 41643 944 41685 953
rect 41643 904 41644 944
rect 41684 904 41685 944
rect 41643 895 41685 904
rect 42027 944 42069 953
rect 42027 904 42028 944
rect 42068 904 42069 944
rect 42027 895 42069 904
rect 42411 944 42453 953
rect 42411 904 42412 944
rect 42452 904 42453 944
rect 42411 895 42453 904
rect 42795 944 42837 953
rect 42795 904 42796 944
rect 42836 904 42837 944
rect 42795 895 42837 904
rect 43179 944 43221 953
rect 43179 904 43180 944
rect 43220 904 43221 944
rect 43179 895 43221 904
rect 43659 944 43701 953
rect 43659 904 43660 944
rect 43700 904 43701 944
rect 43659 895 43701 904
rect 44043 944 44085 953
rect 44043 904 44044 944
rect 44084 904 44085 944
rect 44043 895 44085 904
rect 44427 944 44469 953
rect 44427 904 44428 944
rect 44468 904 44469 944
rect 44427 895 44469 904
rect 44811 944 44853 953
rect 44811 904 44812 944
rect 44852 904 44853 944
rect 44811 895 44853 904
rect 45195 944 45237 953
rect 45195 904 45196 944
rect 45236 904 45237 944
rect 45195 895 45237 904
rect 45579 944 45621 953
rect 45579 904 45580 944
rect 45620 904 45621 944
rect 45579 895 45621 904
rect 45963 944 46005 953
rect 45963 904 45964 944
rect 46004 904 46005 944
rect 45963 895 46005 904
rect 46347 944 46389 953
rect 46347 904 46348 944
rect 46388 904 46389 944
rect 46347 895 46389 904
rect 46731 944 46773 953
rect 46731 904 46732 944
rect 46772 904 46773 944
rect 46731 895 46773 904
rect 47115 944 47157 953
rect 47115 904 47116 944
rect 47156 904 47157 944
rect 47115 895 47157 904
rect 47499 944 47541 953
rect 47499 904 47500 944
rect 47540 904 47541 944
rect 47499 895 47541 904
rect 47883 944 47925 953
rect 47883 904 47884 944
rect 47924 904 47925 944
rect 47883 895 47925 904
rect 48267 944 48309 953
rect 48267 904 48268 944
rect 48308 904 48309 944
rect 48267 895 48309 904
rect 48651 944 48693 953
rect 48651 904 48652 944
rect 48692 904 48693 944
rect 48651 895 48693 904
rect 49035 944 49077 953
rect 49035 904 49036 944
rect 49076 904 49077 944
rect 49035 895 49077 904
rect 49419 944 49461 953
rect 49419 904 49420 944
rect 49460 904 49461 944
rect 49419 895 49461 904
rect 50475 944 50517 953
rect 50475 904 50476 944
rect 50516 904 50517 944
rect 50475 895 50517 904
rect 50763 944 50805 953
rect 50763 904 50764 944
rect 50804 904 50805 944
rect 50763 895 50805 904
rect 51243 944 51285 953
rect 51243 904 51244 944
rect 51284 904 51285 944
rect 51243 895 51285 904
rect 52011 944 52053 953
rect 52011 904 52012 944
rect 52052 904 52053 944
rect 52011 895 52053 904
rect 52587 944 52629 953
rect 52587 904 52588 944
rect 52628 904 52629 944
rect 52587 895 52629 904
rect 53643 944 53685 953
rect 53643 904 53644 944
rect 53684 904 53685 944
rect 53643 895 53685 904
rect 53931 944 53973 953
rect 53931 904 53932 944
rect 53972 904 53973 944
rect 53931 895 53973 904
rect 54411 944 54453 953
rect 54411 904 54412 944
rect 54452 904 54453 944
rect 54411 895 54453 904
rect 54891 944 54933 953
rect 54891 904 54892 944
rect 54932 904 54933 944
rect 54891 895 54933 904
rect 55467 944 55509 953
rect 55467 904 55468 944
rect 55508 904 55509 944
rect 55467 895 55509 904
rect 56331 944 56373 953
rect 56331 904 56332 944
rect 56372 904 56373 944
rect 56331 895 56373 904
rect 56907 944 56949 953
rect 56907 904 56908 944
rect 56948 904 56949 944
rect 56907 895 56949 904
rect 57387 944 57429 953
rect 57387 904 57388 944
rect 57428 904 57429 944
rect 57387 895 57429 904
rect 57963 944 58005 953
rect 57963 904 57964 944
rect 58004 904 58005 944
rect 57963 895 58005 904
rect 58251 944 58293 953
rect 58251 904 58252 944
rect 58292 904 58293 944
rect 58251 895 58293 904
rect 59787 944 59829 953
rect 59787 904 59788 944
rect 59828 904 59829 944
rect 59787 895 59829 904
rect 59979 944 60021 953
rect 59979 904 59980 944
rect 60020 904 60021 944
rect 59979 895 60021 904
rect 60459 944 60501 953
rect 60459 904 60460 944
rect 60500 904 60501 944
rect 60459 895 60501 904
rect 61035 944 61077 953
rect 61035 904 61036 944
rect 61076 904 61077 944
rect 61035 895 61077 904
rect 62763 944 62805 953
rect 62763 904 62764 944
rect 62804 904 62805 944
rect 62763 895 62805 904
rect 63531 944 63573 953
rect 63531 904 63532 944
rect 63572 904 63573 944
rect 63531 895 63573 904
rect 63915 944 63957 953
rect 63915 904 63916 944
rect 63956 904 63957 944
rect 63915 895 63957 904
rect 64299 944 64341 953
rect 64299 904 64300 944
rect 64340 904 64341 944
rect 64299 895 64341 904
rect 64683 944 64725 953
rect 64683 904 64684 944
rect 64724 904 64725 944
rect 64683 895 64725 904
rect 65067 944 65109 953
rect 65067 904 65068 944
rect 65108 904 65109 944
rect 65067 895 65109 904
rect 65451 944 65493 953
rect 65451 904 65452 944
rect 65492 904 65493 944
rect 65451 895 65493 904
rect 65835 944 65877 953
rect 65835 904 65836 944
rect 65876 904 65877 944
rect 65835 895 65877 904
rect 66219 944 66261 953
rect 66219 904 66220 944
rect 66260 904 66261 944
rect 66219 895 66261 904
rect 67371 944 67413 953
rect 67371 904 67372 944
rect 67412 904 67413 944
rect 67371 895 67413 904
rect 68139 944 68181 953
rect 68139 904 68140 944
rect 68180 904 68181 944
rect 68139 895 68181 904
rect 68523 944 68565 953
rect 68523 904 68524 944
rect 68564 904 68565 944
rect 68523 895 68565 904
rect 68907 944 68949 953
rect 68907 904 68908 944
rect 68948 904 68949 944
rect 68907 895 68949 904
rect 69291 944 69333 953
rect 69291 904 69292 944
rect 69332 904 69333 944
rect 69291 895 69333 904
rect 69675 944 69717 953
rect 69675 904 69676 944
rect 69716 904 69717 944
rect 69675 895 69717 904
rect 70059 944 70101 953
rect 70059 904 70060 944
rect 70100 904 70101 944
rect 70059 895 70101 904
rect 70443 944 70485 953
rect 70443 904 70444 944
rect 70484 904 70485 944
rect 70443 895 70485 904
rect 71211 944 71253 953
rect 71211 904 71212 944
rect 71252 904 71253 944
rect 71211 895 71253 904
rect 71595 944 71637 953
rect 71595 904 71596 944
rect 71636 904 71637 944
rect 71595 895 71637 904
rect 71979 944 72021 953
rect 71979 904 71980 944
rect 72020 904 72021 944
rect 71979 895 72021 904
rect 72747 944 72789 953
rect 72747 904 72748 944
rect 72788 904 72789 944
rect 72747 895 72789 904
rect 73131 944 73173 953
rect 73131 904 73132 944
rect 73172 904 73173 944
rect 73131 895 73173 904
rect 73515 944 73557 953
rect 73515 904 73516 944
rect 73556 904 73557 944
rect 73515 895 73557 904
rect 73899 944 73941 953
rect 73899 904 73900 944
rect 73940 904 73941 944
rect 73899 895 73941 904
rect 74283 944 74325 953
rect 74283 904 74284 944
rect 74324 904 74325 944
rect 74283 895 74325 904
rect 74667 944 74709 953
rect 74667 904 74668 944
rect 74708 904 74709 944
rect 74667 895 74709 904
rect 75051 944 75093 953
rect 75051 904 75052 944
rect 75092 904 75093 944
rect 75051 895 75093 904
rect 75435 944 75477 953
rect 75435 904 75436 944
rect 75476 904 75477 944
rect 75435 895 75477 904
rect 75819 944 75861 953
rect 75819 904 75820 944
rect 75860 904 75861 944
rect 75819 895 75861 904
rect 76203 944 76245 953
rect 76203 904 76204 944
rect 76244 904 76245 944
rect 76203 895 76245 904
rect 76587 944 76629 953
rect 76587 904 76588 944
rect 76628 904 76629 944
rect 76587 895 76629 904
rect 76971 944 77013 953
rect 76971 904 76972 944
rect 77012 904 77013 944
rect 76971 895 77013 904
rect 77355 944 77397 953
rect 77355 904 77356 944
rect 77396 904 77397 944
rect 77355 895 77397 904
rect 77739 944 77781 953
rect 77739 904 77740 944
rect 77780 904 77781 944
rect 77739 895 77781 904
rect 78123 944 78165 953
rect 78123 904 78124 944
rect 78164 904 78165 944
rect 78123 895 78165 904
rect 78507 944 78549 953
rect 78507 904 78508 944
rect 78548 904 78549 944
rect 78507 895 78549 904
rect 78891 944 78933 953
rect 78891 904 78892 944
rect 78932 904 78933 944
rect 78891 895 78933 904
rect 79275 944 79317 953
rect 79275 904 79276 944
rect 79316 904 79317 944
rect 79275 895 79317 904
rect 79659 944 79701 953
rect 79659 904 79660 944
rect 79700 904 79701 944
rect 79659 895 79701 904
rect 80043 944 80085 953
rect 80043 904 80044 944
rect 80084 904 80085 944
rect 80043 895 80085 904
rect 80427 944 80469 953
rect 80427 904 80428 944
rect 80468 904 80469 944
rect 80427 895 80469 904
rect 81003 944 81045 953
rect 81003 904 81004 944
rect 81044 904 81045 944
rect 81003 895 81045 904
rect 81387 944 81429 953
rect 81387 904 81388 944
rect 81428 904 81429 944
rect 81387 895 81429 904
rect 81771 944 81813 953
rect 81771 904 81772 944
rect 81812 904 81813 944
rect 81771 895 81813 904
rect 82155 944 82197 953
rect 82155 904 82156 944
rect 82196 904 82197 944
rect 82155 895 82197 904
rect 82539 944 82581 953
rect 82539 904 82540 944
rect 82580 904 82581 944
rect 82539 895 82581 904
rect 83307 944 83349 953
rect 83307 904 83308 944
rect 83348 904 83349 944
rect 83307 895 83349 904
rect 83691 944 83733 953
rect 83691 904 83692 944
rect 83732 904 83733 944
rect 83691 895 83733 904
rect 84075 944 84117 953
rect 84075 904 84076 944
rect 84116 904 84117 944
rect 84075 895 84117 904
rect 84459 944 84501 953
rect 84459 904 84460 944
rect 84500 904 84501 944
rect 84459 895 84501 904
rect 84843 944 84885 953
rect 84843 904 84844 944
rect 84884 904 84885 944
rect 84843 895 84885 904
rect 85227 944 85269 953
rect 85227 904 85228 944
rect 85268 904 85269 944
rect 85227 895 85269 904
rect 86379 944 86421 953
rect 86379 904 86380 944
rect 86420 904 86421 944
rect 86379 895 86421 904
rect 86763 944 86805 953
rect 86763 904 86764 944
rect 86804 904 86805 944
rect 86763 895 86805 904
rect 87147 944 87189 953
rect 87147 904 87148 944
rect 87188 904 87189 944
rect 87147 895 87189 904
rect 87531 944 87573 953
rect 87531 904 87532 944
rect 87572 904 87573 944
rect 87531 895 87573 904
rect 87915 944 87957 953
rect 87915 904 87916 944
rect 87956 904 87957 944
rect 87915 895 87957 904
rect 88299 944 88341 953
rect 88299 904 88300 944
rect 88340 904 88341 944
rect 88299 895 88341 904
rect 88683 944 88725 953
rect 88683 904 88684 944
rect 88724 904 88725 944
rect 88683 895 88725 904
rect 89451 944 89493 953
rect 89451 904 89452 944
rect 89492 904 89493 944
rect 89451 895 89493 904
rect 89835 944 89877 953
rect 89835 904 89836 944
rect 89876 904 89877 944
rect 89835 895 89877 904
rect 90219 944 90261 953
rect 90219 904 90220 944
rect 90260 904 90261 944
rect 90219 895 90261 904
rect 90603 944 90645 953
rect 90603 904 90604 944
rect 90644 904 90645 944
rect 90603 895 90645 904
rect 90987 944 91029 953
rect 90987 904 90988 944
rect 91028 904 91029 944
rect 90987 895 91029 904
rect 91755 944 91797 953
rect 91755 904 91756 944
rect 91796 904 91797 944
rect 91755 895 91797 904
rect 92523 944 92565 953
rect 92523 904 92524 944
rect 92564 904 92565 944
rect 92523 895 92565 904
rect 92907 944 92949 953
rect 92907 904 92908 944
rect 92948 904 92949 944
rect 92907 895 92949 904
rect 93291 944 93333 953
rect 93291 904 93292 944
rect 93332 904 93333 944
rect 93291 895 93333 904
rect 93675 944 93717 953
rect 93675 904 93676 944
rect 93716 904 93717 944
rect 93675 895 93717 904
rect 94059 944 94101 953
rect 94059 904 94060 944
rect 94100 904 94101 944
rect 94059 895 94101 904
rect 94443 944 94485 953
rect 94443 904 94444 944
rect 94484 904 94485 944
rect 94443 895 94485 904
rect 94827 944 94869 953
rect 94827 904 94828 944
rect 94868 904 94869 944
rect 94827 895 94869 904
rect 95211 944 95253 953
rect 95211 904 95212 944
rect 95252 904 95253 944
rect 95211 895 95253 904
rect 95595 944 95637 953
rect 95595 904 95596 944
rect 95636 904 95637 944
rect 95595 895 95637 904
rect 95979 944 96021 953
rect 95979 904 95980 944
rect 96020 904 96021 944
rect 95979 895 96021 904
rect 96363 944 96405 953
rect 96363 904 96364 944
rect 96404 904 96405 944
rect 96363 895 96405 904
rect 96747 944 96789 953
rect 96747 904 96748 944
rect 96788 904 96789 944
rect 96747 895 96789 904
rect 97131 944 97173 953
rect 97131 904 97132 944
rect 97172 904 97173 944
rect 97131 895 97173 904
rect 97515 944 97557 953
rect 97515 904 97516 944
rect 97556 904 97557 944
rect 97515 895 97557 904
rect 98667 944 98709 953
rect 98667 904 98668 944
rect 98708 904 98709 944
rect 98667 895 98709 904
rect 99051 944 99093 953
rect 99051 904 99052 944
rect 99092 904 99093 944
rect 99051 895 99093 904
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 45772 6616 45812 6656
rect 48556 6616 48596 6656
rect 41740 6448 41780 6488
rect 42028 6448 42068 6488
rect 44524 6448 44564 6488
rect 44716 6448 44756 6488
rect 45868 6448 45908 6488
rect 46444 6448 46484 6488
rect 46540 6448 46580 6488
rect 47596 6448 47636 6488
rect 47884 6448 47924 6488
rect 48460 6448 48500 6488
rect 48748 6448 48788 6488
rect 49036 6448 49076 6488
rect 49228 6448 49268 6488
rect 49420 6448 49460 6488
rect 46636 6364 46676 6404
rect 48844 6364 48884 6404
rect 49324 6364 49364 6404
rect 41740 6280 41780 6320
rect 46732 6280 46772 6320
rect 46828 6280 46868 6320
rect 47596 6280 47636 6320
rect 48268 6280 48308 6320
rect 44524 6196 44564 6236
rect 46060 6196 46100 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 53452 5860 53492 5900
rect 41068 5608 41108 5648
rect 41356 5608 41396 5648
rect 41740 5608 41780 5648
rect 41836 5608 41876 5648
rect 44236 5608 44276 5648
rect 44332 5608 44372 5648
rect 44908 5608 44948 5648
rect 45004 5608 45044 5648
rect 46060 5608 46100 5648
rect 46252 5608 46292 5648
rect 46348 5608 46388 5648
rect 50476 5608 50516 5648
rect 50668 5608 50708 5648
rect 51916 5608 51956 5648
rect 52108 5608 52148 5648
rect 52492 5608 52532 5648
rect 52588 5608 52628 5648
rect 53644 5608 53684 5648
rect 53740 5608 53780 5648
rect 54316 5608 54356 5648
rect 54508 5608 54548 5648
rect 55468 5608 55508 5648
rect 55564 5608 55604 5648
rect 56332 5608 56372 5648
rect 56620 5608 56660 5648
rect 56812 5608 56852 5648
rect 58156 5608 58196 5648
rect 58348 5608 58388 5648
rect 61228 5608 61268 5648
rect 61324 5608 61364 5648
rect 61708 5608 61748 5648
rect 61804 5608 61844 5648
rect 61900 5608 61940 5648
rect 61996 5608 62036 5648
rect 41548 5524 41588 5564
rect 44044 5524 44084 5564
rect 44716 5524 44756 5564
rect 50572 5524 50612 5564
rect 52012 5524 52052 5564
rect 52300 5524 52340 5564
rect 54412 5524 54452 5564
rect 55276 5524 55316 5564
rect 56716 5524 56756 5564
rect 61132 5524 61172 5564
rect 41260 5440 41300 5480
rect 41836 5440 41876 5480
rect 44332 5440 44372 5480
rect 45004 5440 45044 5480
rect 46060 5440 46100 5480
rect 52588 5440 52628 5480
rect 53740 5440 53780 5480
rect 55564 5440 55604 5480
rect 56140 5440 56180 5480
rect 56428 5440 56468 5480
rect 58252 5440 58292 5480
rect 60940 5440 60980 5480
rect 61036 5440 61076 5480
rect 61516 5440 61556 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 41452 5104 41492 5144
rect 42124 5104 42164 5144
rect 45868 5104 45908 5144
rect 46636 5104 46676 5144
rect 48076 5104 48116 5144
rect 48844 5104 48884 5144
rect 56620 5104 56660 5144
rect 58060 5104 58100 5144
rect 58732 5104 58772 5144
rect 61900 5104 61940 5144
rect 62188 5020 62228 5060
rect 22444 4936 22484 4976
rect 41356 4936 41396 4976
rect 41452 4936 41492 4976
rect 42028 4936 42068 4976
rect 42124 4936 42164 4976
rect 45868 4936 45908 4976
rect 45964 4936 46004 4976
rect 46540 4936 46580 4976
rect 46636 4936 46676 4976
rect 48076 4936 48116 4976
rect 48172 4936 48212 4976
rect 48748 4936 48788 4976
rect 48844 4936 48884 4976
rect 49324 4936 49364 4976
rect 49516 4936 49556 4976
rect 49612 4936 49652 4976
rect 50380 4936 50420 4976
rect 50668 4936 50708 4976
rect 50860 4947 50900 4987
rect 52396 4936 52436 4976
rect 52685 4947 52725 4987
rect 52876 4936 52916 4976
rect 53548 4936 53588 4976
rect 53740 4936 53780 4976
rect 54892 4936 54932 4976
rect 55180 4936 55220 4976
rect 55372 4936 55412 4976
rect 55948 4936 55988 4976
rect 56140 4936 56180 4976
rect 56332 4936 56372 4976
rect 56428 4936 56468 4976
rect 57964 4936 58004 4976
rect 58060 4936 58100 4976
rect 58636 4936 58676 4976
rect 58732 4936 58772 4976
rect 60460 4936 60500 4976
rect 60844 4936 60884 4976
rect 61036 4936 61076 4976
rect 61228 4936 61268 4976
rect 61324 4936 61364 4976
rect 61516 4936 61556 4976
rect 61900 4936 61940 4976
rect 61996 4936 62036 4976
rect 62380 4936 62420 4976
rect 62572 4936 62612 4976
rect 62668 4936 62708 4976
rect 66892 4936 66932 4976
rect 67180 4936 67220 4976
rect 73324 4936 73364 4976
rect 73612 4936 73652 4976
rect 73804 4936 73844 4976
rect 74092 4936 74132 4976
rect 74284 4936 74324 4976
rect 74476 4936 74516 4976
rect 82156 4936 82196 4976
rect 82348 4936 82388 4976
rect 50764 4852 50804 4892
rect 56044 4852 56084 4892
rect 74380 4852 74420 4892
rect 48556 4768 48596 4808
rect 50380 4768 50420 4808
rect 52396 4768 52436 4808
rect 54892 4768 54932 4808
rect 60460 4768 60500 4808
rect 22348 4684 22388 4724
rect 41164 4684 41204 4724
rect 41836 4684 41876 4724
rect 46156 4684 46196 4724
rect 46348 4684 46388 4724
rect 48364 4684 48404 4724
rect 49516 4684 49556 4724
rect 50188 4684 50228 4724
rect 52204 4684 52244 4724
rect 52684 4684 52724 4724
rect 53644 4684 53684 4724
rect 54700 4684 54740 4724
rect 55180 4684 55220 4724
rect 57772 4684 57812 4724
rect 58444 4684 58484 4724
rect 60652 4684 60692 4724
rect 60844 4684 60884 4724
rect 61324 4684 61364 4724
rect 62380 4684 62420 4724
rect 67180 4684 67220 4724
rect 73324 4684 73364 4724
rect 74092 4684 74132 4724
rect 82156 4684 82196 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 38668 4348 38708 4388
rect 43084 4348 43124 4388
rect 52300 4348 52340 4388
rect 7564 4264 7604 4304
rect 53356 4264 53396 4304
rect 58156 4264 58196 4304
rect 59020 4264 59060 4304
rect 6988 4096 7028 4136
rect 7180 4096 7220 4136
rect 7564 4096 7604 4136
rect 18316 4096 18356 4136
rect 18412 4096 18452 4136
rect 18988 4096 19028 4136
rect 19084 4127 19124 4167
rect 19468 4096 19508 4136
rect 19660 4096 19700 4136
rect 19756 4096 19796 4136
rect 24364 4096 24404 4136
rect 24460 4096 24500 4136
rect 24844 4096 24884 4136
rect 25036 4096 25076 4136
rect 25132 4096 25172 4136
rect 25900 4096 25940 4136
rect 26092 4096 26132 4136
rect 27916 4096 27956 4136
rect 28012 4096 28052 4136
rect 32140 4096 32180 4136
rect 32236 4096 32276 4136
rect 32620 4096 32660 4136
rect 32812 4096 32852 4136
rect 32908 4096 32948 4136
rect 37228 4096 37268 4136
rect 37324 4096 37364 4136
rect 37708 4096 37748 4136
rect 37804 4096 37844 4136
rect 37996 4096 38036 4136
rect 38380 4096 38420 4136
rect 38476 4096 38516 4136
rect 41260 4096 41300 4136
rect 41548 4138 41588 4178
rect 41452 4096 41492 4136
rect 41932 4096 41972 4136
rect 42028 4096 42068 4136
rect 42412 4096 42452 4136
rect 42604 4096 42644 4136
rect 42700 4096 42740 4136
rect 42892 4096 42932 4136
rect 43084 4096 43124 4136
rect 43180 4096 43220 4136
rect 44332 4096 44372 4136
rect 44620 4138 44660 4178
rect 44524 4096 44564 4136
rect 44812 4096 44852 4136
rect 45004 4096 45044 4136
rect 45100 4096 45140 4136
rect 46060 4096 46100 4136
rect 46252 4096 46292 4136
rect 46348 4096 46388 4136
rect 48172 4096 48212 4136
rect 48364 4096 48404 4136
rect 48460 4096 48500 4136
rect 48652 4096 48692 4136
rect 48844 4096 48884 4136
rect 48940 4096 48980 4136
rect 50188 4096 50228 4136
rect 50380 4096 50420 4136
rect 50572 4096 50612 4136
rect 50764 4096 50804 4136
rect 51244 4096 51284 4136
rect 51436 4096 51476 4136
rect 51532 4096 51572 4136
rect 52204 4096 52244 4136
rect 52396 4111 52436 4151
rect 52588 4111 52628 4151
rect 52780 4096 52820 4136
rect 53356 4096 53396 4136
rect 53644 4096 53684 4136
rect 53836 4096 53876 4136
rect 55084 4096 55124 4136
rect 55276 4096 55316 4136
rect 55372 4096 55412 4136
rect 58156 4096 58196 4136
rect 58540 4096 58580 4136
rect 58732 4096 58772 4136
rect 59020 4096 59060 4136
rect 59404 4096 59444 4136
rect 59596 4096 59636 4136
rect 61516 4096 61556 4136
rect 61900 4096 61940 4136
rect 62284 4096 62324 4136
rect 62476 4096 62516 4136
rect 66508 4096 66548 4136
rect 66796 4096 66836 4136
rect 66988 4096 67028 4136
rect 68524 4096 68564 4136
rect 68908 4096 68948 4136
rect 69100 4096 69140 4136
rect 74092 4096 74132 4136
rect 74284 4096 74324 4136
rect 74380 4096 74420 4136
rect 74764 4096 74804 4136
rect 74860 4096 74900 4136
rect 80332 4096 80372 4136
rect 80524 4096 80564 4136
rect 80812 4096 80852 4136
rect 86668 4096 86708 4136
rect 87052 4096 87092 4136
rect 87244 4096 87284 4136
rect 91564 4096 91604 4136
rect 91756 4096 91796 4136
rect 92044 4096 92084 4136
rect 18124 4012 18164 4052
rect 18796 4012 18836 4052
rect 24652 4012 24692 4052
rect 31948 4012 31988 4052
rect 37516 4012 37556 4052
rect 41740 4012 41780 4052
rect 50284 4012 50324 4052
rect 50668 4012 50708 4052
rect 52684 4012 52724 4052
rect 58636 4012 58676 4052
rect 62380 4012 62420 4052
rect 66892 4012 66932 4052
rect 69004 4012 69044 4052
rect 75052 4012 75092 4052
rect 80428 4012 80468 4052
rect 87148 4012 87188 4052
rect 91660 4012 91700 4052
rect 7084 3928 7124 3968
rect 7372 3928 7412 3968
rect 18412 3928 18452 3968
rect 19084 3928 19124 3968
rect 19468 3928 19508 3968
rect 24364 3928 24404 3968
rect 24844 3928 24884 3968
rect 25996 3928 26036 3968
rect 27724 3928 27764 3968
rect 32236 3928 32276 3968
rect 32620 3928 32660 3968
rect 37228 3928 37268 3968
rect 37996 3928 38036 3968
rect 38380 3928 38420 3968
rect 41260 3928 41300 3968
rect 42028 3928 42068 3968
rect 42412 3928 42452 3968
rect 44332 3928 44372 3968
rect 44812 3928 44852 3968
rect 46060 3928 46100 3968
rect 48172 3928 48212 3968
rect 48652 3928 48692 3968
rect 51244 3928 51284 3968
rect 53164 3928 53204 3968
rect 53740 3928 53780 3968
rect 55084 3928 55124 3968
rect 58348 3928 58388 3968
rect 59212 3928 59252 3968
rect 59500 3928 59540 3968
rect 61324 3928 61364 3968
rect 61612 3928 61652 3968
rect 61804 3928 61844 3968
rect 62092 3928 62132 3968
rect 66316 3928 66356 3968
rect 66604 3928 66644 3968
rect 68428 3928 68468 3968
rect 68716 3928 68756 3968
rect 74092 3928 74132 3968
rect 74764 3928 74804 3968
rect 80716 3928 80756 3968
rect 81004 3928 81044 3968
rect 86572 3928 86612 3968
rect 86860 3928 86900 3968
rect 91948 3928 91988 3968
rect 92236 3928 92276 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 33676 3508 33716 3548
rect 1900 3424 1940 3464
rect 2092 3424 2132 3464
rect 4204 3424 4244 3464
rect 4396 3424 4436 3464
rect 4588 3424 4628 3464
rect 4780 3424 4820 3464
rect 4972 3424 5012 3464
rect 5164 3424 5204 3464
rect 5740 3424 5780 3464
rect 5932 3424 5972 3464
rect 6892 3424 6932 3464
rect 7084 3424 7124 3464
rect 7276 3445 7316 3485
rect 7468 3424 7508 3464
rect 7660 3424 7700 3464
rect 7852 3424 7892 3464
rect 8428 3424 8468 3464
rect 8620 3424 8660 3464
rect 8812 3424 8852 3464
rect 9004 3424 9044 3464
rect 9196 3424 9236 3464
rect 9388 3424 9428 3464
rect 9580 3424 9620 3464
rect 9772 3424 9812 3464
rect 9964 3424 10004 3464
rect 10156 3424 10196 3464
rect 10348 3424 10388 3464
rect 10540 3424 10580 3464
rect 10732 3424 10772 3464
rect 10924 3424 10964 3464
rect 11116 3424 11156 3464
rect 11308 3424 11348 3464
rect 11500 3424 11540 3464
rect 11692 3424 11732 3464
rect 11884 3424 11924 3464
rect 12076 3424 12116 3464
rect 12268 3424 12308 3464
rect 12460 3424 12500 3464
rect 13036 3424 13076 3464
rect 13228 3424 13268 3464
rect 13420 3424 13460 3464
rect 13612 3424 13652 3464
rect 13804 3424 13844 3464
rect 13996 3424 14036 3464
rect 14284 3424 14324 3464
rect 14476 3424 14516 3464
rect 14668 3424 14708 3464
rect 14860 3424 14900 3464
rect 15052 3424 15092 3464
rect 15244 3424 15284 3464
rect 15436 3424 15476 3464
rect 15628 3424 15668 3464
rect 15820 3424 15860 3464
rect 16012 3424 16052 3464
rect 16204 3424 16244 3464
rect 16396 3424 16436 3464
rect 16588 3424 16628 3464
rect 16780 3424 16820 3464
rect 16972 3424 17012 3464
rect 17164 3424 17204 3464
rect 17356 3424 17396 3464
rect 17548 3424 17588 3464
rect 17740 3424 17780 3464
rect 17932 3424 17972 3464
rect 18124 3424 18164 3464
rect 18316 3424 18356 3464
rect 18508 3424 18548 3464
rect 18700 3424 18740 3464
rect 18892 3424 18932 3464
rect 19084 3424 19124 3464
rect 19180 3424 19220 3464
rect 19948 3424 19988 3464
rect 20149 3409 20189 3449
rect 20716 3424 20756 3464
rect 20908 3424 20948 3464
rect 21100 3424 21140 3464
rect 21292 3424 21332 3464
rect 21484 3424 21524 3464
rect 21676 3424 21716 3464
rect 22156 3424 22196 3464
rect 22348 3424 22388 3464
rect 22540 3424 22580 3464
rect 22732 3424 22772 3464
rect 22924 3424 22964 3464
rect 23116 3424 23156 3464
rect 23596 3424 23636 3464
rect 23788 3424 23828 3464
rect 23980 3424 24020 3464
rect 24172 3424 24212 3464
rect 24364 3424 24404 3464
rect 24556 3424 24596 3464
rect 25324 3424 25364 3464
rect 25516 3424 25556 3464
rect 25708 3424 25748 3464
rect 25900 3424 25940 3464
rect 26092 3424 26132 3464
rect 26284 3424 26324 3464
rect 26764 3424 26804 3464
rect 26956 3424 26996 3464
rect 27148 3424 27188 3464
rect 27340 3424 27380 3464
rect 27628 3424 27668 3464
rect 27820 3424 27860 3464
rect 28396 3424 28436 3464
rect 28588 3424 28628 3464
rect 28780 3424 28820 3464
rect 28972 3424 29012 3464
rect 29164 3424 29204 3464
rect 29356 3424 29396 3464
rect 29644 3424 29684 3464
rect 29836 3424 29876 3464
rect 30028 3424 30068 3464
rect 30220 3424 30260 3464
rect 30412 3424 30452 3464
rect 30604 3424 30644 3464
rect 31276 3424 31316 3464
rect 31468 3424 31508 3464
rect 31660 3424 31700 3464
rect 31852 3424 31892 3464
rect 32044 3424 32084 3464
rect 32236 3424 32276 3464
rect 32428 3424 32468 3464
rect 32620 3424 32660 3464
rect 32812 3424 32852 3464
rect 33004 3424 33044 3464
rect 33196 3424 33236 3464
rect 33388 3424 33428 3464
rect 33580 3424 33620 3464
rect 33772 3424 33812 3464
rect 33964 3424 34004 3464
rect 34156 3424 34196 3464
rect 34348 3424 34388 3464
rect 34540 3424 34580 3464
rect 34732 3424 34772 3464
rect 34924 3424 34964 3464
rect 35116 3424 35156 3464
rect 35308 3424 35348 3464
rect 35500 3424 35540 3464
rect 35692 3424 35732 3464
rect 35884 3424 35924 3464
rect 36076 3424 36116 3464
rect 36268 3424 36308 3464
rect 36460 3424 36500 3464
rect 36652 3424 36692 3464
rect 36844 3424 36884 3464
rect 37804 3424 37844 3464
rect 37996 3424 38036 3464
rect 38092 3424 38132 3464
rect 38284 3424 38324 3464
rect 38476 3424 38516 3464
rect 38860 3424 38900 3464
rect 39052 3424 39092 3464
rect 39244 3424 39284 3464
rect 39436 3424 39476 3464
rect 39628 3424 39668 3464
rect 39820 3424 39860 3464
rect 40300 3424 40340 3464
rect 40492 3424 40532 3464
rect 40780 3424 40820 3464
rect 40972 3424 41012 3464
rect 41164 3424 41204 3464
rect 41356 3424 41396 3464
rect 41932 3424 41972 3464
rect 42124 3424 42164 3464
rect 42316 3424 42356 3464
rect 42508 3424 42548 3464
rect 42604 3424 42644 3464
rect 42796 3424 42836 3464
rect 42988 3424 43028 3464
rect 44428 3424 44468 3464
rect 44620 3424 44660 3464
rect 45196 3424 45236 3464
rect 45388 3424 45428 3464
rect 45580 3424 45620 3464
rect 45772 3424 45812 3464
rect 45964 3424 46004 3464
rect 46156 3424 46196 3464
rect 46828 3424 46868 3464
rect 47020 3424 47060 3464
rect 47212 3424 47252 3464
rect 47404 3424 47444 3464
rect 47596 3424 47636 3464
rect 47788 3424 47828 3464
rect 48940 3424 48980 3464
rect 49132 3424 49172 3464
rect 50092 3424 50132 3464
rect 50284 3424 50324 3464
rect 50668 3424 50708 3464
rect 50956 3424 50996 3464
rect 51148 3424 51188 3464
rect 52588 3424 52628 3464
rect 52780 3424 52820 3464
rect 53260 3424 53300 3464
rect 53452 3424 53492 3464
rect 54892 3424 54932 3464
rect 55084 3424 55124 3464
rect 55276 3424 55316 3464
rect 55468 3424 55508 3464
rect 56620 3424 56660 3464
rect 56908 3424 56948 3464
rect 57100 3424 57140 3464
rect 58156 3424 58196 3464
rect 58348 3424 58388 3464
rect 58540 3411 58580 3451
rect 58636 3424 58676 3464
rect 58828 3424 58868 3464
rect 59020 3424 59060 3464
rect 59116 3424 59156 3464
rect 59308 3424 59348 3464
rect 61612 3424 61652 3464
rect 61804 3424 61844 3464
rect 63148 3424 63188 3464
rect 63340 3424 63380 3464
rect 63820 3424 63860 3464
rect 64012 3424 64052 3464
rect 64204 3424 64244 3464
rect 64396 3424 64436 3464
rect 64588 3424 64628 3464
rect 64780 3424 64820 3464
rect 65260 3424 65300 3464
rect 65452 3424 65492 3464
rect 65644 3424 65684 3464
rect 65836 3424 65876 3464
rect 66028 3424 66068 3464
rect 66220 3424 66260 3464
rect 66796 3424 66836 3464
rect 66988 3424 67028 3464
rect 67180 3424 67220 3464
rect 67372 3424 67412 3464
rect 68620 3424 68660 3464
rect 68812 3424 68852 3464
rect 69004 3424 69044 3464
rect 69196 3424 69236 3464
rect 69388 3424 69428 3464
rect 69580 3424 69620 3464
rect 69772 3424 69812 3464
rect 69964 3424 70004 3464
rect 70156 3424 70196 3464
rect 70348 3424 70388 3464
rect 70540 3424 70580 3464
rect 70732 3424 70772 3464
rect 70924 3424 70964 3464
rect 71116 3424 71156 3464
rect 71308 3424 71348 3464
rect 71500 3424 71540 3464
rect 71692 3424 71732 3464
rect 71884 3424 71924 3464
rect 72076 3424 72116 3464
rect 72268 3424 72308 3464
rect 72460 3424 72500 3464
rect 72652 3424 72692 3464
rect 72844 3424 72884 3464
rect 73036 3424 73076 3464
rect 74956 3424 74996 3464
rect 75148 3424 75188 3464
rect 75340 3424 75380 3464
rect 75532 3424 75572 3464
rect 76012 3424 76052 3464
rect 76204 3424 76244 3464
rect 76396 3424 76436 3464
rect 76588 3424 76628 3464
rect 76780 3424 76820 3464
rect 76972 3424 77012 3464
rect 77452 3424 77492 3464
rect 77644 3424 77684 3464
rect 77932 3424 77972 3464
rect 78124 3424 78164 3464
rect 78316 3424 78356 3464
rect 78508 3424 78548 3464
rect 78988 3424 79028 3464
rect 79180 3424 79220 3464
rect 79372 3424 79412 3464
rect 79564 3424 79604 3464
rect 79756 3424 79796 3464
rect 79948 3424 79988 3464
rect 80140 3424 80180 3464
rect 80332 3424 80372 3464
rect 81100 3424 81140 3464
rect 81292 3424 81332 3464
rect 81484 3424 81524 3464
rect 81676 3424 81716 3464
rect 82156 3424 82196 3464
rect 82348 3424 82388 3464
rect 82540 3424 82580 3464
rect 82732 3424 82772 3464
rect 82924 3424 82964 3464
rect 83116 3424 83156 3464
rect 83596 3424 83636 3464
rect 83788 3424 83828 3464
rect 83980 3424 84020 3464
rect 84172 3424 84212 3464
rect 84364 3424 84404 3464
rect 84556 3424 84596 3464
rect 86860 3424 86900 3464
rect 87052 3424 87092 3464
rect 87244 3424 87284 3464
rect 87436 3424 87476 3464
rect 87628 3424 87668 3464
rect 87820 3424 87860 3464
rect 88012 3424 88052 3464
rect 88204 3424 88244 3464
rect 88396 3424 88436 3464
rect 88588 3424 88628 3464
rect 88780 3424 88820 3464
rect 88972 3424 89012 3464
rect 89164 3424 89204 3464
rect 89356 3424 89396 3464
rect 89548 3424 89588 3464
rect 89740 3424 89780 3464
rect 89932 3424 89972 3464
rect 90124 3424 90164 3464
rect 90316 3424 90356 3464
rect 90508 3424 90548 3464
rect 90700 3424 90740 3464
rect 90892 3424 90932 3464
rect 91084 3424 91124 3464
rect 91276 3424 91316 3464
rect 91468 3424 91508 3464
rect 91660 3424 91700 3464
rect 91852 3424 91892 3464
rect 92044 3424 92084 3464
rect 92236 3424 92276 3464
rect 92428 3424 92468 3464
rect 92620 3424 92660 3464
rect 92812 3424 92852 3464
rect 93292 3424 93332 3464
rect 93484 3424 93524 3464
rect 94060 3424 94100 3464
rect 94252 3424 94292 3464
rect 94444 3424 94484 3464
rect 94636 3424 94676 3464
rect 94828 3424 94868 3464
rect 95020 3424 95060 3464
rect 95500 3424 95540 3464
rect 95692 3424 95732 3464
rect 95980 3424 96020 3464
rect 96172 3424 96212 3464
rect 50668 3256 50708 3296
rect 52684 3256 52724 3296
rect 56620 3256 56660 3296
rect 1996 3172 2036 3212
rect 4300 3172 4340 3212
rect 4684 3172 4724 3212
rect 5068 3172 5108 3212
rect 5836 3172 5876 3212
rect 6988 3172 7028 3212
rect 7372 3172 7412 3212
rect 7756 3172 7796 3212
rect 8524 3172 8564 3212
rect 8908 3172 8948 3212
rect 9292 3172 9332 3212
rect 9676 3172 9716 3212
rect 10060 3172 10100 3212
rect 10444 3172 10484 3212
rect 10828 3172 10868 3212
rect 11212 3172 11252 3212
rect 11596 3172 11636 3212
rect 11980 3172 12020 3212
rect 12364 3172 12404 3212
rect 13132 3172 13172 3212
rect 13516 3172 13556 3212
rect 13900 3172 13940 3212
rect 14380 3172 14420 3212
rect 14764 3172 14804 3212
rect 15148 3172 15188 3212
rect 15532 3172 15572 3212
rect 15916 3172 15956 3212
rect 16300 3172 16340 3212
rect 16684 3172 16724 3212
rect 17068 3172 17108 3212
rect 17452 3172 17492 3212
rect 17836 3172 17876 3212
rect 18220 3172 18260 3212
rect 18604 3172 18644 3212
rect 18892 3172 18932 3212
rect 20044 3172 20084 3212
rect 20812 3172 20852 3212
rect 21196 3172 21236 3212
rect 21580 3172 21620 3212
rect 22252 3172 22292 3212
rect 22636 3172 22676 3212
rect 23020 3172 23060 3212
rect 23692 3172 23732 3212
rect 24076 3172 24116 3212
rect 24460 3172 24500 3212
rect 25420 3172 25460 3212
rect 25804 3172 25844 3212
rect 26188 3172 26228 3212
rect 26860 3172 26900 3212
rect 27244 3172 27284 3212
rect 27724 3172 27764 3212
rect 28492 3172 28532 3212
rect 28876 3172 28916 3212
rect 29260 3172 29300 3212
rect 29740 3172 29780 3212
rect 30124 3172 30164 3212
rect 30508 3172 30548 3212
rect 31372 3172 31412 3212
rect 31756 3172 31796 3212
rect 32140 3172 32180 3212
rect 32524 3172 32564 3212
rect 32908 3172 32948 3212
rect 33292 3172 33332 3212
rect 34060 3172 34100 3212
rect 34444 3172 34484 3212
rect 34828 3172 34868 3212
rect 35212 3172 35252 3212
rect 35596 3172 35636 3212
rect 35980 3172 36020 3212
rect 36364 3172 36404 3212
rect 36748 3172 36788 3212
rect 37804 3172 37844 3212
rect 38380 3172 38420 3212
rect 38956 3172 38996 3212
rect 39340 3172 39380 3212
rect 39724 3172 39764 3212
rect 40396 3172 40436 3212
rect 40876 3172 40916 3212
rect 41260 3172 41300 3212
rect 42028 3172 42068 3212
rect 42316 3172 42356 3212
rect 42892 3172 42932 3212
rect 44524 3172 44564 3212
rect 45292 3172 45332 3212
rect 45676 3172 45716 3212
rect 46060 3172 46100 3212
rect 46924 3172 46964 3212
rect 47308 3172 47348 3212
rect 47692 3172 47732 3212
rect 49036 3172 49076 3212
rect 50284 3172 50324 3212
rect 50476 3172 50516 3212
rect 51052 3172 51092 3212
rect 53356 3172 53396 3212
rect 54988 3172 55028 3212
rect 55372 3172 55412 3212
rect 56428 3172 56468 3212
rect 56908 3172 56948 3212
rect 58252 3172 58292 3212
rect 58828 3172 58868 3212
rect 59308 3172 59348 3212
rect 61708 3172 61748 3212
rect 63244 3172 63284 3212
rect 63916 3172 63956 3212
rect 64300 3172 64340 3212
rect 64684 3172 64724 3212
rect 65356 3172 65396 3212
rect 65740 3172 65780 3212
rect 66124 3172 66164 3212
rect 66892 3172 66932 3212
rect 67276 3172 67316 3212
rect 68716 3172 68756 3212
rect 69100 3172 69140 3212
rect 69484 3172 69524 3212
rect 69868 3172 69908 3212
rect 70252 3172 70292 3212
rect 70636 3172 70676 3212
rect 71020 3172 71060 3212
rect 71404 3172 71444 3212
rect 71788 3172 71828 3212
rect 72172 3172 72212 3212
rect 72556 3172 72596 3212
rect 72940 3172 72980 3212
rect 75052 3172 75092 3212
rect 75436 3172 75476 3212
rect 76108 3172 76148 3212
rect 76492 3172 76532 3212
rect 76876 3172 76916 3212
rect 77548 3172 77588 3212
rect 78028 3172 78068 3212
rect 78412 3172 78452 3212
rect 79084 3172 79124 3212
rect 79468 3172 79508 3212
rect 79852 3172 79892 3212
rect 80236 3172 80276 3212
rect 81196 3172 81236 3212
rect 81580 3172 81620 3212
rect 82252 3172 82292 3212
rect 82636 3172 82676 3212
rect 83020 3172 83060 3212
rect 83692 3172 83732 3212
rect 84076 3172 84116 3212
rect 84460 3172 84500 3212
rect 86956 3172 86996 3212
rect 87340 3172 87380 3212
rect 87724 3172 87764 3212
rect 88108 3172 88148 3212
rect 88492 3172 88532 3212
rect 88876 3172 88916 3212
rect 89260 3172 89300 3212
rect 89644 3172 89684 3212
rect 90028 3172 90068 3212
rect 90412 3172 90452 3212
rect 90796 3172 90836 3212
rect 91180 3172 91220 3212
rect 91564 3172 91604 3212
rect 91948 3172 91988 3212
rect 92332 3172 92372 3212
rect 92716 3172 92756 3212
rect 93388 3172 93428 3212
rect 94156 3172 94196 3212
rect 94540 3172 94580 3212
rect 94924 3172 94964 3212
rect 95596 3172 95636 3212
rect 96076 3172 96116 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 54892 2752 54932 2792
rect 55276 2726 55316 2766
rect 55756 2752 55796 2792
rect 58636 2752 58676 2792
rect 60940 2752 60980 2792
rect 61420 2752 61460 2792
rect 1612 2584 1652 2624
rect 1804 2584 1844 2624
rect 2092 2584 2132 2624
rect 2284 2584 2324 2624
rect 2476 2584 2516 2624
rect 2668 2584 2708 2624
rect 2956 2584 2996 2624
rect 3148 2584 3188 2624
rect 3340 2584 3380 2624
rect 3532 2584 3572 2624
rect 3724 2584 3764 2624
rect 3916 2584 3956 2624
rect 6124 2584 6164 2624
rect 6316 2584 6356 2624
rect 6604 2584 6644 2624
rect 6796 2584 6836 2624
rect 6988 2584 7028 2624
rect 7180 2584 7220 2624
rect 8044 2584 8084 2624
rect 8236 2584 8276 2624
rect 12556 2584 12596 2624
rect 12748 2584 12788 2624
rect 14092 2584 14132 2624
rect 14284 2584 14324 2624
rect 19660 2584 19700 2624
rect 19852 2584 19892 2624
rect 20236 2584 20276 2624
rect 20428 2584 20468 2624
rect 21868 2584 21908 2624
rect 22060 2584 22100 2624
rect 23404 2584 23444 2624
rect 23596 2584 23636 2624
rect 26380 2584 26420 2624
rect 26572 2584 26612 2624
rect 27916 2584 27956 2624
rect 28108 2584 28148 2624
rect 29548 2584 29588 2624
rect 29740 2584 29780 2624
rect 30700 2584 30740 2624
rect 30892 2584 30932 2624
rect 31660 2584 31700 2624
rect 31852 2584 31892 2624
rect 37612 2584 37652 2624
rect 37804 2584 37844 2624
rect 38188 2571 38228 2611
rect 38380 2584 38420 2624
rect 38572 2584 38612 2624
rect 38764 2584 38804 2624
rect 40012 2584 40052 2624
rect 40204 2584 40244 2624
rect 41644 2584 41684 2624
rect 41836 2584 41876 2624
rect 42028 2584 42068 2624
rect 42220 2584 42260 2624
rect 42796 2584 42836 2624
rect 42988 2584 43028 2624
rect 44044 2584 44084 2624
rect 44236 2584 44276 2624
rect 44812 2584 44852 2624
rect 45004 2584 45044 2624
rect 46348 2584 46388 2624
rect 46540 2584 46580 2624
rect 47884 2584 47924 2624
rect 48076 2584 48116 2624
rect 48268 2584 48308 2624
rect 48460 2584 48500 2624
rect 48652 2584 48692 2624
rect 48844 2584 48884 2624
rect 49132 2584 49172 2624
rect 49324 2584 49364 2624
rect 54700 2584 54740 2624
rect 54892 2573 54932 2613
rect 55276 2576 55316 2616
rect 55756 2584 55796 2624
rect 56044 2584 56084 2624
rect 56236 2584 56276 2624
rect 58636 2584 58676 2624
rect 60460 2584 60500 2624
rect 60652 2584 60692 2624
rect 60940 2584 60980 2624
rect 61420 2584 61460 2624
rect 61804 2584 61844 2624
rect 61996 2584 62036 2624
rect 62860 2584 62900 2624
rect 63052 2584 63092 2624
rect 63340 2584 63380 2624
rect 63532 2584 63572 2624
rect 67372 2584 67412 2624
rect 67564 2584 67604 2624
rect 72940 2584 72980 2624
rect 73132 2584 73172 2624
rect 73324 2584 73364 2624
rect 73516 2584 73556 2624
rect 73708 2584 73748 2624
rect 73901 2607 73941 2647
rect 74092 2584 74132 2624
rect 74284 2563 74324 2603
rect 74764 2584 74804 2624
rect 74956 2584 74996 2624
rect 75628 2584 75668 2624
rect 75820 2584 75860 2624
rect 77068 2584 77108 2624
rect 77260 2584 77300 2624
rect 78604 2584 78644 2624
rect 78796 2584 78836 2624
rect 81676 2584 81716 2624
rect 81868 2584 81908 2624
rect 83212 2584 83252 2624
rect 83404 2584 83444 2624
rect 84748 2584 84788 2624
rect 84940 2584 84980 2624
rect 85132 2584 85172 2624
rect 85324 2584 85364 2624
rect 85516 2584 85556 2624
rect 85708 2584 85748 2624
rect 85900 2584 85940 2624
rect 86092 2584 86132 2624
rect 86284 2584 86324 2624
rect 86476 2584 86516 2624
rect 92908 2584 92948 2624
rect 93100 2584 93140 2624
rect 93580 2584 93620 2624
rect 93772 2584 93812 2624
rect 95116 2584 95156 2624
rect 95308 2584 95348 2624
rect 96364 2584 96404 2624
rect 96556 2584 96596 2624
rect 96748 2584 96788 2624
rect 96940 2584 96980 2624
rect 97132 2584 97172 2624
rect 97324 2584 97364 2624
rect 97516 2584 97556 2624
rect 97709 2607 97749 2647
rect 97900 2584 97940 2624
rect 98092 2584 98132 2624
rect 1708 2500 1748 2540
rect 2188 2500 2228 2540
rect 2572 2500 2612 2540
rect 3052 2500 3092 2540
rect 3436 2500 3476 2540
rect 3820 2500 3860 2540
rect 6220 2500 6260 2540
rect 6700 2500 6740 2540
rect 7084 2500 7124 2540
rect 8140 2500 8180 2540
rect 12652 2500 12692 2540
rect 14188 2500 14228 2540
rect 19756 2500 19796 2540
rect 20332 2500 20372 2540
rect 21964 2500 22004 2540
rect 23500 2500 23540 2540
rect 26476 2500 26516 2540
rect 28012 2500 28052 2540
rect 29644 2500 29684 2540
rect 30796 2500 30836 2540
rect 31756 2500 31796 2540
rect 37708 2500 37748 2540
rect 38284 2500 38324 2540
rect 38668 2500 38708 2540
rect 40108 2500 40148 2540
rect 41740 2500 41780 2540
rect 42124 2500 42164 2540
rect 42892 2500 42932 2540
rect 44140 2500 44180 2540
rect 44908 2500 44948 2540
rect 46444 2500 46484 2540
rect 47980 2500 48020 2540
rect 48364 2500 48404 2540
rect 48748 2500 48788 2540
rect 49228 2500 49268 2540
rect 62956 2500 62996 2540
rect 63436 2500 63476 2540
rect 67468 2500 67508 2540
rect 73036 2500 73076 2540
rect 73420 2500 73460 2540
rect 73804 2500 73844 2540
rect 74188 2500 74228 2540
rect 74860 2500 74900 2540
rect 75724 2500 75764 2540
rect 77164 2500 77204 2540
rect 78700 2500 78740 2540
rect 81772 2500 81812 2540
rect 83308 2500 83348 2540
rect 84844 2500 84884 2540
rect 85228 2500 85268 2540
rect 85612 2500 85652 2540
rect 85996 2500 86036 2540
rect 86380 2500 86420 2540
rect 93004 2500 93044 2540
rect 93676 2500 93716 2540
rect 95212 2500 95252 2540
rect 96460 2500 96500 2540
rect 96844 2500 96884 2540
rect 97228 2500 97268 2540
rect 97612 2500 97652 2540
rect 97996 2500 98036 2540
rect 55084 2416 55124 2456
rect 55564 2416 55604 2456
rect 56140 2416 56180 2456
rect 58828 2416 58868 2456
rect 60556 2416 60596 2456
rect 61132 2416 61172 2456
rect 61612 2416 61652 2456
rect 61900 2416 61940 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 1516 1912 1556 1952
rect 1708 1912 1748 1952
rect 5356 1912 5396 1952
rect 5548 1912 5588 1952
rect 6796 1912 6836 1952
rect 6988 1912 7028 1952
rect 19372 1912 19412 1952
rect 19564 1912 19604 1952
rect 24652 1912 24692 1952
rect 24844 1912 24884 1952
rect 25900 1912 25940 1952
rect 26092 1912 26132 1952
rect 31948 1912 31988 1952
rect 32140 1912 32180 1952
rect 43660 1912 43700 1952
rect 43852 1912 43892 1952
rect 51244 1912 51284 1952
rect 51436 1912 51476 1952
rect 51820 1912 51860 1952
rect 52108 1912 52148 1952
rect 52300 1912 52340 1952
rect 52876 1912 52916 1952
rect 53164 1912 53204 1952
rect 53356 1912 53396 1952
rect 54316 1912 54356 1952
rect 54508 1912 54548 1952
rect 57004 1912 57044 1952
rect 57196 1912 57236 1952
rect 57484 1912 57524 1952
rect 57868 1912 57908 1952
rect 58060 1912 58100 1952
rect 58732 1912 58772 1952
rect 58924 1912 58964 1952
rect 59980 1912 60020 1952
rect 60172 1912 60212 1952
rect 62572 1912 62612 1952
rect 62764 1912 62804 1952
rect 64876 1912 64916 1952
rect 65068 1912 65108 1952
rect 66412 1912 66452 1952
rect 66604 1912 66644 1952
rect 67660 1912 67700 1952
rect 67852 1912 67892 1952
rect 79948 1912 79988 1952
rect 80140 1912 80180 1952
rect 80812 1912 80852 1952
rect 81004 1912 81044 1952
rect 92524 1912 92564 1952
rect 92716 1912 92756 1952
rect 97900 1912 97940 1952
rect 98092 1933 98132 1973
rect 25996 1828 26036 1868
rect 51340 1828 51380 1868
rect 60076 1828 60116 1868
rect 51820 1744 51860 1784
rect 52876 1744 52916 1784
rect 57484 1744 57524 1784
rect 1612 1660 1652 1700
rect 5452 1660 5492 1700
rect 6796 1660 6836 1700
rect 19468 1660 19508 1700
rect 24748 1660 24788 1700
rect 31948 1660 31988 1700
rect 43756 1660 43796 1700
rect 51628 1660 51668 1700
rect 52108 1660 52148 1700
rect 52684 1660 52724 1700
rect 53164 1660 53204 1700
rect 54508 1660 54548 1700
rect 57196 1660 57236 1700
rect 57676 1660 57716 1700
rect 57868 1660 57908 1700
rect 58732 1660 58772 1700
rect 62668 1660 62708 1700
rect 64972 1660 65012 1700
rect 66508 1660 66548 1700
rect 67756 1660 67796 1700
rect 80140 1660 80180 1700
rect 80908 1660 80948 1700
rect 92620 1660 92660 1700
rect 97996 1660 98036 1700
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 6988 1324 7028 1364
rect 14284 1324 14324 1364
rect 16588 1324 16628 1364
rect 20428 1324 20468 1364
rect 24652 1324 24692 1364
rect 30700 1324 30740 1364
rect 63052 1324 63092 1364
rect 66892 1324 66932 1364
rect 70732 1324 70772 1364
rect 72268 1324 72308 1364
rect 82828 1324 82868 1364
rect 85516 1324 85556 1364
rect 85900 1324 85940 1364
rect 98380 1324 98420 1364
rect 31660 1240 31700 1280
rect 50956 1240 50996 1280
rect 51436 1214 51476 1254
rect 52204 1240 52244 1280
rect 54124 1240 54164 1280
rect 54604 1240 54644 1280
rect 55084 1240 55124 1280
rect 56716 1240 56756 1280
rect 57196 1240 57236 1280
rect 57772 1240 57812 1280
rect 59308 1240 59348 1280
rect 59596 1240 59636 1280
rect 60172 1240 60212 1280
rect 60652 1240 60692 1280
rect 66604 1156 66644 1196
rect 1036 1072 1076 1112
rect 1228 1072 1268 1112
rect 1420 1072 1460 1112
rect 1612 1072 1652 1112
rect 1804 1072 1844 1112
rect 1996 1072 2036 1112
rect 2188 1072 2228 1112
rect 2380 1072 2420 1112
rect 2572 1072 2612 1112
rect 2764 1072 2804 1112
rect 2956 1072 2996 1112
rect 3148 1072 3188 1112
rect 3340 1072 3380 1112
rect 3532 1072 3572 1112
rect 3724 1072 3764 1112
rect 3916 1072 3956 1112
rect 4108 1085 4148 1125
rect 4300 1072 4340 1112
rect 4493 1085 4533 1125
rect 4684 1072 4724 1112
rect 4876 1072 4916 1112
rect 5068 1072 5108 1112
rect 5260 1072 5300 1112
rect 5452 1072 5492 1112
rect 5644 1072 5684 1112
rect 5836 1072 5876 1112
rect 6038 1061 6078 1101
rect 6217 1061 6257 1101
rect 6412 1072 6452 1112
rect 6604 1072 6644 1112
rect 6807 1061 6847 1101
rect 6995 1085 7035 1125
rect 7180 1072 7220 1112
rect 7372 1072 7412 1112
rect 7564 1072 7604 1112
rect 7756 1072 7796 1112
rect 7948 1072 7988 1112
rect 8140 1072 8180 1112
rect 8332 1072 8372 1112
rect 8524 1072 8564 1112
rect 8716 1072 8756 1112
rect 8908 1072 8948 1112
rect 9100 1072 9140 1112
rect 9292 1072 9332 1112
rect 9484 1072 9524 1112
rect 9676 1072 9716 1112
rect 9868 1072 9908 1112
rect 10060 1072 10100 1112
rect 10252 1072 10292 1112
rect 10444 1072 10484 1112
rect 10636 1072 10676 1112
rect 10828 1072 10868 1112
rect 11020 1072 11060 1112
rect 11212 1072 11252 1112
rect 11404 1072 11444 1112
rect 11596 1085 11636 1125
rect 11788 1072 11828 1112
rect 11980 1072 12020 1112
rect 12172 1072 12212 1112
rect 12364 1072 12404 1112
rect 12556 1072 12596 1112
rect 12748 1069 12788 1109
rect 12940 1072 12980 1112
rect 13132 1072 13172 1112
rect 13324 1072 13364 1112
rect 13516 1072 13556 1112
rect 13708 1072 13748 1112
rect 13900 1072 13940 1112
rect 14092 1072 14132 1112
rect 14284 1072 14324 1112
rect 14476 1072 14516 1112
rect 14668 1072 14708 1112
rect 14860 1072 14900 1112
rect 15052 1072 15092 1112
rect 15244 1072 15284 1112
rect 15436 1072 15476 1112
rect 15628 1072 15668 1112
rect 15820 1072 15860 1112
rect 16012 1072 16052 1112
rect 16204 1072 16244 1112
rect 16396 1072 16436 1112
rect 16588 1085 16628 1125
rect 16780 1085 16820 1125
rect 16972 1072 17012 1112
rect 17164 1072 17204 1112
rect 17356 1072 17396 1112
rect 17548 1072 17588 1112
rect 17740 1072 17780 1112
rect 17932 1072 17972 1112
rect 18114 1069 18154 1109
rect 18316 1072 18356 1112
rect 18508 1072 18548 1112
rect 18700 1072 18740 1112
rect 18892 1072 18932 1112
rect 19084 1072 19124 1112
rect 19276 1085 19316 1125
rect 19468 1072 19508 1112
rect 19660 1072 19700 1112
rect 19852 1072 19892 1112
rect 20044 1072 20084 1112
rect 20236 1072 20276 1112
rect 20428 1072 20468 1112
rect 20620 1061 20660 1101
rect 20812 1072 20852 1112
rect 21004 1072 21044 1112
rect 21196 1072 21236 1112
rect 21388 1072 21428 1112
rect 21580 1085 21620 1125
rect 21772 1072 21812 1112
rect 21964 1072 22004 1112
rect 22156 1072 22196 1112
rect 22348 1072 22388 1112
rect 22540 1072 22580 1112
rect 22732 1072 22772 1112
rect 22924 1072 22964 1112
rect 23116 1072 23156 1112
rect 23308 1072 23348 1112
rect 23500 1072 23540 1112
rect 23692 1072 23732 1112
rect 23884 1072 23924 1112
rect 24076 1072 24116 1112
rect 24268 1072 24308 1112
rect 24460 1072 24500 1112
rect 24652 1072 24692 1112
rect 24844 1072 24884 1112
rect 25036 1072 25076 1112
rect 25516 1072 25556 1112
rect 25708 1072 25748 1112
rect 25900 1072 25940 1112
rect 26092 1072 26132 1112
rect 26284 1072 26324 1112
rect 26476 1072 26516 1112
rect 26668 1072 26708 1112
rect 26860 1072 26900 1112
rect 27052 1072 27092 1112
rect 27244 1072 27284 1112
rect 27436 1072 27476 1112
rect 27628 1072 27668 1112
rect 27820 1072 27860 1112
rect 28012 1072 28052 1112
rect 28204 1072 28244 1112
rect 28396 1072 28436 1112
rect 28588 1072 28628 1112
rect 28780 1072 28820 1112
rect 28972 1072 29012 1112
rect 29164 1072 29204 1112
rect 29356 1072 29396 1112
rect 29548 1072 29588 1112
rect 29740 1072 29780 1112
rect 29932 1072 29972 1112
rect 30124 1072 30164 1112
rect 30316 1072 30356 1112
rect 30508 1072 30548 1112
rect 30700 1072 30740 1112
rect 30892 1072 30932 1112
rect 31084 1072 31124 1112
rect 31468 1072 31508 1112
rect 31660 1072 31700 1112
rect 31852 1072 31892 1112
rect 32044 1072 32084 1112
rect 32236 1085 32276 1125
rect 32428 1072 32468 1112
rect 32620 1072 32660 1112
rect 32812 1072 32852 1112
rect 33004 1061 33044 1101
rect 33196 1072 33236 1112
rect 33388 1072 33428 1112
rect 33580 1072 33620 1112
rect 33772 1072 33812 1112
rect 33964 1072 34004 1112
rect 34156 1085 34196 1125
rect 34348 1072 34388 1112
rect 34540 1072 34580 1112
rect 34732 1072 34772 1112
rect 34924 1072 34964 1112
rect 35116 1085 35156 1125
rect 35308 1072 35348 1112
rect 35500 1072 35540 1112
rect 35692 1072 35732 1112
rect 35884 1072 35924 1112
rect 36076 1072 36116 1112
rect 36268 1072 36308 1112
rect 36460 1072 36500 1112
rect 36652 1072 36692 1112
rect 36844 1072 36884 1112
rect 37036 1072 37076 1112
rect 37324 1072 37364 1112
rect 37516 1072 37556 1112
rect 37708 1072 37748 1112
rect 37900 1072 37940 1112
rect 38092 1072 38132 1112
rect 38284 1072 38324 1112
rect 38476 1072 38516 1112
rect 38668 1072 38708 1112
rect 38860 1072 38900 1112
rect 39052 1072 39092 1112
rect 39244 1072 39284 1112
rect 39436 1072 39476 1112
rect 39628 1072 39668 1112
rect 39820 1072 39860 1112
rect 40012 1072 40052 1112
rect 40204 1072 40244 1112
rect 40396 1072 40436 1112
rect 40588 1072 40628 1112
rect 40780 1072 40820 1112
rect 40972 1072 41012 1112
rect 41164 1072 41204 1112
rect 41356 1072 41396 1112
rect 41548 1072 41588 1112
rect 41740 1072 41780 1112
rect 41943 1061 41983 1101
rect 42124 1072 42164 1112
rect 42316 1072 42356 1112
rect 42508 1072 42548 1112
rect 42700 1072 42740 1112
rect 42892 1072 42932 1112
rect 43084 1072 43124 1112
rect 43276 1072 43316 1112
rect 43564 1072 43604 1112
rect 43756 1072 43796 1112
rect 43948 1072 43988 1112
rect 44140 1072 44180 1112
rect 44343 1085 44383 1125
rect 44524 1072 44564 1112
rect 44716 1072 44756 1112
rect 44908 1072 44948 1112
rect 45100 1072 45140 1112
rect 45292 1072 45332 1112
rect 45484 1072 45524 1112
rect 45676 1072 45716 1112
rect 45868 1072 45908 1112
rect 46060 1072 46100 1112
rect 46252 1072 46292 1112
rect 46444 1072 46484 1112
rect 46636 1072 46676 1112
rect 46828 1072 46868 1112
rect 47020 1072 47060 1112
rect 47212 1072 47252 1112
rect 47404 1072 47444 1112
rect 47596 1072 47636 1112
rect 47788 1072 47828 1112
rect 47980 1072 48020 1112
rect 48172 1072 48212 1112
rect 48364 1072 48404 1112
rect 48556 1072 48596 1112
rect 48748 1072 48788 1112
rect 48940 1072 48980 1112
rect 49132 1072 49172 1112
rect 49324 1072 49364 1112
rect 49516 1072 49556 1112
rect 50380 1072 50420 1112
rect 50572 1072 50612 1112
rect 50956 1072 50996 1112
rect 51436 1072 51476 1112
rect 52204 1072 52244 1112
rect 52492 1072 52532 1112
rect 52684 1072 52724 1112
rect 53548 1072 53588 1112
rect 53740 1072 53780 1112
rect 54124 1072 54164 1112
rect 54604 1084 54644 1124
rect 55084 1072 55124 1112
rect 55372 1072 55412 1112
rect 55564 1072 55604 1112
rect 56236 1072 56276 1112
rect 56428 1072 56468 1112
rect 56716 1075 56756 1115
rect 57196 1072 57236 1112
rect 57772 1072 57812 1112
rect 58156 1072 58196 1112
rect 58348 1072 58388 1112
rect 59116 1072 59156 1112
rect 59308 1072 59348 1112
rect 59596 1072 59636 1112
rect 60172 1072 60212 1112
rect 60652 1072 60692 1112
rect 60940 1072 60980 1112
rect 61132 1072 61172 1112
rect 62668 1072 62708 1112
rect 62860 1061 62900 1101
rect 63052 1072 63092 1112
rect 63244 1072 63284 1112
rect 63436 1072 63476 1112
rect 63628 1072 63668 1112
rect 63820 1085 63860 1125
rect 64012 1072 64052 1112
rect 64204 1072 64244 1112
rect 64396 1072 64436 1112
rect 64588 1072 64628 1112
rect 64780 1072 64820 1112
rect 64972 1072 65012 1112
rect 65164 1072 65204 1112
rect 65356 1072 65396 1112
rect 65548 1072 65588 1112
rect 65740 1072 65780 1112
rect 65932 1072 65972 1112
rect 66124 1072 66164 1112
rect 66316 1072 66356 1112
rect 66508 1072 66548 1112
rect 66700 1072 66740 1112
rect 66885 1085 66925 1125
rect 67084 1072 67124 1112
rect 67276 1072 67316 1112
rect 67468 1072 67508 1112
rect 67660 1072 67700 1112
rect 67852 1072 67892 1112
rect 68044 1072 68084 1112
rect 68236 1072 68276 1112
rect 68428 1072 68468 1112
rect 68620 1072 68660 1112
rect 68812 1072 68852 1112
rect 69004 1072 69044 1112
rect 69196 1072 69236 1112
rect 69388 1072 69428 1112
rect 69590 1069 69630 1109
rect 69772 1072 69812 1112
rect 69964 1072 70004 1112
rect 70156 1072 70196 1112
rect 70348 1072 70388 1112
rect 70521 1077 70561 1117
rect 70732 1072 70772 1112
rect 70924 1072 70964 1112
rect 71116 1072 71156 1112
rect 71308 1072 71348 1112
rect 71500 1072 71540 1112
rect 71692 1072 71732 1112
rect 71884 1072 71924 1112
rect 72076 1072 72116 1112
rect 72268 1072 72308 1112
rect 72460 1072 72500 1112
rect 72652 1072 72692 1112
rect 72844 1072 72884 1112
rect 73036 1072 73076 1112
rect 73228 1072 73268 1112
rect 73420 1072 73460 1112
rect 73612 1072 73652 1112
rect 73804 1072 73844 1112
rect 73996 1072 74036 1112
rect 74188 1072 74228 1112
rect 74380 1072 74420 1112
rect 74572 1072 74612 1112
rect 74764 1072 74804 1112
rect 74956 1072 74996 1112
rect 75148 1072 75188 1112
rect 75340 1073 75380 1113
rect 75532 1072 75572 1112
rect 75724 1072 75764 1112
rect 75916 1072 75956 1112
rect 76108 1072 76148 1112
rect 76300 1072 76340 1112
rect 76492 1061 76532 1101
rect 76684 1072 76724 1112
rect 76876 1072 76916 1112
rect 77068 1072 77108 1112
rect 77260 1072 77300 1112
rect 77452 1072 77492 1112
rect 77644 1072 77684 1112
rect 77836 1072 77876 1112
rect 78028 1072 78068 1112
rect 78220 1072 78260 1112
rect 78412 1072 78452 1112
rect 78604 1072 78644 1112
rect 78796 1072 78836 1112
rect 78988 1072 79028 1112
rect 79180 1072 79220 1112
rect 79372 1072 79412 1112
rect 79564 1072 79604 1112
rect 79756 1072 79796 1112
rect 79948 1072 79988 1112
rect 80140 1072 80180 1112
rect 80332 1072 80372 1112
rect 80524 1072 80564 1112
rect 80908 1072 80948 1112
rect 81100 1072 81140 1112
rect 81292 1072 81332 1112
rect 81484 1072 81524 1112
rect 81676 1072 81716 1112
rect 81868 1072 81908 1112
rect 82060 1072 82100 1112
rect 82252 1072 82292 1112
rect 82444 1072 82484 1112
rect 82636 1072 82676 1112
rect 82828 1072 82868 1112
rect 83020 1072 83060 1112
rect 83212 1072 83252 1112
rect 83393 1069 83433 1109
rect 83596 1072 83636 1112
rect 83793 1069 83833 1109
rect 83980 1072 84020 1112
rect 84172 1072 84212 1112
rect 84364 1072 84404 1112
rect 84556 1072 84596 1112
rect 84748 1072 84788 1112
rect 84940 1072 84980 1112
rect 85132 1072 85172 1112
rect 85324 1072 85364 1112
rect 85516 1072 85556 1112
rect 85708 1072 85748 1112
rect 85900 1085 85940 1125
rect 86092 1072 86132 1112
rect 86284 1072 86324 1112
rect 86476 1072 86516 1112
rect 86668 1072 86708 1112
rect 86860 1072 86900 1112
rect 87052 1072 87092 1112
rect 87244 1072 87284 1112
rect 87436 1072 87476 1112
rect 87628 1072 87668 1112
rect 87820 1072 87860 1112
rect 88012 1072 88052 1112
rect 88204 1072 88244 1112
rect 88396 1085 88436 1125
rect 88588 1072 88628 1112
rect 88780 1072 88820 1112
rect 88972 1072 89012 1112
rect 89164 1072 89204 1112
rect 89356 1072 89396 1112
rect 89548 1072 89588 1112
rect 89740 1072 89780 1112
rect 89932 1072 89972 1112
rect 90124 1072 90164 1112
rect 90316 1072 90356 1112
rect 90508 1072 90548 1112
rect 90700 1061 90740 1101
rect 90892 1072 90932 1112
rect 91084 1072 91124 1112
rect 91276 1072 91316 1112
rect 91468 1072 91508 1112
rect 91660 1072 91700 1112
rect 91852 1072 91892 1112
rect 92044 1072 92084 1112
rect 92236 1072 92276 1112
rect 92428 1072 92468 1112
rect 92620 1072 92660 1112
rect 92812 1072 92852 1112
rect 93004 1072 93044 1112
rect 93196 1072 93236 1112
rect 93388 1072 93428 1112
rect 93580 1072 93620 1112
rect 93772 1072 93812 1112
rect 93964 1072 94004 1112
rect 94156 1072 94196 1112
rect 94348 1072 94388 1112
rect 94540 1061 94580 1101
rect 94732 1069 94772 1109
rect 94924 1061 94964 1101
rect 95116 1061 95156 1101
rect 95308 1061 95348 1101
rect 95500 1072 95540 1112
rect 95699 1069 95739 1109
rect 95884 1072 95924 1112
rect 96076 1072 96116 1112
rect 96268 1072 96308 1112
rect 96460 1072 96500 1112
rect 96652 1072 96692 1112
rect 96844 1072 96884 1112
rect 97036 1072 97076 1112
rect 97227 1085 97267 1125
rect 97420 1072 97460 1112
rect 97612 1072 97652 1112
rect 97804 1072 97844 1112
rect 97995 1085 98035 1125
rect 98188 1072 98228 1112
rect 98380 1072 98420 1112
rect 98572 1072 98612 1112
rect 98764 1072 98804 1112
rect 98956 1072 98996 1112
rect 99148 1072 99188 1112
rect 5356 988 5396 1028
rect 35020 988 35060 1028
rect 67756 988 67796 1028
rect 89068 988 89108 1028
rect 91372 988 91412 1028
rect 92140 988 92180 1028
rect 97900 988 97940 1028
rect 1132 904 1172 944
rect 1516 904 1556 944
rect 1900 904 1940 944
rect 2284 904 2324 944
rect 2668 904 2708 944
rect 3052 904 3092 944
rect 3436 904 3476 944
rect 3820 904 3860 944
rect 4204 904 4244 944
rect 4588 904 4628 944
rect 4972 904 5012 944
rect 5740 904 5780 944
rect 6124 904 6164 944
rect 6508 904 6548 944
rect 7276 904 7316 944
rect 7660 904 7700 944
rect 8044 904 8084 944
rect 8428 904 8468 944
rect 8812 904 8852 944
rect 9196 904 9236 944
rect 9580 904 9620 944
rect 9964 904 10004 944
rect 10348 904 10388 944
rect 10732 904 10772 944
rect 11116 904 11156 944
rect 11500 904 11540 944
rect 11884 904 11924 944
rect 12268 904 12308 944
rect 12652 904 12692 944
rect 13036 904 13076 944
rect 13420 904 13460 944
rect 13804 904 13844 944
rect 14572 904 14612 944
rect 14956 904 14996 944
rect 15340 904 15380 944
rect 15724 904 15764 944
rect 16108 904 16148 944
rect 16876 904 16916 944
rect 17260 904 17300 944
rect 17644 904 17684 944
rect 18028 904 18068 944
rect 18412 904 18452 944
rect 18796 904 18836 944
rect 19180 904 19220 944
rect 19564 904 19604 944
rect 19948 904 19988 944
rect 20716 904 20756 944
rect 21100 904 21140 944
rect 21484 904 21524 944
rect 21868 904 21908 944
rect 22252 904 22292 944
rect 22636 904 22676 944
rect 23020 904 23060 944
rect 23404 904 23444 944
rect 23788 904 23828 944
rect 24172 904 24212 944
rect 24940 904 24980 944
rect 25612 904 25652 944
rect 25996 904 26036 944
rect 26380 904 26420 944
rect 26764 904 26804 944
rect 27148 904 27188 944
rect 27532 904 27572 944
rect 27916 904 27956 944
rect 28300 904 28340 944
rect 28684 904 28724 944
rect 29068 904 29108 944
rect 29452 904 29492 944
rect 29836 904 29876 944
rect 30220 904 30260 944
rect 30988 904 31028 944
rect 31948 904 31988 944
rect 32332 904 32372 944
rect 32716 904 32756 944
rect 33100 904 33140 944
rect 33484 904 33524 944
rect 33868 904 33908 944
rect 34252 904 34292 944
rect 34636 904 34676 944
rect 35404 904 35444 944
rect 35788 904 35828 944
rect 36172 904 36212 944
rect 36556 904 36596 944
rect 36940 904 36980 944
rect 37420 904 37460 944
rect 37804 904 37844 944
rect 38188 904 38228 944
rect 38572 904 38612 944
rect 38956 904 38996 944
rect 39340 904 39380 944
rect 39724 904 39764 944
rect 40108 904 40148 944
rect 40492 904 40532 944
rect 40876 904 40916 944
rect 41260 904 41300 944
rect 41644 904 41684 944
rect 42028 904 42068 944
rect 42412 904 42452 944
rect 42796 904 42836 944
rect 43180 904 43220 944
rect 43660 904 43700 944
rect 44044 904 44084 944
rect 44428 904 44468 944
rect 44812 904 44852 944
rect 45196 904 45236 944
rect 45580 904 45620 944
rect 45964 904 46004 944
rect 46348 904 46388 944
rect 46732 904 46772 944
rect 47116 904 47156 944
rect 47500 904 47540 944
rect 47884 904 47924 944
rect 48268 904 48308 944
rect 48652 904 48692 944
rect 49036 904 49076 944
rect 49420 904 49460 944
rect 50476 904 50516 944
rect 50764 904 50804 944
rect 51244 904 51284 944
rect 52012 904 52052 944
rect 52588 904 52628 944
rect 53644 904 53684 944
rect 53932 904 53972 944
rect 54412 904 54452 944
rect 54892 904 54932 944
rect 55468 904 55508 944
rect 56332 904 56372 944
rect 56908 904 56948 944
rect 57388 904 57428 944
rect 57964 904 58004 944
rect 58252 904 58292 944
rect 59788 904 59828 944
rect 59980 904 60020 944
rect 60460 904 60500 944
rect 61036 904 61076 944
rect 62764 904 62804 944
rect 63532 904 63572 944
rect 63916 904 63956 944
rect 64300 904 64340 944
rect 64684 904 64724 944
rect 65068 904 65108 944
rect 65452 904 65492 944
rect 65836 904 65876 944
rect 66220 904 66260 944
rect 67372 904 67412 944
rect 68140 904 68180 944
rect 68524 904 68564 944
rect 68908 904 68948 944
rect 69292 904 69332 944
rect 69676 904 69716 944
rect 70060 904 70100 944
rect 70444 904 70484 944
rect 71212 904 71252 944
rect 71596 904 71636 944
rect 71980 904 72020 944
rect 72748 904 72788 944
rect 73132 904 73172 944
rect 73516 904 73556 944
rect 73900 904 73940 944
rect 74284 904 74324 944
rect 74668 904 74708 944
rect 75052 904 75092 944
rect 75436 904 75476 944
rect 75820 904 75860 944
rect 76204 904 76244 944
rect 76588 904 76628 944
rect 76972 904 77012 944
rect 77356 904 77396 944
rect 77740 904 77780 944
rect 78124 904 78164 944
rect 78508 904 78548 944
rect 78892 904 78932 944
rect 79276 904 79316 944
rect 79660 904 79700 944
rect 80044 904 80084 944
rect 80428 904 80468 944
rect 81004 904 81044 944
rect 81388 904 81428 944
rect 81772 904 81812 944
rect 82156 904 82196 944
rect 82540 904 82580 944
rect 83308 904 83348 944
rect 83692 904 83732 944
rect 84076 904 84116 944
rect 84460 904 84500 944
rect 84844 904 84884 944
rect 85228 904 85268 944
rect 86380 904 86420 944
rect 86764 904 86804 944
rect 87148 904 87188 944
rect 87532 904 87572 944
rect 87916 904 87956 944
rect 88300 904 88340 944
rect 88684 904 88724 944
rect 89452 904 89492 944
rect 89836 904 89876 944
rect 90220 904 90260 944
rect 90604 904 90644 944
rect 90988 904 91028 944
rect 91756 904 91796 944
rect 92524 904 92564 944
rect 92908 904 92948 944
rect 93292 904 93332 944
rect 93676 904 93716 944
rect 94060 904 94100 944
rect 94444 904 94484 944
rect 94828 904 94868 944
rect 95212 904 95252 944
rect 95596 904 95636 944
rect 95980 904 96020 944
rect 96364 904 96404 944
rect 96748 904 96788 944
rect 97132 904 97172 944
rect 97516 904 97556 944
rect 98668 904 98708 944
rect 99052 904 99092 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 6200 9920 6280 10000
rect 17144 9920 17224 10000
rect 28088 9920 28168 10000
rect 39032 9920 39112 10000
rect 49420 9940 49844 9980
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 6220 7001 6260 9920
rect 6219 6992 6261 7001
rect 6219 6952 6220 6992
rect 6260 6952 6261 6992
rect 6219 6943 6261 6952
rect 17164 6917 17204 9920
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 28108 7001 28148 9920
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 24555 6992 24597 7001
rect 24555 6952 24556 6992
rect 24596 6952 24597 6992
rect 24555 6943 24597 6952
rect 28107 6992 28149 7001
rect 28107 6952 28108 6992
rect 28148 6952 28149 6992
rect 28107 6943 28149 6952
rect 17163 6908 17205 6917
rect 17163 6868 17164 6908
rect 17204 6868 17205 6908
rect 17163 6859 17205 6868
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 24556 5657 24596 6943
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 39052 6665 39092 9920
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 41067 6992 41109 7001
rect 41067 6952 41068 6992
rect 41108 6952 41109 6992
rect 41067 6943 41109 6952
rect 41739 6992 41781 7001
rect 41739 6952 41740 6992
rect 41780 6952 41781 6992
rect 41739 6943 41781 6952
rect 39051 6656 39093 6665
rect 39051 6616 39052 6656
rect 39092 6616 39093 6656
rect 39051 6607 39093 6616
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 24555 5648 24597 5657
rect 24555 5608 24556 5648
rect 24596 5608 24597 5648
rect 24555 5599 24597 5608
rect 41068 5648 41108 6943
rect 41355 6908 41397 6917
rect 41355 6868 41356 6908
rect 41396 6868 41397 6908
rect 41355 6859 41397 6868
rect 41068 5599 41108 5608
rect 41356 5648 41396 6859
rect 41740 6581 41780 6943
rect 42027 6908 42069 6917
rect 42027 6868 42028 6908
rect 42068 6868 42069 6908
rect 42027 6859 42069 6868
rect 41739 6572 41781 6581
rect 41739 6532 41740 6572
rect 41780 6532 41781 6572
rect 41739 6523 41781 6532
rect 41740 6488 41780 6523
rect 42028 6497 42068 6859
rect 45772 6656 45812 6667
rect 44524 6497 44564 6582
rect 45772 6581 45812 6616
rect 46731 6656 46773 6665
rect 46731 6616 46732 6656
rect 46772 6616 46773 6656
rect 46731 6607 46773 6616
rect 47595 6656 47637 6665
rect 47595 6616 47596 6656
rect 47636 6616 47637 6656
rect 47595 6607 47637 6616
rect 48459 6656 48501 6665
rect 48459 6616 48460 6656
rect 48500 6616 48501 6656
rect 48459 6607 48501 6616
rect 48556 6656 48596 6665
rect 44715 6572 44757 6581
rect 44715 6532 44716 6572
rect 44756 6532 44757 6572
rect 44715 6523 44757 6532
rect 45771 6572 45813 6581
rect 45771 6532 45772 6572
rect 45812 6532 45813 6572
rect 45771 6523 45813 6532
rect 46347 6572 46389 6581
rect 46539 6572 46581 6581
rect 46347 6532 46348 6572
rect 46388 6532 46484 6572
rect 46347 6523 46389 6532
rect 41740 6438 41780 6448
rect 42027 6488 42069 6497
rect 42027 6448 42028 6488
rect 42068 6448 42069 6488
rect 42027 6439 42069 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44716 6488 44756 6523
rect 42028 6354 42068 6439
rect 44716 6437 44756 6448
rect 45867 6488 45909 6497
rect 45867 6448 45868 6488
rect 45908 6448 45909 6488
rect 45867 6439 45909 6448
rect 46444 6488 46484 6532
rect 46539 6532 46540 6572
rect 46580 6532 46581 6572
rect 46539 6523 46581 6532
rect 46444 6439 46484 6448
rect 46540 6488 46580 6523
rect 45868 6354 45908 6439
rect 46540 6437 46580 6448
rect 46635 6488 46677 6497
rect 46635 6448 46636 6488
rect 46676 6448 46677 6488
rect 46635 6439 46677 6448
rect 46636 6404 46676 6439
rect 46636 6353 46676 6364
rect 41740 6320 41780 6329
rect 41644 6280 41740 6320
rect 41356 5599 41396 5608
rect 41451 5648 41493 5657
rect 41451 5608 41452 5648
rect 41492 5608 41493 5648
rect 41451 5599 41493 5608
rect 41452 5489 41492 5599
rect 41548 5564 41588 5573
rect 41260 5480 41300 5489
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 22444 4976 22484 4985
rect 22348 4724 22388 4733
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 18891 4556 18933 4565
rect 18891 4516 18892 4556
rect 18932 4516 18933 4556
rect 18891 4507 18933 4516
rect 19467 4556 19509 4565
rect 19467 4516 19468 4556
rect 19508 4516 19509 4556
rect 19467 4507 19509 4516
rect 20043 4556 20085 4565
rect 20043 4516 20044 4556
rect 20084 4516 20085 4556
rect 20043 4507 20085 4516
rect 7564 4313 7604 4398
rect 18507 4388 18549 4397
rect 18507 4348 18508 4388
rect 18548 4348 18549 4388
rect 18507 4339 18549 4348
rect 6987 4304 7029 4313
rect 6987 4264 6988 4304
rect 7028 4264 7029 4304
rect 6987 4255 7029 4264
rect 7563 4304 7605 4313
rect 7563 4264 7564 4304
rect 7604 4264 7605 4304
rect 7563 4255 7605 4264
rect 6988 4136 7028 4255
rect 6988 4087 7028 4096
rect 7179 4136 7221 4145
rect 7179 4096 7180 4136
rect 7220 4096 7221 4136
rect 7179 4087 7221 4096
rect 7563 4136 7605 4145
rect 7563 4096 7564 4136
rect 7604 4096 7605 4136
rect 7563 4087 7605 4096
rect 18315 4136 18357 4145
rect 18315 4096 18316 4136
rect 18356 4096 18357 4136
rect 18315 4087 18357 4096
rect 18412 4136 18452 4145
rect 18508 4136 18548 4339
rect 18452 4096 18548 4136
rect 18412 4087 18452 4096
rect 7180 4002 7220 4087
rect 7564 4002 7604 4087
rect 18124 4052 18164 4061
rect 7084 3968 7124 3977
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4395 3632 4437 3641
rect 4395 3592 4396 3632
rect 4436 3592 4437 3632
rect 7084 3632 7124 3928
rect 7372 3968 7412 3977
rect 7084 3592 7220 3632
rect 4395 3583 4437 3592
rect 1900 3464 1940 3473
rect 1804 3424 1900 3464
rect 1611 3128 1653 3137
rect 1611 3088 1612 3128
rect 1652 3088 1653 3128
rect 1611 3079 1653 3088
rect 1612 2624 1652 3079
rect 1612 2575 1652 2584
rect 1804 2624 1844 3424
rect 1900 3415 1940 3424
rect 2091 3464 2133 3473
rect 2091 3424 2092 3464
rect 2132 3424 2133 3464
rect 2091 3415 2133 3424
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 4203 3464 4245 3473
rect 4203 3424 4204 3464
rect 4244 3424 4245 3464
rect 4203 3415 4245 3424
rect 4396 3464 4436 3583
rect 6411 3548 6453 3557
rect 6411 3508 6412 3548
rect 6452 3508 6453 3548
rect 6411 3499 6453 3508
rect 4396 3415 4436 3424
rect 4587 3464 4629 3473
rect 4587 3424 4588 3464
rect 4628 3424 4629 3464
rect 4587 3415 4629 3424
rect 4780 3464 4820 3473
rect 4971 3464 5013 3473
rect 4820 3424 4916 3464
rect 4780 3415 4820 3424
rect 2092 3330 2132 3415
rect 2667 3296 2709 3305
rect 2667 3256 2668 3296
rect 2708 3256 2709 3296
rect 2667 3247 2709 3256
rect 1996 3212 2036 3221
rect 1708 2540 1748 2549
rect 1708 2120 1748 2500
rect 1804 2465 1844 2584
rect 1900 3172 1996 3212
rect 1803 2456 1845 2465
rect 1803 2416 1804 2456
rect 1844 2416 1845 2456
rect 1803 2407 1845 2416
rect 1324 2080 1748 2120
rect 1035 1280 1077 1289
rect 1035 1240 1036 1280
rect 1076 1240 1077 1280
rect 1035 1231 1077 1240
rect 843 1196 885 1205
rect 843 1156 844 1196
rect 884 1156 885 1196
rect 843 1147 885 1156
rect 844 80 884 1147
rect 1036 1112 1076 1231
rect 1228 1121 1268 1206
rect 1036 1063 1076 1072
rect 1227 1112 1269 1121
rect 1227 1072 1228 1112
rect 1268 1072 1269 1112
rect 1227 1063 1269 1072
rect 1132 944 1172 953
rect 1324 944 1364 2080
rect 1515 1952 1557 1961
rect 1515 1912 1516 1952
rect 1556 1912 1557 1952
rect 1515 1903 1557 1912
rect 1708 1952 1748 1961
rect 1804 1952 1844 2407
rect 1748 1912 1844 1952
rect 1708 1903 1748 1912
rect 1516 1818 1556 1903
rect 1612 1700 1652 1709
rect 1516 1660 1612 1700
rect 1419 1280 1461 1289
rect 1419 1240 1420 1280
rect 1460 1240 1461 1280
rect 1419 1231 1461 1240
rect 1420 1112 1460 1231
rect 1516 1205 1556 1660
rect 1612 1651 1652 1660
rect 1900 1448 1940 3172
rect 1996 3163 2036 3172
rect 2092 2624 2132 2635
rect 2092 2465 2132 2584
rect 2283 2624 2325 2633
rect 2283 2584 2284 2624
rect 2324 2584 2325 2624
rect 2283 2575 2325 2584
rect 2476 2624 2516 2635
rect 2188 2540 2228 2549
rect 2091 2456 2133 2465
rect 2091 2416 2092 2456
rect 2132 2416 2133 2456
rect 2091 2407 2133 2416
rect 2188 1448 2228 2500
rect 2284 2490 2324 2575
rect 2476 2465 2516 2584
rect 2668 2624 2708 3247
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 3147 2792 3189 2801
rect 3147 2752 3148 2792
rect 3188 2752 3189 2792
rect 3147 2743 3189 2752
rect 2668 2575 2708 2584
rect 2956 2624 2996 2635
rect 2572 2540 2612 2549
rect 2475 2456 2517 2465
rect 2475 2416 2476 2456
rect 2516 2416 2517 2456
rect 2475 2407 2517 2416
rect 1708 1408 1940 1448
rect 2092 1408 2228 1448
rect 1515 1196 1557 1205
rect 1515 1156 1516 1196
rect 1556 1156 1557 1196
rect 1515 1147 1557 1156
rect 1612 1121 1652 1206
rect 1420 1063 1460 1072
rect 1611 1112 1653 1121
rect 1611 1072 1612 1112
rect 1652 1072 1653 1112
rect 1611 1063 1653 1072
rect 1516 944 1556 953
rect 1708 944 1748 1408
rect 1803 1196 1845 1205
rect 1803 1156 1804 1196
rect 1844 1156 1845 1196
rect 1803 1147 1845 1156
rect 1804 1112 1844 1147
rect 1804 1061 1844 1072
rect 1995 1112 2037 1121
rect 1995 1072 1996 1112
rect 2036 1072 2037 1112
rect 1995 1063 2037 1072
rect 1996 978 2036 1063
rect 1900 944 1940 953
rect 1036 904 1132 944
rect 1036 80 1076 904
rect 1132 895 1172 904
rect 1228 904 1364 944
rect 1420 904 1516 944
rect 1228 80 1268 904
rect 1420 80 1460 904
rect 1516 895 1556 904
rect 1612 904 1748 944
rect 1804 904 1900 944
rect 1612 80 1652 904
rect 1804 80 1844 904
rect 1900 895 1940 904
rect 2092 860 2132 1408
rect 2572 1364 2612 2500
rect 2859 2540 2901 2549
rect 2956 2540 2996 2584
rect 3148 2624 3188 2743
rect 3148 2575 3188 2584
rect 3340 2624 3380 2635
rect 2859 2500 2860 2540
rect 2900 2500 2996 2540
rect 3052 2540 3092 2549
rect 2859 2491 2901 2500
rect 3052 1700 3092 2500
rect 3243 2540 3285 2549
rect 3340 2540 3380 2584
rect 3531 2624 3573 2633
rect 3531 2584 3532 2624
rect 3572 2584 3573 2624
rect 3531 2575 3573 2584
rect 3724 2624 3764 3415
rect 4204 3330 4244 3415
rect 4588 3330 4628 3415
rect 4876 3221 4916 3424
rect 4971 3424 4972 3464
rect 5012 3424 5013 3464
rect 4971 3415 5013 3424
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 5740 3464 5780 3473
rect 4300 3212 4340 3221
rect 4204 3172 4300 3212
rect 3243 2500 3244 2540
rect 3284 2500 3380 2540
rect 3436 2540 3476 2549
rect 3243 2491 3285 2500
rect 2476 1324 2612 1364
rect 2860 1660 3092 1700
rect 3436 1700 3476 2500
rect 3532 2490 3572 2575
rect 3627 2540 3669 2549
rect 3724 2540 3764 2584
rect 3915 2624 3957 2633
rect 3915 2584 3916 2624
rect 3956 2584 3957 2624
rect 3915 2575 3957 2584
rect 3627 2500 3628 2540
rect 3668 2500 3764 2540
rect 3820 2540 3860 2549
rect 3627 2491 3669 2500
rect 3820 1952 3860 2500
rect 3916 2490 3956 2575
rect 4204 2540 4244 3172
rect 4300 3163 4340 3172
rect 4683 3212 4725 3221
rect 4683 3172 4684 3212
rect 4724 3172 4725 3212
rect 4683 3163 4725 3172
rect 4875 3212 4917 3221
rect 4875 3172 4876 3212
rect 4916 3172 4917 3212
rect 4875 3163 4917 3172
rect 4684 3078 4724 3163
rect 4972 3053 5012 3415
rect 5164 3330 5204 3415
rect 5068 3212 5108 3221
rect 4971 3044 5013 3053
rect 4971 3004 4972 3044
rect 5012 3004 5013 3044
rect 4971 2995 5013 3004
rect 4012 2500 4244 2540
rect 3628 1912 3860 1952
rect 3436 1660 3572 1700
rect 2188 1121 2228 1206
rect 2187 1112 2229 1121
rect 2187 1072 2188 1112
rect 2228 1072 2229 1112
rect 2187 1063 2229 1072
rect 2380 1112 2420 1121
rect 2284 944 2324 953
rect 1996 820 2132 860
rect 2188 904 2284 944
rect 1996 80 2036 820
rect 2188 80 2228 904
rect 2284 895 2324 904
rect 2380 701 2420 1072
rect 2379 692 2421 701
rect 2379 652 2380 692
rect 2420 652 2421 692
rect 2379 643 2421 652
rect 2476 524 2516 1324
rect 2571 1196 2613 1205
rect 2571 1156 2572 1196
rect 2612 1156 2613 1196
rect 2571 1147 2613 1156
rect 2572 1112 2612 1147
rect 2764 1121 2804 1206
rect 2572 1061 2612 1072
rect 2763 1112 2805 1121
rect 2763 1072 2764 1112
rect 2804 1072 2805 1112
rect 2763 1063 2805 1072
rect 2668 944 2708 953
rect 2860 944 2900 1660
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 3532 1364 3572 1660
rect 3244 1324 3572 1364
rect 2955 1196 2997 1205
rect 2955 1156 2956 1196
rect 2996 1156 2997 1196
rect 2955 1147 2997 1156
rect 2956 1112 2996 1147
rect 3148 1121 3188 1206
rect 2956 1061 2996 1072
rect 3147 1112 3189 1121
rect 3147 1072 3148 1112
rect 3188 1072 3189 1112
rect 3147 1063 3189 1072
rect 3052 944 3092 953
rect 2380 484 2516 524
rect 2572 904 2668 944
rect 2380 80 2420 484
rect 2572 80 2612 904
rect 2668 895 2708 904
rect 2764 904 2900 944
rect 2956 904 3052 944
rect 2764 80 2804 904
rect 2956 80 2996 904
rect 3052 895 3092 904
rect 3244 776 3284 1324
rect 3339 1196 3381 1205
rect 3339 1156 3340 1196
rect 3380 1156 3381 1196
rect 3339 1147 3381 1156
rect 3340 1112 3380 1147
rect 3532 1121 3572 1206
rect 3340 1061 3380 1072
rect 3531 1112 3573 1121
rect 3531 1072 3532 1112
rect 3572 1072 3573 1112
rect 3531 1063 3573 1072
rect 3436 944 3476 953
rect 3628 944 3668 1912
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 3724 1112 3764 1231
rect 3916 1121 3956 1206
rect 3724 1063 3764 1072
rect 3915 1112 3957 1121
rect 3915 1072 3916 1112
rect 3956 1072 3957 1112
rect 3915 1063 3957 1072
rect 3820 944 3860 953
rect 4012 944 4052 2500
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 5068 1289 5108 3172
rect 5740 3053 5780 3424
rect 5931 3464 5973 3473
rect 5931 3424 5932 3464
rect 5972 3424 5973 3464
rect 5931 3415 5973 3424
rect 5932 3330 5972 3415
rect 5836 3212 5876 3221
rect 5739 3044 5781 3053
rect 5739 3004 5740 3044
rect 5780 3004 5781 3044
rect 5739 2995 5781 3004
rect 5740 2633 5780 2995
rect 5355 2624 5397 2633
rect 5355 2584 5356 2624
rect 5396 2584 5397 2624
rect 5355 2575 5397 2584
rect 5739 2624 5781 2633
rect 5739 2584 5740 2624
rect 5780 2584 5781 2624
rect 5739 2575 5781 2584
rect 5356 1952 5396 2575
rect 5547 2288 5589 2297
rect 5547 2248 5548 2288
rect 5588 2248 5589 2288
rect 5547 2239 5589 2248
rect 5356 1903 5396 1912
rect 5548 1952 5588 2239
rect 5548 1903 5588 1912
rect 5452 1700 5492 1709
rect 5164 1660 5452 1700
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 5067 1280 5109 1289
rect 5067 1240 5068 1280
rect 5108 1240 5109 1280
rect 5067 1231 5109 1240
rect 4108 1125 4148 1231
rect 4300 1121 4340 1206
rect 4491 1196 4533 1205
rect 4491 1156 4492 1196
rect 4532 1156 4533 1196
rect 4491 1147 4533 1156
rect 4493 1125 4533 1147
rect 4108 1076 4148 1085
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 4684 1121 4724 1206
rect 4875 1196 4917 1205
rect 4875 1156 4876 1196
rect 4916 1156 4917 1196
rect 4875 1147 4917 1156
rect 4493 1062 4533 1085
rect 4683 1112 4725 1121
rect 4683 1072 4684 1112
rect 4724 1072 4725 1112
rect 4683 1063 4725 1072
rect 4876 1112 4916 1147
rect 4876 1061 4916 1072
rect 5068 1112 5108 1121
rect 4204 944 4244 953
rect 3145 736 3284 776
rect 3340 904 3436 944
rect 3145 692 3185 736
rect 3145 652 3188 692
rect 3148 80 3188 652
rect 3340 80 3380 904
rect 3436 895 3476 904
rect 3532 904 3668 944
rect 3724 904 3820 944
rect 3532 80 3572 904
rect 3724 80 3764 904
rect 3820 895 3860 904
rect 3916 904 4052 944
rect 4108 904 4204 944
rect 3916 80 3956 904
rect 4108 80 4148 904
rect 4204 895 4244 904
rect 4588 944 4628 953
rect 4972 944 5012 953
rect 4628 904 4820 944
rect 4588 895 4628 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 4299 608 4341 617
rect 4299 568 4300 608
rect 4340 568 4341 608
rect 4299 559 4341 568
rect 4300 80 4340 559
rect 4780 524 4820 904
rect 4492 484 4820 524
rect 4876 904 4972 944
rect 4492 80 4532 484
rect 4683 356 4725 365
rect 4683 316 4684 356
rect 4724 316 4725 356
rect 4683 307 4725 316
rect 4684 80 4724 307
rect 4876 80 4916 904
rect 4972 895 5012 904
rect 5068 617 5108 1072
rect 5067 608 5109 617
rect 5067 568 5068 608
rect 5108 568 5109 608
rect 5067 559 5109 568
rect 5164 188 5204 1660
rect 5452 1651 5492 1660
rect 5836 1364 5876 3172
rect 6412 3137 6452 3499
rect 6699 3464 6741 3473
rect 6699 3424 6700 3464
rect 6740 3424 6741 3464
rect 6699 3415 6741 3424
rect 6891 3464 6933 3473
rect 6891 3424 6892 3464
rect 6932 3424 6933 3464
rect 6891 3415 6933 3424
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 6411 3128 6453 3137
rect 6411 3088 6412 3128
rect 6452 3088 6453 3128
rect 6411 3079 6453 3088
rect 6315 3044 6357 3053
rect 6315 3004 6316 3044
rect 6356 3004 6357 3044
rect 6315 2995 6357 3004
rect 6123 2624 6165 2633
rect 6123 2584 6124 2624
rect 6164 2584 6165 2624
rect 6123 2575 6165 2584
rect 6316 2624 6356 2995
rect 6316 2575 6356 2584
rect 6124 2490 6164 2575
rect 6220 2540 6260 2549
rect 6220 1373 6260 2500
rect 6412 2465 6452 3079
rect 6700 2969 6740 3415
rect 6892 3330 6932 3415
rect 7084 3330 7124 3415
rect 6988 3212 7028 3221
rect 6892 3172 6988 3212
rect 6795 3128 6837 3137
rect 6795 3088 6796 3128
rect 6836 3088 6837 3128
rect 6795 3079 6837 3088
rect 6699 2960 6741 2969
rect 6699 2920 6700 2960
rect 6740 2920 6741 2960
rect 6699 2911 6741 2920
rect 6603 2624 6645 2633
rect 6603 2584 6604 2624
rect 6644 2584 6645 2624
rect 6603 2575 6645 2584
rect 6796 2624 6836 3079
rect 6796 2575 6836 2584
rect 6604 2490 6644 2575
rect 6700 2540 6740 2549
rect 6411 2456 6453 2465
rect 6411 2416 6412 2456
rect 6452 2416 6453 2456
rect 6411 2407 6453 2416
rect 6411 2036 6453 2045
rect 6411 1996 6412 2036
rect 6452 1996 6453 2036
rect 6411 1987 6453 1996
rect 5548 1324 5876 1364
rect 6219 1364 6261 1373
rect 6219 1324 6220 1364
rect 6260 1324 6261 1364
rect 5259 1196 5301 1205
rect 5259 1156 5260 1196
rect 5300 1156 5301 1196
rect 5259 1147 5301 1156
rect 5260 1112 5300 1147
rect 5260 1061 5300 1072
rect 5452 1112 5492 1121
rect 5356 1028 5396 1037
rect 5452 1028 5492 1072
rect 5356 944 5396 988
rect 5068 148 5204 188
rect 5260 904 5396 944
rect 5445 988 5492 1028
rect 5548 1028 5588 1324
rect 6219 1315 6261 1324
rect 6412 1205 6452 1987
rect 6700 1289 6740 2500
rect 6795 2036 6837 2045
rect 6795 1996 6796 2036
rect 6836 1996 6837 2036
rect 6795 1987 6837 1996
rect 6796 1952 6836 1987
rect 6796 1901 6836 1912
rect 6796 1700 6836 1709
rect 6796 1457 6836 1660
rect 6795 1448 6837 1457
rect 6795 1408 6796 1448
rect 6836 1408 6837 1448
rect 6795 1399 6837 1408
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 5643 1196 5685 1205
rect 5643 1156 5644 1196
rect 5684 1156 5685 1196
rect 5643 1147 5685 1156
rect 6123 1196 6165 1205
rect 6123 1156 6124 1196
rect 6164 1156 6165 1196
rect 6123 1147 6165 1156
rect 6411 1196 6453 1205
rect 6411 1156 6412 1196
rect 6452 1156 6453 1196
rect 6411 1147 6453 1156
rect 5644 1112 5684 1147
rect 5644 1061 5684 1072
rect 5836 1112 5876 1121
rect 5876 1072 5972 1112
rect 5836 1063 5876 1072
rect 5548 988 5591 1028
rect 5068 80 5108 148
rect 5260 80 5300 904
rect 5445 860 5485 988
rect 5356 820 5485 860
rect 5356 701 5396 820
rect 5551 776 5591 988
rect 5740 944 5780 953
rect 5452 736 5591 776
rect 5644 904 5740 944
rect 5355 692 5397 701
rect 5355 652 5356 692
rect 5396 652 5397 692
rect 5355 643 5397 652
rect 5452 80 5492 736
rect 5644 80 5684 904
rect 5740 895 5780 904
rect 5835 524 5877 533
rect 5835 484 5836 524
rect 5876 484 5877 524
rect 5835 475 5877 484
rect 5836 80 5876 475
rect 5932 281 5972 1072
rect 6038 1101 6078 1110
rect 6124 1101 6164 1147
rect 6412 1112 6452 1147
rect 6078 1061 6164 1101
rect 6217 1101 6257 1110
rect 6412 1063 6452 1072
rect 6507 1112 6549 1121
rect 6604 1112 6644 1121
rect 6507 1072 6508 1112
rect 6548 1072 6604 1112
rect 6507 1063 6549 1072
rect 6604 1063 6644 1072
rect 6807 1101 6847 1110
rect 6038 1052 6078 1061
rect 6217 1028 6257 1061
rect 6217 988 6260 1028
rect 6124 944 6164 953
rect 6028 904 6124 944
rect 5931 272 5973 281
rect 5931 232 5932 272
rect 5972 232 5973 272
rect 5931 223 5973 232
rect 6028 80 6068 904
rect 6124 895 6164 904
rect 6220 785 6260 988
rect 6807 953 6847 1061
rect 6892 1028 6932 3172
rect 6988 3163 7028 3172
rect 7180 2960 7220 3592
rect 7276 3557 7316 3580
rect 7275 3548 7317 3557
rect 7275 3508 7276 3548
rect 7316 3508 7317 3548
rect 7275 3499 7317 3508
rect 7276 3485 7316 3499
rect 7276 3436 7316 3445
rect 7372 3380 7412 3928
rect 9195 3800 9237 3809
rect 9195 3760 9196 3800
rect 9236 3760 9237 3800
rect 9195 3751 9237 3760
rect 15243 3800 15285 3809
rect 15243 3760 15244 3800
rect 15284 3760 15285 3800
rect 15243 3751 15285 3760
rect 8427 3716 8469 3725
rect 8427 3676 8428 3716
rect 8468 3676 8469 3716
rect 8427 3667 8469 3676
rect 7467 3464 7509 3473
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7660 3464 7700 3473
rect 6988 2920 7220 2960
rect 7276 3340 7412 3380
rect 6988 2633 7028 2920
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 6988 2490 7028 2575
rect 7083 2540 7125 2549
rect 7083 2500 7084 2540
rect 7124 2500 7125 2540
rect 7083 2491 7125 2500
rect 7084 2406 7124 2491
rect 7180 2490 7220 2575
rect 6987 2120 7029 2129
rect 6987 2080 6988 2120
rect 7028 2080 7029 2120
rect 6987 2071 7029 2080
rect 6988 1952 7028 2071
rect 7276 2045 7316 3340
rect 7468 3330 7508 3415
rect 7372 3212 7412 3221
rect 7412 3172 7508 3212
rect 7372 3163 7412 3172
rect 7275 2036 7317 2045
rect 7275 1996 7276 2036
rect 7316 1996 7317 2036
rect 7275 1987 7317 1996
rect 6988 1903 7028 1912
rect 6988 1364 7028 1373
rect 7028 1324 7124 1364
rect 6988 1315 7028 1324
rect 6988 1205 7028 1213
rect 6987 1196 7029 1205
rect 6987 1156 6988 1196
rect 7028 1156 7035 1196
rect 6987 1147 7035 1156
rect 6995 1125 7035 1147
rect 6995 1076 7035 1085
rect 6892 988 7028 1028
rect 6411 944 6453 953
rect 6411 904 6412 944
rect 6452 904 6453 944
rect 6411 895 6453 904
rect 6508 944 6548 953
rect 6219 776 6261 785
rect 6219 736 6220 776
rect 6260 736 6261 776
rect 6219 727 6261 736
rect 6219 524 6261 533
rect 6219 484 6220 524
rect 6260 484 6261 524
rect 6219 475 6261 484
rect 6220 80 6260 475
rect 6412 80 6452 895
rect 6508 365 6548 904
rect 6806 944 6848 953
rect 6806 904 6807 944
rect 6847 904 6848 944
rect 6806 895 6848 904
rect 6507 356 6549 365
rect 6507 316 6508 356
rect 6548 316 6549 356
rect 6507 307 6549 316
rect 6795 356 6837 365
rect 6795 316 6796 356
rect 6836 316 6837 356
rect 6795 307 6837 316
rect 6603 188 6645 197
rect 6603 148 6604 188
rect 6644 148 6645 188
rect 6603 139 6645 148
rect 6604 80 6644 139
rect 6796 80 6836 307
rect 6988 80 7028 988
rect 7084 524 7124 1324
rect 7179 1196 7221 1205
rect 7179 1156 7180 1196
rect 7220 1156 7221 1196
rect 7179 1147 7221 1156
rect 7371 1196 7413 1205
rect 7371 1156 7372 1196
rect 7412 1156 7413 1196
rect 7371 1147 7413 1156
rect 7180 1112 7220 1147
rect 7180 1061 7220 1072
rect 7372 1112 7412 1147
rect 7372 1061 7412 1072
rect 7275 944 7317 953
rect 7468 944 7508 3172
rect 7660 2969 7700 3424
rect 7851 3464 7893 3473
rect 7851 3424 7852 3464
rect 7892 3424 7893 3464
rect 7851 3415 7893 3424
rect 8235 3464 8277 3473
rect 8235 3424 8236 3464
rect 8276 3424 8277 3464
rect 8235 3415 8277 3424
rect 8428 3464 8468 3667
rect 7852 3330 7892 3415
rect 7756 3212 7796 3221
rect 7796 3172 7892 3212
rect 7756 3163 7796 3172
rect 7659 2960 7701 2969
rect 7659 2920 7660 2960
rect 7700 2920 7701 2960
rect 7659 2911 7701 2920
rect 7564 1205 7604 1207
rect 7563 1196 7605 1205
rect 7563 1156 7564 1196
rect 7604 1156 7605 1196
rect 7563 1147 7605 1156
rect 7564 1112 7604 1147
rect 7756 1121 7796 1206
rect 7564 1063 7604 1072
rect 7755 1112 7797 1121
rect 7755 1072 7756 1112
rect 7796 1072 7797 1112
rect 7755 1063 7797 1072
rect 7275 904 7276 944
rect 7316 904 7317 944
rect 7275 895 7317 904
rect 7372 904 7508 944
rect 7563 944 7605 953
rect 7563 904 7564 944
rect 7604 904 7605 944
rect 7276 810 7316 895
rect 7084 484 7220 524
rect 7180 80 7220 484
rect 7372 80 7412 904
rect 7563 895 7605 904
rect 7660 944 7700 953
rect 7852 944 7892 3172
rect 8043 2624 8085 2633
rect 8043 2584 8044 2624
rect 8084 2584 8085 2624
rect 8043 2575 8085 2584
rect 8236 2624 8276 3415
rect 8428 3305 8468 3424
rect 8619 3464 8661 3473
rect 8619 3424 8620 3464
rect 8660 3424 8661 3464
rect 8619 3415 8661 3424
rect 8812 3464 8852 3473
rect 8620 3330 8660 3415
rect 8427 3296 8469 3305
rect 8427 3256 8428 3296
rect 8468 3256 8469 3296
rect 8427 3247 8469 3256
rect 8524 3212 8564 3221
rect 8564 3172 8660 3212
rect 8524 3163 8564 3172
rect 8236 2575 8276 2584
rect 8044 2490 8084 2575
rect 8140 2540 8180 2549
rect 8140 1364 8180 2500
rect 8140 1324 8276 1364
rect 8140 1121 8180 1206
rect 7564 80 7604 895
rect 7660 533 7700 904
rect 7756 904 7892 944
rect 7948 1112 7988 1121
rect 7659 524 7701 533
rect 7659 484 7660 524
rect 7700 484 7701 524
rect 7659 475 7701 484
rect 7756 80 7796 904
rect 7948 860 7988 1072
rect 8139 1112 8181 1121
rect 8139 1072 8140 1112
rect 8180 1072 8181 1112
rect 8139 1063 8181 1072
rect 8043 944 8085 953
rect 8236 944 8276 1324
rect 8332 1205 8372 1207
rect 8331 1196 8373 1205
rect 8331 1156 8332 1196
rect 8372 1156 8373 1196
rect 8331 1147 8373 1156
rect 8523 1196 8565 1205
rect 8523 1156 8524 1196
rect 8564 1156 8565 1196
rect 8523 1147 8565 1156
rect 8332 1112 8372 1147
rect 8332 1063 8372 1072
rect 8524 1112 8564 1147
rect 8524 1061 8564 1072
rect 8043 904 8044 944
rect 8084 904 8085 944
rect 8043 895 8085 904
rect 8140 904 8276 944
rect 8331 944 8373 953
rect 8331 904 8332 944
rect 8372 904 8373 944
rect 7852 820 7988 860
rect 7852 281 7892 820
rect 8044 810 8084 895
rect 7947 524 7989 533
rect 7947 484 7948 524
rect 7988 484 7989 524
rect 7947 475 7989 484
rect 7851 272 7893 281
rect 7851 232 7852 272
rect 7892 232 7893 272
rect 7851 223 7893 232
rect 7948 80 7988 475
rect 8140 80 8180 904
rect 8331 895 8373 904
rect 8428 944 8468 953
rect 8620 944 8660 3172
rect 8812 2801 8852 3424
rect 9003 3464 9045 3473
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9196 3464 9236 3751
rect 12075 3716 12117 3725
rect 12075 3676 12076 3716
rect 12116 3676 12117 3716
rect 12075 3667 12117 3676
rect 12459 3716 12501 3725
rect 12459 3676 12460 3716
rect 12500 3676 12501 3716
rect 12459 3667 12501 3676
rect 10155 3632 10197 3641
rect 10155 3592 10156 3632
rect 10196 3592 10197 3632
rect 10155 3583 10197 3592
rect 10539 3632 10581 3641
rect 10539 3592 10540 3632
rect 10580 3592 10581 3632
rect 10539 3583 10581 3592
rect 10923 3632 10965 3641
rect 10923 3592 10924 3632
rect 10964 3592 10965 3632
rect 10923 3583 10965 3592
rect 11307 3632 11349 3641
rect 11307 3592 11308 3632
rect 11348 3592 11349 3632
rect 11307 3583 11349 3592
rect 11691 3632 11733 3641
rect 11691 3592 11692 3632
rect 11732 3592 11733 3632
rect 11691 3583 11733 3592
rect 9579 3548 9621 3557
rect 9579 3508 9580 3548
rect 9620 3508 9621 3548
rect 9579 3499 9621 3508
rect 9963 3548 10005 3557
rect 9963 3508 9964 3548
rect 10004 3508 10005 3548
rect 9963 3499 10005 3508
rect 9004 3330 9044 3415
rect 8908 3212 8948 3221
rect 8948 3172 9044 3212
rect 8908 3163 8948 3172
rect 8811 2792 8853 2801
rect 8811 2752 8812 2792
rect 8852 2752 8853 2792
rect 8811 2743 8853 2752
rect 8907 1196 8949 1205
rect 8907 1156 8908 1196
rect 8948 1156 8949 1196
rect 8907 1147 8949 1156
rect 8332 80 8372 895
rect 8428 533 8468 904
rect 8524 904 8660 944
rect 8716 1112 8756 1121
rect 8427 524 8469 533
rect 8427 484 8428 524
rect 8468 484 8469 524
rect 8427 475 8469 484
rect 8524 80 8564 904
rect 8716 860 8756 1072
rect 8908 1112 8948 1147
rect 8908 1061 8948 1072
rect 8811 944 8853 953
rect 9004 944 9044 3172
rect 9196 2717 9236 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 9580 3464 9620 3499
rect 9388 3330 9428 3415
rect 9580 3413 9620 3424
rect 9771 3464 9813 3473
rect 9771 3424 9772 3464
rect 9812 3424 9813 3464
rect 9771 3415 9813 3424
rect 9964 3464 10004 3499
rect 10156 3473 10196 3583
rect 9772 3330 9812 3415
rect 9964 3413 10004 3424
rect 10155 3464 10197 3473
rect 10155 3424 10156 3464
rect 10196 3424 10197 3464
rect 10155 3415 10197 3424
rect 10348 3464 10388 3473
rect 10156 3330 10196 3415
rect 10348 3305 10388 3424
rect 10540 3464 10580 3583
rect 10540 3415 10580 3424
rect 10732 3464 10772 3475
rect 10732 3389 10772 3424
rect 10924 3464 10964 3583
rect 10924 3415 10964 3424
rect 11115 3464 11157 3473
rect 11115 3424 11116 3464
rect 11156 3424 11157 3464
rect 11115 3415 11157 3424
rect 11308 3464 11348 3583
rect 11692 3473 11732 3583
rect 12076 3473 12116 3667
rect 11308 3415 11348 3424
rect 11499 3464 11541 3473
rect 11499 3424 11500 3464
rect 11540 3424 11541 3464
rect 11499 3415 11541 3424
rect 11691 3464 11733 3473
rect 11691 3424 11692 3464
rect 11732 3424 11733 3464
rect 11691 3415 11733 3424
rect 11884 3464 11924 3473
rect 10731 3380 10773 3389
rect 10731 3340 10732 3380
rect 10772 3340 10773 3380
rect 10731 3331 10773 3340
rect 10347 3296 10389 3305
rect 10347 3256 10348 3296
rect 10388 3256 10389 3296
rect 10347 3247 10389 3256
rect 9292 3212 9332 3221
rect 9676 3212 9716 3221
rect 10060 3212 10100 3221
rect 9332 3172 9428 3212
rect 9292 3163 9332 3172
rect 9195 2708 9237 2717
rect 9195 2668 9196 2708
rect 9236 2668 9237 2708
rect 9195 2659 9237 2668
rect 9099 1280 9141 1289
rect 9099 1240 9100 1280
rect 9140 1240 9141 1280
rect 9099 1231 9141 1240
rect 9100 1121 9140 1231
rect 9291 1196 9333 1205
rect 9291 1156 9292 1196
rect 9332 1156 9333 1196
rect 9291 1147 9333 1156
rect 9099 1112 9141 1121
rect 9099 1072 9100 1112
rect 9140 1072 9141 1112
rect 9099 1063 9141 1072
rect 9292 1112 9332 1147
rect 9292 1061 9332 1072
rect 8811 904 8812 944
rect 8852 904 8853 944
rect 8811 895 8853 904
rect 8908 904 9044 944
rect 9099 944 9141 953
rect 9099 904 9100 944
rect 9140 904 9141 944
rect 8620 820 8756 860
rect 8620 449 8660 820
rect 8812 810 8852 895
rect 8715 524 8757 533
rect 8715 484 8716 524
rect 8756 484 8757 524
rect 8715 475 8757 484
rect 8619 440 8661 449
rect 8619 400 8620 440
rect 8660 400 8661 440
rect 8619 391 8661 400
rect 8716 80 8756 475
rect 8908 80 8948 904
rect 9099 895 9141 904
rect 9196 944 9236 953
rect 9388 944 9428 3172
rect 9716 3172 9812 3212
rect 9676 3163 9716 3172
rect 9675 1196 9717 1205
rect 9675 1156 9676 1196
rect 9716 1156 9717 1196
rect 9675 1147 9717 1156
rect 9484 1112 9524 1121
rect 9484 1037 9524 1072
rect 9676 1112 9716 1147
rect 9676 1061 9716 1072
rect 9483 1028 9525 1037
rect 9483 988 9484 1028
rect 9524 988 9525 1028
rect 9483 979 9525 988
rect 9100 80 9140 895
rect 9196 533 9236 904
rect 9292 904 9428 944
rect 9195 524 9237 533
rect 9195 484 9196 524
rect 9236 484 9237 524
rect 9195 475 9237 484
rect 9292 80 9332 904
rect 9484 869 9524 979
rect 9579 944 9621 953
rect 9772 944 9812 3172
rect 10060 2540 10100 3172
rect 10444 3212 10484 3221
rect 10828 3212 10868 3221
rect 10484 3172 10580 3212
rect 10444 3163 10484 3172
rect 10060 2500 10196 2540
rect 9868 1121 9908 1206
rect 10059 1196 10101 1205
rect 10059 1156 10060 1196
rect 10100 1156 10101 1196
rect 10059 1147 10101 1156
rect 9867 1112 9909 1121
rect 9867 1072 9868 1112
rect 9908 1072 9909 1112
rect 9867 1063 9909 1072
rect 10060 1112 10100 1147
rect 10060 1061 10100 1072
rect 9579 904 9580 944
rect 9620 904 9621 944
rect 9579 895 9621 904
rect 9676 904 9812 944
rect 9867 944 9909 953
rect 9867 904 9868 944
rect 9908 904 9909 944
rect 9483 860 9525 869
rect 9483 820 9484 860
rect 9524 820 9525 860
rect 9483 811 9525 820
rect 9580 810 9620 895
rect 9483 524 9525 533
rect 9483 484 9484 524
rect 9524 484 9525 524
rect 9483 475 9525 484
rect 9484 80 9524 475
rect 9676 80 9716 904
rect 9867 895 9909 904
rect 9964 944 10004 953
rect 10156 944 10196 2500
rect 10443 1196 10485 1205
rect 10443 1156 10444 1196
rect 10484 1156 10485 1196
rect 10443 1147 10485 1156
rect 10251 1112 10293 1121
rect 10251 1072 10252 1112
rect 10292 1072 10293 1112
rect 10251 1063 10293 1072
rect 10444 1112 10484 1147
rect 10252 978 10292 1063
rect 10444 1061 10484 1072
rect 9868 80 9908 895
rect 9964 533 10004 904
rect 10060 904 10196 944
rect 10347 944 10389 953
rect 10540 944 10580 3172
rect 10868 3172 10964 3212
rect 10828 3163 10868 3172
rect 10636 1121 10676 1206
rect 10827 1196 10869 1205
rect 10827 1156 10828 1196
rect 10868 1156 10869 1196
rect 10827 1147 10869 1156
rect 10635 1112 10677 1121
rect 10635 1072 10636 1112
rect 10676 1072 10677 1112
rect 10635 1063 10677 1072
rect 10828 1112 10868 1147
rect 10828 1061 10868 1072
rect 10347 904 10348 944
rect 10388 904 10389 944
rect 9963 524 10005 533
rect 9963 484 9964 524
rect 10004 484 10005 524
rect 9963 475 10005 484
rect 10060 80 10100 904
rect 10347 895 10389 904
rect 10444 904 10580 944
rect 10635 944 10677 953
rect 10635 904 10636 944
rect 10676 904 10677 944
rect 10348 810 10388 895
rect 10251 524 10293 533
rect 10251 484 10252 524
rect 10292 484 10293 524
rect 10251 475 10293 484
rect 10252 80 10292 475
rect 10444 80 10484 904
rect 10635 895 10677 904
rect 10732 944 10772 953
rect 10924 944 10964 3172
rect 11116 2297 11156 3415
rect 11500 3330 11540 3415
rect 11691 3296 11733 3305
rect 11691 3256 11692 3296
rect 11732 3256 11733 3296
rect 11691 3247 11733 3256
rect 11212 3212 11252 3221
rect 11596 3212 11636 3221
rect 11252 3172 11348 3212
rect 11212 3163 11252 3172
rect 11115 2288 11157 2297
rect 11115 2248 11116 2288
rect 11156 2248 11157 2288
rect 11115 2239 11157 2248
rect 11211 1196 11253 1205
rect 11211 1156 11212 1196
rect 11252 1156 11253 1196
rect 11211 1147 11253 1156
rect 10636 80 10676 895
rect 10732 281 10772 904
rect 10828 904 10964 944
rect 11020 1112 11060 1121
rect 10731 272 10773 281
rect 10731 232 10732 272
rect 10772 232 10773 272
rect 10731 223 10773 232
rect 10828 80 10868 904
rect 11020 701 11060 1072
rect 11212 1112 11252 1147
rect 11212 1061 11252 1072
rect 11115 944 11157 953
rect 11308 944 11348 3172
rect 11596 2540 11636 3172
rect 11692 2885 11732 3247
rect 11884 3221 11924 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 12268 3464 12308 3473
rect 12076 3330 12116 3415
rect 12268 3305 12308 3424
rect 12460 3464 12500 3667
rect 15244 3641 15284 3751
rect 16779 3716 16821 3725
rect 16779 3676 16780 3716
rect 16820 3676 16821 3716
rect 16779 3667 16821 3676
rect 14475 3632 14517 3641
rect 14475 3592 14476 3632
rect 14516 3592 14517 3632
rect 14475 3583 14517 3592
rect 15243 3632 15285 3641
rect 15243 3592 15244 3632
rect 15284 3592 15285 3632
rect 15243 3583 15285 3592
rect 13227 3548 13269 3557
rect 13227 3508 13228 3548
rect 13268 3508 13269 3548
rect 13227 3499 13269 3508
rect 13611 3548 13653 3557
rect 13611 3508 13612 3548
rect 13652 3508 13653 3548
rect 13611 3499 13653 3508
rect 13995 3548 14037 3557
rect 13995 3508 13996 3548
rect 14036 3508 14037 3548
rect 13995 3499 14037 3508
rect 14283 3548 14325 3557
rect 14283 3508 14284 3548
rect 14324 3508 14325 3548
rect 14283 3499 14325 3508
rect 13035 3464 13077 3473
rect 12500 3424 12596 3464
rect 12460 3415 12500 3424
rect 12267 3296 12309 3305
rect 12267 3256 12268 3296
rect 12308 3256 12309 3296
rect 12267 3247 12309 3256
rect 11883 3212 11925 3221
rect 11883 3172 11884 3212
rect 11924 3172 11925 3212
rect 11883 3163 11925 3172
rect 11980 3212 12020 3221
rect 11691 2876 11733 2885
rect 11691 2836 11692 2876
rect 11732 2836 11733 2876
rect 11691 2827 11733 2836
rect 11980 2540 12020 3172
rect 12268 3137 12308 3247
rect 12364 3212 12404 3221
rect 12267 3128 12309 3137
rect 12267 3088 12268 3128
rect 12308 3088 12309 3128
rect 12267 3079 12309 3088
rect 12364 2540 12404 3172
rect 12556 2624 12596 3424
rect 13035 3424 13036 3464
rect 13076 3424 13077 3464
rect 13035 3415 13077 3424
rect 13228 3464 13268 3499
rect 13036 3330 13076 3415
rect 13228 3413 13268 3424
rect 13420 3464 13460 3473
rect 13132 3212 13172 3221
rect 12748 2633 12788 2718
rect 12556 2575 12596 2584
rect 12747 2624 12789 2633
rect 12747 2584 12748 2624
rect 12788 2584 12789 2624
rect 12747 2575 12789 2584
rect 12652 2540 12692 2549
rect 11596 2500 11732 2540
rect 11980 2500 12116 2540
rect 12364 2500 12500 2540
rect 11596 1205 11636 1220
rect 11595 1196 11637 1205
rect 11595 1156 11596 1196
rect 11636 1156 11637 1196
rect 11595 1147 11637 1156
rect 11596 1125 11636 1147
rect 11404 1112 11444 1121
rect 11499 1112 11541 1121
rect 11444 1072 11500 1112
rect 11540 1072 11541 1112
rect 11596 1076 11636 1085
rect 11404 1063 11444 1072
rect 11499 1063 11541 1072
rect 11692 1028 11732 2500
rect 11979 1196 12021 1205
rect 11979 1156 11980 1196
rect 12020 1156 12021 1196
rect 11979 1147 12021 1156
rect 11596 988 11732 1028
rect 11788 1112 11828 1121
rect 11115 904 11116 944
rect 11156 904 11157 944
rect 11115 895 11157 904
rect 11212 904 11348 944
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11116 810 11156 895
rect 11019 692 11061 701
rect 11019 652 11020 692
rect 11060 652 11061 692
rect 11019 643 11061 652
rect 11020 449 11060 643
rect 11019 440 11061 449
rect 11019 400 11020 440
rect 11060 400 11061 440
rect 11019 391 11061 400
rect 11019 272 11061 281
rect 11019 232 11020 272
rect 11060 232 11061 272
rect 11019 223 11061 232
rect 11020 80 11060 223
rect 11212 80 11252 904
rect 11403 895 11445 904
rect 11500 944 11540 953
rect 11404 80 11444 895
rect 11500 197 11540 904
rect 11499 188 11541 197
rect 11499 148 11500 188
rect 11540 148 11541 188
rect 11499 139 11541 148
rect 11596 80 11636 988
rect 11788 944 11828 1072
rect 11980 1112 12020 1147
rect 11980 1061 12020 1072
rect 11884 944 11924 953
rect 12076 944 12116 2500
rect 12171 2120 12213 2129
rect 12171 2080 12172 2120
rect 12212 2080 12213 2120
rect 12171 2071 12213 2080
rect 12172 1121 12212 2071
rect 12363 1196 12405 1205
rect 12363 1156 12364 1196
rect 12404 1156 12405 1196
rect 12363 1147 12405 1156
rect 12171 1112 12213 1121
rect 12171 1072 12172 1112
rect 12212 1072 12213 1112
rect 12171 1063 12213 1072
rect 12364 1112 12404 1147
rect 12172 978 12212 1063
rect 12364 1061 12404 1072
rect 11788 904 11831 944
rect 11692 869 11732 888
rect 11691 860 11733 869
rect 11791 860 11831 904
rect 11691 820 11692 860
rect 11732 820 11831 860
rect 11691 811 11733 820
rect 11788 449 11828 820
rect 11884 533 11924 904
rect 11980 904 12116 944
rect 12267 944 12309 953
rect 12460 944 12500 2500
rect 13132 2540 13172 3172
rect 13132 2500 13268 2540
rect 12652 1364 12692 2500
rect 13035 1616 13077 1625
rect 13035 1576 13036 1616
rect 13076 1576 13077 1616
rect 13035 1567 13077 1576
rect 12652 1324 12884 1364
rect 12556 1121 12596 1206
rect 12651 1196 12693 1205
rect 12651 1156 12652 1196
rect 12692 1156 12788 1196
rect 12651 1147 12693 1156
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12748 1109 12788 1156
rect 12748 1060 12788 1069
rect 12267 904 12268 944
rect 12308 904 12309 944
rect 11883 524 11925 533
rect 11883 484 11884 524
rect 11924 484 11925 524
rect 11883 475 11925 484
rect 11787 440 11829 449
rect 11787 400 11788 440
rect 11828 400 11829 440
rect 11787 391 11829 400
rect 11787 188 11829 197
rect 11787 148 11788 188
rect 11828 148 11829 188
rect 11787 139 11829 148
rect 11788 80 11828 139
rect 11980 80 12020 904
rect 12267 895 12309 904
rect 12364 904 12500 944
rect 12555 944 12597 953
rect 12555 904 12556 944
rect 12596 904 12597 944
rect 12268 810 12308 895
rect 12171 524 12213 533
rect 12171 484 12172 524
rect 12212 484 12213 524
rect 12171 475 12213 484
rect 12172 80 12212 475
rect 12364 80 12404 904
rect 12555 895 12597 904
rect 12652 944 12692 953
rect 12844 944 12884 1324
rect 12940 1121 12980 1206
rect 13036 1205 13076 1567
rect 13035 1196 13077 1205
rect 13035 1156 13036 1196
rect 13076 1156 13077 1196
rect 13035 1147 13077 1156
rect 13132 1121 13172 1206
rect 12939 1112 12981 1121
rect 12939 1072 12940 1112
rect 12980 1072 12981 1112
rect 12939 1063 12981 1072
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 13131 1063 13173 1072
rect 12556 80 12596 895
rect 12652 533 12692 904
rect 12748 904 12884 944
rect 13035 944 13077 953
rect 13228 944 13268 2500
rect 13420 2465 13460 3424
rect 13612 3464 13652 3499
rect 13612 3413 13652 3424
rect 13804 3464 13844 3473
rect 13516 3212 13556 3221
rect 13516 2540 13556 3172
rect 13804 2969 13844 3424
rect 13996 3464 14036 3499
rect 13900 3212 13940 3221
rect 13803 2960 13845 2969
rect 13803 2920 13804 2960
rect 13844 2920 13845 2960
rect 13803 2911 13845 2920
rect 13516 2500 13652 2540
rect 13419 2456 13461 2465
rect 13419 2416 13420 2456
rect 13460 2416 13461 2456
rect 13419 2407 13461 2416
rect 13324 1205 13364 1207
rect 13323 1196 13365 1205
rect 13323 1156 13324 1196
rect 13364 1156 13365 1196
rect 13323 1147 13365 1156
rect 13324 1112 13364 1147
rect 13516 1121 13556 1206
rect 13324 1063 13364 1072
rect 13515 1112 13557 1121
rect 13515 1072 13516 1112
rect 13556 1072 13557 1112
rect 13515 1063 13557 1072
rect 13035 904 13036 944
rect 13076 904 13077 944
rect 12651 524 12693 533
rect 12651 484 12652 524
rect 12692 484 12693 524
rect 12651 475 12693 484
rect 12748 80 12788 904
rect 13035 895 13077 904
rect 13132 904 13268 944
rect 13323 944 13365 953
rect 13323 904 13324 944
rect 13364 904 13365 944
rect 13036 810 13076 895
rect 12939 524 12981 533
rect 12939 484 12940 524
rect 12980 484 12981 524
rect 12939 475 12981 484
rect 12940 80 12980 475
rect 13132 80 13172 904
rect 13323 895 13365 904
rect 13420 944 13460 953
rect 13612 944 13652 2500
rect 13804 2465 13844 2911
rect 13900 2540 13940 3172
rect 13996 2624 14036 3424
rect 14284 3464 14324 3499
rect 14284 3413 14324 3424
rect 14476 3464 14516 3583
rect 14667 3548 14709 3557
rect 14667 3508 14668 3548
rect 14708 3508 14709 3548
rect 14667 3499 14709 3508
rect 15051 3548 15093 3557
rect 15051 3508 15052 3548
rect 15092 3508 15093 3548
rect 15051 3499 15093 3508
rect 14380 3212 14420 3221
rect 14284 2717 14324 2719
rect 14283 2708 14325 2717
rect 14283 2668 14284 2708
rect 14324 2668 14325 2708
rect 14283 2659 14325 2668
rect 14092 2624 14132 2633
rect 13996 2584 14092 2624
rect 14092 2575 14132 2584
rect 14284 2624 14324 2659
rect 14188 2540 14228 2549
rect 13900 2500 14036 2540
rect 13803 2456 13845 2465
rect 13803 2416 13804 2456
rect 13844 2416 13845 2456
rect 13803 2407 13845 2416
rect 13900 1121 13940 1206
rect 13324 80 13364 895
rect 13420 533 13460 904
rect 13516 904 13652 944
rect 13708 1112 13748 1121
rect 13419 524 13461 533
rect 13419 484 13420 524
rect 13460 484 13461 524
rect 13419 475 13461 484
rect 13516 80 13556 904
rect 13708 785 13748 1072
rect 13899 1112 13941 1121
rect 13899 1072 13900 1112
rect 13940 1072 13941 1112
rect 13899 1063 13941 1072
rect 13803 944 13845 953
rect 13996 944 14036 2500
rect 14092 1205 14132 1207
rect 14091 1196 14133 1205
rect 14091 1156 14092 1196
rect 14132 1156 14133 1196
rect 14091 1147 14133 1156
rect 14092 1112 14132 1147
rect 14092 1063 14132 1072
rect 13803 904 13804 944
rect 13844 904 13845 944
rect 13803 895 13845 904
rect 13900 904 14036 944
rect 14091 944 14133 953
rect 14091 904 14092 944
rect 14132 904 14133 944
rect 13804 810 13844 895
rect 13707 776 13749 785
rect 13707 736 13708 776
rect 13748 736 13749 776
rect 13707 727 13749 736
rect 13707 524 13749 533
rect 13707 484 13708 524
rect 13748 484 13749 524
rect 13707 475 13749 484
rect 13708 80 13748 475
rect 13900 80 13940 904
rect 14091 895 14133 904
rect 14092 80 14132 895
rect 14188 776 14228 2500
rect 14284 2381 14324 2584
rect 14380 2540 14420 3172
rect 14476 2717 14516 3424
rect 14668 3464 14708 3499
rect 14668 3413 14708 3424
rect 14860 3464 14900 3473
rect 14764 3212 14804 3221
rect 14475 2708 14517 2717
rect 14475 2668 14476 2708
rect 14516 2668 14517 2708
rect 14475 2659 14517 2668
rect 14764 2540 14804 3172
rect 14860 2801 14900 3424
rect 15052 3464 15092 3499
rect 15052 3413 15092 3424
rect 15244 3464 15284 3583
rect 15435 3548 15477 3557
rect 15435 3508 15436 3548
rect 15476 3508 15477 3548
rect 15435 3499 15477 3508
rect 15819 3548 15861 3557
rect 15819 3508 15820 3548
rect 15860 3508 15861 3548
rect 15819 3499 15861 3508
rect 16203 3548 16245 3557
rect 16203 3508 16204 3548
rect 16244 3508 16245 3548
rect 16203 3499 16245 3508
rect 16587 3548 16629 3557
rect 16587 3508 16588 3548
rect 16628 3508 16629 3548
rect 16587 3499 16629 3508
rect 15244 3415 15284 3424
rect 15436 3464 15476 3499
rect 15436 3413 15476 3424
rect 15628 3464 15668 3473
rect 15628 3296 15668 3424
rect 15820 3464 15860 3499
rect 15820 3413 15860 3424
rect 16011 3464 16053 3473
rect 16011 3424 16012 3464
rect 16052 3424 16053 3464
rect 16011 3415 16053 3424
rect 16204 3464 16244 3499
rect 16012 3330 16052 3415
rect 16204 3413 16244 3424
rect 16396 3464 16436 3473
rect 15819 3296 15861 3305
rect 15628 3256 15820 3296
rect 15860 3256 15861 3296
rect 15819 3247 15861 3256
rect 15148 3212 15188 3221
rect 14859 2792 14901 2801
rect 14859 2752 14860 2792
rect 14900 2752 14901 2792
rect 14859 2743 14901 2752
rect 15148 2540 15188 3172
rect 15532 3212 15572 3221
rect 15916 3212 15956 3221
rect 16300 3212 16340 3221
rect 15572 3172 15764 3212
rect 15532 3163 15572 3172
rect 15724 2540 15764 3172
rect 15956 3172 16244 3212
rect 15916 3163 15956 3172
rect 14380 2500 14612 2540
rect 14764 2500 14996 2540
rect 15148 2500 15572 2540
rect 15724 2500 15956 2540
rect 14283 2372 14325 2381
rect 14283 2332 14284 2372
rect 14324 2332 14325 2372
rect 14283 2323 14325 2332
rect 14283 1364 14325 1373
rect 14283 1324 14284 1364
rect 14324 1324 14325 1364
rect 14572 1364 14612 2500
rect 14956 1364 14996 2500
rect 14572 1324 14804 1364
rect 14956 1324 15188 1364
rect 14283 1315 14325 1324
rect 14284 1230 14324 1315
rect 14668 1121 14708 1206
rect 14283 1112 14325 1121
rect 14476 1112 14516 1121
rect 14283 1072 14284 1112
rect 14324 1072 14325 1112
rect 14283 1063 14325 1072
rect 14380 1072 14476 1112
rect 14284 978 14324 1063
rect 14380 869 14420 1072
rect 14476 1063 14516 1072
rect 14667 1112 14709 1121
rect 14667 1072 14668 1112
rect 14708 1072 14709 1112
rect 14667 1063 14709 1072
rect 14572 953 14612 1038
rect 14571 944 14613 953
rect 14764 944 14804 1324
rect 14859 1196 14901 1205
rect 14859 1156 14860 1196
rect 14900 1156 14901 1196
rect 14859 1147 14901 1156
rect 15051 1196 15093 1205
rect 15051 1156 15052 1196
rect 15092 1156 15093 1196
rect 15051 1147 15093 1156
rect 14860 1112 14900 1147
rect 14860 1061 14900 1072
rect 15052 1112 15092 1147
rect 15052 1061 15092 1072
rect 14571 904 14572 944
rect 14612 904 14613 944
rect 14571 895 14613 904
rect 14668 904 14804 944
rect 14859 944 14901 953
rect 14859 904 14860 944
rect 14900 904 14901 944
rect 14379 860 14421 869
rect 14379 820 14380 860
rect 14420 820 14421 860
rect 14379 811 14421 820
rect 14571 776 14613 785
rect 14188 736 14324 776
rect 14284 80 14324 736
rect 14571 736 14572 776
rect 14612 736 14613 776
rect 14571 727 14613 736
rect 14475 692 14517 701
rect 14475 652 14476 692
rect 14516 652 14517 692
rect 14475 643 14517 652
rect 14476 80 14516 643
rect 14572 281 14612 727
rect 14571 272 14613 281
rect 14571 232 14572 272
rect 14612 232 14613 272
rect 14571 223 14613 232
rect 14668 80 14708 904
rect 14859 895 14901 904
rect 14956 944 14996 953
rect 15148 944 15188 1324
rect 15243 1280 15285 1289
rect 15243 1240 15244 1280
rect 15284 1240 15285 1280
rect 15243 1231 15285 1240
rect 14860 80 14900 895
rect 14956 281 14996 904
rect 15052 904 15188 944
rect 15244 1112 15284 1231
rect 15435 1196 15477 1205
rect 15435 1156 15436 1196
rect 15476 1156 15477 1196
rect 15435 1147 15477 1156
rect 14955 272 14997 281
rect 14955 232 14956 272
rect 14996 232 14997 272
rect 14955 223 14997 232
rect 15052 80 15092 904
rect 15244 701 15284 1072
rect 15436 1112 15476 1147
rect 15436 1061 15476 1072
rect 15340 944 15380 953
rect 15243 692 15285 701
rect 15243 652 15244 692
rect 15284 652 15285 692
rect 15243 643 15285 652
rect 15340 281 15380 904
rect 15532 860 15572 2500
rect 15819 1196 15861 1205
rect 15819 1156 15820 1196
rect 15860 1156 15861 1196
rect 15819 1147 15861 1156
rect 15628 1112 15668 1123
rect 15628 1037 15668 1072
rect 15820 1112 15860 1147
rect 15820 1061 15860 1072
rect 15627 1028 15669 1037
rect 15627 988 15628 1028
rect 15668 988 15669 1028
rect 15627 979 15669 988
rect 15723 944 15765 953
rect 15916 944 15956 2500
rect 16204 1364 16244 3172
rect 16300 1448 16340 3172
rect 16396 2885 16436 3424
rect 16588 3464 16628 3499
rect 16588 3413 16628 3424
rect 16780 3464 16820 3667
rect 16971 3548 17013 3557
rect 16971 3508 16972 3548
rect 17012 3508 17013 3548
rect 16971 3499 17013 3508
rect 17355 3548 17397 3557
rect 17355 3508 17356 3548
rect 17396 3508 17397 3548
rect 17355 3499 17397 3508
rect 17931 3548 17973 3557
rect 17931 3508 17932 3548
rect 17972 3508 17973 3548
rect 17931 3499 17973 3508
rect 16780 3305 16820 3424
rect 16972 3464 17012 3499
rect 16972 3413 17012 3424
rect 17163 3464 17205 3473
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 17356 3464 17396 3499
rect 17164 3330 17204 3415
rect 17356 3413 17396 3424
rect 17547 3464 17589 3473
rect 17547 3424 17548 3464
rect 17588 3424 17589 3464
rect 17547 3415 17589 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 17932 3464 17972 3499
rect 18124 3473 18164 4012
rect 18316 4002 18356 4087
rect 18411 3968 18453 3977
rect 18411 3928 18412 3968
rect 18452 3928 18453 3968
rect 18411 3919 18453 3928
rect 18412 3834 18452 3919
rect 18508 3893 18548 4096
rect 18796 4052 18836 4061
rect 18507 3884 18549 3893
rect 18507 3844 18508 3884
rect 18548 3844 18549 3884
rect 18507 3835 18549 3844
rect 18796 3809 18836 4012
rect 18892 3977 18932 4507
rect 19083 4388 19125 4397
rect 19083 4348 19084 4388
rect 19124 4348 19125 4388
rect 19083 4339 19125 4348
rect 19084 4167 19124 4339
rect 18988 4136 19028 4147
rect 19084 4118 19124 4127
rect 19468 4136 19508 4507
rect 19755 4388 19797 4397
rect 19755 4348 19756 4388
rect 19796 4348 19797 4388
rect 19755 4339 19797 4348
rect 19756 4145 19796 4339
rect 18988 4061 19028 4096
rect 19468 4087 19508 4096
rect 19660 4136 19700 4145
rect 18987 4052 19029 4061
rect 18987 4012 18988 4052
rect 19028 4012 19029 4052
rect 18987 4003 19029 4012
rect 19084 3977 19124 4062
rect 19179 4052 19221 4061
rect 19179 4012 19180 4052
rect 19220 4012 19221 4052
rect 19179 4003 19221 4012
rect 18891 3968 18933 3977
rect 18891 3928 18892 3968
rect 18932 3928 18933 3968
rect 18891 3919 18933 3928
rect 19083 3968 19125 3977
rect 19083 3928 19084 3968
rect 19124 3928 19125 3968
rect 19083 3919 19125 3928
rect 18795 3800 18837 3809
rect 18795 3760 18796 3800
rect 18836 3760 18837 3800
rect 18795 3751 18837 3760
rect 17548 3330 17588 3415
rect 17740 3330 17780 3415
rect 16779 3296 16821 3305
rect 16779 3256 16780 3296
rect 16820 3256 16821 3296
rect 16779 3247 16821 3256
rect 17932 3221 17972 3424
rect 18123 3464 18165 3473
rect 18123 3424 18124 3464
rect 18164 3424 18165 3464
rect 18123 3415 18165 3424
rect 18316 3464 18356 3473
rect 18124 3330 18164 3415
rect 18316 3221 18356 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18699 3464 18741 3473
rect 18699 3424 18700 3464
rect 18740 3424 18741 3464
rect 18699 3415 18741 3424
rect 18892 3464 18932 3919
rect 19083 3800 19125 3809
rect 19083 3760 19084 3800
rect 19124 3760 19125 3800
rect 19083 3751 19125 3760
rect 18892 3415 18932 3424
rect 19084 3464 19124 3751
rect 19084 3415 19124 3424
rect 19180 3464 19220 4003
rect 19660 3977 19700 4096
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 19756 4002 19796 4087
rect 19948 3977 19988 4087
rect 19468 3968 19508 3977
rect 19180 3415 19220 3424
rect 19276 3928 19468 3968
rect 18508 3330 18548 3415
rect 18700 3330 18740 3415
rect 16684 3212 16724 3221
rect 16395 2876 16437 2885
rect 16395 2836 16396 2876
rect 16436 2836 16437 2876
rect 16395 2827 16437 2836
rect 16684 2540 16724 3172
rect 17068 3212 17108 3221
rect 17452 3212 17492 3221
rect 17836 3212 17876 3221
rect 17108 3172 17300 3212
rect 17068 3163 17108 3172
rect 17260 2540 17300 3172
rect 17492 3172 17588 3212
rect 17452 3163 17492 3172
rect 16684 2500 17108 2540
rect 17260 2500 17492 2540
rect 16300 1408 16532 1448
rect 16204 1324 16340 1364
rect 16012 1121 16052 1206
rect 16203 1196 16245 1205
rect 16203 1156 16204 1196
rect 16244 1156 16245 1196
rect 16203 1147 16245 1156
rect 16011 1112 16053 1121
rect 16011 1072 16012 1112
rect 16052 1072 16053 1112
rect 16011 1063 16053 1072
rect 16204 1112 16244 1147
rect 16204 1061 16244 1072
rect 15723 904 15724 944
rect 15764 904 15765 944
rect 15723 895 15765 904
rect 15820 904 15956 944
rect 16011 944 16053 953
rect 16011 904 16012 944
rect 16052 904 16053 944
rect 15436 820 15572 860
rect 15147 272 15189 281
rect 15339 272 15381 281
rect 15147 232 15148 272
rect 15188 232 15284 272
rect 15147 223 15189 232
rect 15244 80 15284 232
rect 15339 232 15340 272
rect 15380 232 15381 272
rect 15339 223 15381 232
rect 15436 80 15476 820
rect 15724 810 15764 895
rect 15627 272 15669 281
rect 15627 232 15628 272
rect 15668 232 15669 272
rect 15627 223 15669 232
rect 15628 80 15668 223
rect 15820 80 15860 904
rect 16011 895 16053 904
rect 16108 944 16148 953
rect 16300 944 16340 1324
rect 16395 1280 16437 1289
rect 16395 1240 16396 1280
rect 16436 1240 16437 1280
rect 16395 1231 16437 1240
rect 16396 1112 16436 1231
rect 16396 1037 16436 1072
rect 16395 1028 16437 1037
rect 16395 988 16396 1028
rect 16436 988 16437 1028
rect 16395 979 16437 988
rect 16012 80 16052 895
rect 16108 281 16148 904
rect 16204 904 16340 944
rect 16492 944 16532 1408
rect 16588 1364 16628 1373
rect 16628 1324 16724 1364
rect 16588 1315 16628 1324
rect 16588 1205 16628 1220
rect 16587 1196 16629 1205
rect 16587 1156 16588 1196
rect 16628 1156 16629 1196
rect 16587 1147 16629 1156
rect 16588 1125 16628 1147
rect 16588 1076 16628 1085
rect 16684 1028 16724 1324
rect 16779 1280 16821 1289
rect 16779 1240 16780 1280
rect 16820 1240 16821 1280
rect 16779 1231 16821 1240
rect 16780 1125 16820 1231
rect 16971 1196 17013 1205
rect 16971 1156 16972 1196
rect 17012 1156 17013 1196
rect 16971 1147 17013 1156
rect 16780 1076 16820 1085
rect 16972 1112 17012 1147
rect 16972 1061 17012 1072
rect 16684 988 16820 1028
rect 16492 904 16628 944
rect 16107 272 16149 281
rect 16107 232 16108 272
rect 16148 232 16149 272
rect 16107 223 16149 232
rect 16204 80 16244 904
rect 16395 272 16437 281
rect 16395 232 16396 272
rect 16436 232 16437 272
rect 16395 223 16437 232
rect 16396 80 16436 223
rect 16588 80 16628 904
rect 16683 860 16725 869
rect 16683 820 16684 860
rect 16724 820 16725 860
rect 16683 811 16725 820
rect 16684 281 16724 811
rect 16683 272 16725 281
rect 16683 232 16684 272
rect 16724 232 16725 272
rect 16683 223 16725 232
rect 16780 80 16820 988
rect 16875 944 16917 953
rect 17068 944 17108 2500
rect 17164 1121 17204 1206
rect 17355 1196 17397 1205
rect 17355 1156 17356 1196
rect 17396 1156 17397 1196
rect 17355 1147 17397 1156
rect 17163 1112 17205 1121
rect 17163 1072 17164 1112
rect 17204 1072 17205 1112
rect 17163 1063 17205 1072
rect 17356 1112 17396 1147
rect 17356 1061 17396 1072
rect 16875 904 16876 944
rect 16916 904 16917 944
rect 16875 895 16917 904
rect 16972 904 17108 944
rect 17163 944 17205 953
rect 17163 904 17164 944
rect 17204 904 17205 944
rect 16876 810 16916 895
rect 16972 80 17012 904
rect 17163 895 17205 904
rect 17260 944 17300 953
rect 17452 944 17492 2500
rect 17548 1280 17588 3172
rect 17836 2540 17876 3172
rect 17931 3212 17973 3221
rect 18220 3212 18260 3221
rect 17931 3172 17932 3212
rect 17972 3172 17973 3212
rect 17931 3163 17973 3172
rect 18124 3172 18220 3212
rect 18124 2876 18164 3172
rect 18220 3163 18260 3172
rect 18315 3212 18357 3221
rect 18315 3172 18316 3212
rect 18356 3172 18357 3212
rect 18315 3163 18357 3172
rect 18604 3212 18644 3221
rect 18892 3212 18932 3221
rect 18644 3172 18836 3212
rect 18604 3163 18644 3172
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 18124 2836 18740 2876
rect 17836 2500 18164 2540
rect 18124 1364 18164 2500
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 18124 1324 18260 1364
rect 17548 1240 17684 1280
rect 17644 1121 17684 1240
rect 17548 1112 17588 1121
rect 17548 953 17588 1072
rect 17643 1112 17685 1121
rect 17643 1072 17644 1112
rect 17684 1072 17685 1112
rect 17643 1063 17685 1072
rect 17740 1112 17780 1121
rect 17835 1112 17877 1121
rect 17780 1072 17836 1112
rect 17876 1072 17877 1112
rect 17740 1063 17780 1072
rect 17835 1063 17877 1072
rect 17932 1112 17972 1123
rect 17932 1037 17972 1072
rect 18027 1112 18069 1121
rect 18114 1112 18154 1118
rect 18027 1072 18028 1112
rect 18068 1109 18154 1112
rect 18068 1072 18114 1109
rect 18027 1063 18069 1072
rect 18114 1060 18154 1069
rect 17931 1028 17973 1037
rect 17931 988 17932 1028
rect 17972 988 17973 1028
rect 17931 979 17973 988
rect 17164 80 17204 895
rect 17260 533 17300 904
rect 17356 904 17492 944
rect 17547 944 17589 953
rect 17547 904 17548 944
rect 17588 904 17589 944
rect 17259 524 17301 533
rect 17259 484 17260 524
rect 17300 484 17301 524
rect 17259 475 17301 484
rect 17356 80 17396 904
rect 17547 895 17589 904
rect 17644 944 17684 953
rect 17739 944 17781 953
rect 17684 904 17740 944
rect 17780 904 17781 944
rect 17644 895 17684 904
rect 17739 895 17781 904
rect 18027 944 18069 953
rect 18220 944 18260 1324
rect 18700 1280 18740 2836
rect 18796 1364 18836 3172
rect 18892 1625 18932 3172
rect 18987 3128 19029 3137
rect 18987 3088 18988 3128
rect 19028 3088 19029 3128
rect 18987 3079 19029 3088
rect 18988 2801 19028 3079
rect 18987 2792 19029 2801
rect 18987 2752 18988 2792
rect 19028 2752 19029 2792
rect 18987 2743 19029 2752
rect 19276 2540 19316 3928
rect 19468 3919 19508 3928
rect 19659 3968 19701 3977
rect 19659 3928 19660 3968
rect 19700 3928 19701 3968
rect 19659 3919 19701 3928
rect 19947 3968 19989 3977
rect 19947 3928 19948 3968
rect 19988 3928 19989 3968
rect 20044 3968 20084 4507
rect 22348 4229 22388 4684
rect 22347 4220 22389 4229
rect 22347 4180 22348 4220
rect 22388 4180 22389 4220
rect 22347 4171 22389 4180
rect 22444 4061 22484 4936
rect 41164 4724 41204 4733
rect 40972 4684 41164 4724
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 38667 4556 38709 4565
rect 38667 4516 38668 4556
rect 38708 4516 38709 4556
rect 38667 4507 38709 4516
rect 37323 4388 37365 4397
rect 37323 4348 37324 4388
rect 37364 4348 37365 4388
rect 37323 4339 37365 4348
rect 38187 4388 38229 4397
rect 38187 4348 38188 4388
rect 38228 4348 38229 4388
rect 38187 4339 38229 4348
rect 38668 4388 38708 4507
rect 38955 4472 38997 4481
rect 38955 4432 38956 4472
rect 38996 4432 38997 4472
rect 38955 4423 38997 4432
rect 38668 4339 38708 4348
rect 25899 4304 25941 4313
rect 25899 4264 25900 4304
rect 25940 4264 25941 4304
rect 25899 4255 25941 4264
rect 28011 4304 28053 4313
rect 28011 4264 28012 4304
rect 28052 4264 28053 4304
rect 28011 4255 28053 4264
rect 24459 4220 24501 4229
rect 24268 4180 24404 4220
rect 24268 4061 24308 4180
rect 24364 4136 24404 4180
rect 24459 4180 24460 4220
rect 24500 4180 24501 4220
rect 24459 4171 24501 4180
rect 25131 4220 25173 4229
rect 25131 4180 25132 4220
rect 25172 4180 25173 4220
rect 25131 4171 25173 4180
rect 24364 4087 24404 4096
rect 24460 4136 24500 4171
rect 24460 4085 24500 4096
rect 24844 4136 24884 4145
rect 25036 4136 25076 4147
rect 24884 4096 24980 4136
rect 24844 4087 24884 4096
rect 22443 4052 22485 4061
rect 22443 4012 22444 4052
rect 22484 4012 22485 4052
rect 22443 4003 22485 4012
rect 24267 4052 24309 4061
rect 24267 4012 24268 4052
rect 24308 4012 24309 4052
rect 24267 4003 24309 4012
rect 24652 4052 24692 4061
rect 20235 3968 20277 3977
rect 20044 3928 20236 3968
rect 20276 3928 20277 3968
rect 19947 3919 19989 3928
rect 20235 3919 20277 3928
rect 24363 3968 24405 3977
rect 24363 3928 24364 3968
rect 24404 3928 24405 3968
rect 24363 3919 24405 3928
rect 24364 3834 24404 3919
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 21099 3800 21141 3809
rect 21099 3760 21100 3800
rect 21140 3760 21141 3800
rect 21099 3751 21141 3760
rect 19371 3548 19413 3557
rect 19371 3508 19372 3548
rect 19412 3508 19413 3548
rect 19371 3499 19413 3508
rect 19372 3221 19412 3499
rect 20149 3473 20189 3573
rect 20715 3548 20757 3557
rect 20715 3508 20716 3548
rect 20756 3508 20757 3548
rect 20715 3499 20757 3508
rect 19947 3464 19989 3473
rect 19947 3424 19948 3464
rect 19988 3424 19989 3464
rect 19947 3415 19989 3424
rect 20148 3464 20190 3473
rect 20148 3415 20149 3464
rect 19948 3330 19988 3415
rect 20189 3415 20190 3464
rect 20716 3464 20756 3499
rect 19371 3212 19413 3221
rect 19371 3172 19372 3212
rect 19412 3172 19413 3212
rect 19371 3163 19413 3172
rect 20044 3212 20084 3221
rect 20149 3212 20189 3409
rect 20149 3172 20276 3212
rect 20044 2885 20084 3172
rect 20043 2876 20085 2885
rect 20043 2836 20044 2876
rect 20084 2836 20085 2876
rect 20043 2827 20085 2836
rect 19851 2792 19893 2801
rect 19851 2752 19852 2792
rect 19892 2752 19893 2792
rect 19851 2743 19893 2752
rect 19660 2633 19700 2718
rect 19467 2624 19509 2633
rect 19467 2584 19468 2624
rect 19508 2584 19509 2624
rect 19467 2575 19509 2584
rect 19659 2624 19701 2633
rect 19659 2584 19660 2624
rect 19700 2584 19701 2624
rect 19659 2575 19701 2584
rect 19852 2624 19892 2743
rect 20236 2633 20276 3172
rect 20428 2633 20468 2718
rect 20716 2717 20756 3424
rect 20907 3464 20949 3473
rect 20907 3424 20908 3464
rect 20948 3424 20949 3464
rect 20907 3415 20949 3424
rect 21100 3464 21140 3751
rect 21675 3716 21717 3725
rect 21580 3676 21676 3716
rect 21716 3676 21717 3716
rect 21387 3632 21429 3641
rect 21387 3592 21388 3632
rect 21428 3592 21524 3632
rect 21387 3583 21429 3592
rect 20908 3330 20948 3415
rect 20812 3212 20852 3221
rect 20715 2708 20757 2717
rect 20715 2668 20716 2708
rect 20756 2668 20757 2708
rect 20715 2659 20757 2668
rect 19180 2500 19316 2540
rect 18891 1616 18933 1625
rect 18891 1576 18892 1616
rect 18932 1576 18933 1616
rect 18891 1567 18933 1576
rect 18796 1324 19028 1364
rect 18604 1240 18740 1280
rect 18316 1205 18356 1207
rect 18315 1196 18357 1205
rect 18315 1156 18316 1196
rect 18356 1156 18357 1196
rect 18315 1147 18357 1156
rect 18316 1112 18356 1147
rect 18316 1063 18356 1072
rect 18507 1112 18549 1121
rect 18507 1072 18508 1112
rect 18548 1072 18549 1112
rect 18507 1063 18549 1072
rect 18508 978 18548 1063
rect 18027 904 18028 944
rect 18068 904 18069 944
rect 18027 895 18069 904
rect 18124 904 18260 944
rect 18315 944 18357 953
rect 18315 904 18316 944
rect 18356 904 18357 944
rect 17931 860 17973 869
rect 17931 820 17932 860
rect 17972 820 17973 860
rect 17931 811 17973 820
rect 17739 776 17781 785
rect 17739 736 17740 776
rect 17780 736 17781 776
rect 17739 727 17781 736
rect 17547 524 17589 533
rect 17547 484 17548 524
rect 17588 484 17589 524
rect 17547 475 17589 484
rect 17548 80 17588 475
rect 17740 80 17780 727
rect 17932 80 17972 811
rect 18028 810 18068 895
rect 18124 80 18164 904
rect 18315 895 18357 904
rect 18412 944 18452 953
rect 18316 80 18356 895
rect 18412 533 18452 904
rect 18604 860 18644 1240
rect 18700 1112 18740 1123
rect 18700 1037 18740 1072
rect 18891 1112 18933 1121
rect 18891 1072 18892 1112
rect 18932 1072 18933 1112
rect 18891 1063 18933 1072
rect 18699 1028 18741 1037
rect 18699 988 18700 1028
rect 18740 988 18741 1028
rect 18699 979 18741 988
rect 18892 978 18932 1063
rect 18795 944 18837 953
rect 18795 904 18796 944
rect 18836 904 18837 944
rect 18795 895 18837 904
rect 18508 820 18644 860
rect 18699 860 18741 869
rect 18699 820 18700 860
rect 18740 820 18741 860
rect 18411 524 18453 533
rect 18411 484 18412 524
rect 18452 484 18453 524
rect 18411 475 18453 484
rect 18508 80 18548 820
rect 18699 811 18741 820
rect 18700 692 18740 811
rect 18796 810 18836 895
rect 18988 860 19028 1324
rect 19083 1280 19125 1289
rect 19083 1240 19084 1280
rect 19124 1240 19125 1280
rect 19083 1231 19125 1240
rect 19084 1112 19124 1231
rect 19180 1121 19220 2500
rect 19468 2456 19508 2575
rect 19372 2416 19508 2456
rect 19756 2540 19796 2549
rect 19852 2540 19892 2584
rect 20235 2624 20277 2633
rect 20235 2584 20236 2624
rect 20276 2584 20277 2624
rect 20235 2575 20277 2584
rect 20427 2624 20469 2633
rect 20427 2584 20428 2624
rect 20468 2584 20469 2624
rect 20427 2575 20469 2584
rect 20332 2540 20372 2549
rect 19852 2500 20084 2540
rect 19756 2456 19796 2500
rect 19756 2416 19988 2456
rect 19372 2297 19412 2416
rect 19371 2288 19413 2297
rect 19371 2248 19372 2288
rect 19412 2248 19413 2288
rect 19371 2239 19413 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 19371 1952 19413 1961
rect 19371 1912 19372 1952
rect 19412 1912 19413 1952
rect 19371 1903 19413 1912
rect 19563 1952 19605 1961
rect 19563 1912 19564 1952
rect 19604 1912 19605 1952
rect 19563 1903 19605 1912
rect 19372 1818 19412 1903
rect 19564 1818 19604 1903
rect 19468 1700 19508 1709
rect 19372 1660 19468 1700
rect 19276 1205 19316 1220
rect 19275 1196 19317 1205
rect 19275 1156 19276 1196
rect 19316 1156 19317 1196
rect 19275 1147 19317 1156
rect 19276 1125 19316 1147
rect 19084 1063 19124 1072
rect 19179 1112 19221 1121
rect 19179 1072 19180 1112
rect 19220 1072 19221 1112
rect 19276 1076 19316 1085
rect 19179 1063 19221 1072
rect 19083 944 19125 953
rect 19083 904 19084 944
rect 19124 904 19125 944
rect 19083 895 19125 904
rect 19180 944 19220 953
rect 18892 820 19028 860
rect 18700 652 18836 692
rect 18699 524 18741 533
rect 18699 484 18700 524
rect 18740 484 18741 524
rect 18699 475 18741 484
rect 18700 80 18740 475
rect 18796 449 18836 652
rect 18795 440 18837 449
rect 18795 400 18796 440
rect 18836 400 18837 440
rect 18795 391 18837 400
rect 18892 80 18932 820
rect 19084 80 19124 895
rect 19180 533 19220 904
rect 19372 860 19412 1660
rect 19468 1651 19508 1660
rect 19467 1448 19509 1457
rect 19467 1408 19468 1448
rect 19508 1408 19509 1448
rect 19467 1399 19509 1408
rect 19468 1289 19508 1399
rect 19467 1280 19509 1289
rect 19467 1240 19468 1280
rect 19508 1240 19509 1280
rect 19467 1231 19509 1240
rect 19851 1280 19893 1289
rect 19851 1240 19852 1280
rect 19892 1240 19893 1280
rect 19851 1231 19893 1240
rect 19468 1112 19508 1231
rect 19660 1121 19700 1206
rect 19468 1063 19508 1072
rect 19659 1112 19701 1121
rect 19659 1072 19660 1112
rect 19700 1072 19701 1112
rect 19659 1063 19701 1072
rect 19852 1112 19892 1231
rect 19948 1205 19988 2416
rect 20044 1961 20084 2500
rect 20812 2540 20852 3172
rect 21100 3137 21140 3424
rect 21291 3464 21333 3473
rect 21291 3424 21292 3464
rect 21332 3424 21333 3464
rect 21291 3415 21333 3424
rect 21484 3464 21524 3592
rect 21580 3464 21620 3676
rect 21675 3667 21717 3676
rect 23115 3632 23157 3641
rect 23115 3592 23116 3632
rect 23156 3592 23157 3632
rect 23115 3583 23157 3592
rect 21524 3424 21620 3464
rect 21675 3464 21717 3473
rect 21675 3424 21676 3464
rect 21716 3424 21717 3464
rect 21484 3415 21524 3424
rect 21675 3415 21717 3424
rect 22059 3464 22101 3473
rect 22156 3464 22196 3492
rect 22059 3424 22060 3464
rect 22100 3424 22156 3464
rect 22059 3415 22101 3424
rect 22156 3415 22196 3424
rect 22348 3464 22388 3475
rect 21292 3330 21332 3415
rect 21676 3330 21716 3415
rect 21196 3212 21236 3221
rect 21099 3128 21141 3137
rect 21099 3088 21100 3128
rect 21140 3088 21141 3128
rect 21099 3079 21141 3088
rect 21196 2540 21236 3172
rect 21580 3212 21620 3221
rect 21580 2540 21620 3172
rect 21868 2633 21908 2718
rect 21867 2624 21909 2633
rect 21867 2584 21868 2624
rect 21908 2584 21909 2624
rect 21867 2575 21909 2584
rect 22060 2624 22100 3415
rect 22348 3389 22388 3424
rect 22539 3464 22581 3473
rect 22539 3424 22540 3464
rect 22580 3424 22581 3464
rect 22539 3415 22581 3424
rect 22732 3464 22772 3473
rect 22347 3380 22389 3389
rect 22347 3340 22348 3380
rect 22388 3340 22389 3380
rect 22347 3331 22389 3340
rect 22540 3330 22580 3415
rect 22060 2575 22100 2584
rect 22252 3212 22292 3221
rect 21964 2540 22004 2549
rect 20812 2500 20948 2540
rect 21196 2500 21332 2540
rect 21580 2500 21716 2540
rect 20043 1952 20085 1961
rect 20043 1912 20044 1952
rect 20084 1912 20085 1952
rect 20043 1903 20085 1912
rect 20236 1205 20276 1207
rect 19947 1196 19989 1205
rect 19947 1156 19948 1196
rect 19988 1156 19989 1196
rect 19947 1147 19989 1156
rect 20235 1196 20277 1205
rect 20235 1156 20236 1196
rect 20276 1156 20277 1196
rect 20235 1147 20277 1156
rect 19564 953 19604 1038
rect 19852 1037 19892 1072
rect 20043 1112 20085 1121
rect 20043 1072 20044 1112
rect 20084 1072 20085 1112
rect 20043 1063 20085 1072
rect 20236 1112 20276 1147
rect 20236 1063 20276 1072
rect 19851 1028 19893 1037
rect 19851 988 19852 1028
rect 19892 988 19893 1028
rect 19851 979 19893 988
rect 20044 978 20084 1063
rect 19563 944 19605 953
rect 19563 904 19564 944
rect 19604 904 19605 944
rect 19563 895 19605 904
rect 19947 944 19989 953
rect 19947 904 19948 944
rect 19988 904 19989 944
rect 19947 895 19989 904
rect 20235 944 20277 953
rect 20235 904 20236 944
rect 20276 904 20277 944
rect 20235 895 20277 904
rect 19276 820 19412 860
rect 19276 692 19316 820
rect 19948 810 19988 895
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 19275 652 19316 692
rect 19275 608 19315 652
rect 19275 568 19316 608
rect 19179 524 19221 533
rect 19276 524 19316 568
rect 19179 484 19180 524
rect 19220 484 19221 524
rect 19179 475 19221 484
rect 19275 484 19316 524
rect 19467 524 19509 533
rect 19947 524 19989 533
rect 19467 484 19468 524
rect 19508 484 19511 524
rect 19275 440 19315 484
rect 19467 475 19511 484
rect 19947 484 19948 524
rect 19988 484 19989 524
rect 19947 475 19989 484
rect 19275 400 19412 440
rect 19372 356 19412 400
rect 19471 356 19511 475
rect 19948 356 19988 475
rect 19369 316 19412 356
rect 19468 316 19511 356
rect 19659 316 19988 356
rect 19369 272 19409 316
rect 19283 232 19409 272
rect 19283 104 19323 232
rect 19276 80 19323 104
rect 19468 80 19508 316
rect 19659 188 19699 316
rect 19659 148 19700 188
rect 19660 80 19700 148
rect 19851 104 19893 113
rect 19851 80 19852 104
rect 824 0 904 80
rect 1016 0 1096 80
rect 1208 0 1288 80
rect 1400 0 1480 80
rect 1592 0 1672 80
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 64 19852 80
rect 19892 80 19893 104
rect 20043 104 20085 113
rect 20043 80 20044 104
rect 19892 64 19912 80
rect 19832 0 19912 64
rect 20024 64 20044 80
rect 20084 80 20085 104
rect 20236 80 20276 895
rect 20332 776 20372 2500
rect 20427 1532 20469 1541
rect 20427 1492 20428 1532
rect 20468 1492 20469 1532
rect 20427 1483 20469 1492
rect 20428 1364 20468 1483
rect 20428 1315 20468 1324
rect 20812 1121 20852 1206
rect 20427 1112 20469 1121
rect 20427 1072 20428 1112
rect 20468 1072 20469 1112
rect 20811 1112 20853 1121
rect 20427 1063 20469 1072
rect 20620 1101 20660 1110
rect 20428 978 20468 1063
rect 20811 1072 20812 1112
rect 20852 1072 20853 1112
rect 20811 1063 20853 1072
rect 20620 1037 20660 1061
rect 20619 1028 20661 1037
rect 20619 988 20620 1028
rect 20660 988 20661 1028
rect 20619 979 20661 988
rect 20620 966 20660 979
rect 20715 944 20757 953
rect 20908 944 20948 2500
rect 21004 1205 21044 1207
rect 21003 1196 21045 1205
rect 21003 1156 21004 1196
rect 21044 1156 21045 1196
rect 21003 1147 21045 1156
rect 21195 1196 21237 1205
rect 21195 1156 21196 1196
rect 21236 1156 21237 1196
rect 21195 1147 21237 1156
rect 21004 1112 21044 1147
rect 21004 1063 21044 1072
rect 21196 1112 21236 1147
rect 21196 1061 21236 1072
rect 20715 904 20716 944
rect 20756 904 20757 944
rect 20715 895 20757 904
rect 20812 904 20948 944
rect 21003 944 21045 953
rect 21003 904 21004 944
rect 21044 904 21045 944
rect 20716 810 20756 895
rect 20332 736 20468 776
rect 20428 80 20468 736
rect 20619 524 20661 533
rect 20619 484 20620 524
rect 20660 484 20661 524
rect 20619 475 20661 484
rect 20620 80 20660 475
rect 20812 80 20852 904
rect 21003 895 21045 904
rect 21100 944 21140 953
rect 21292 944 21332 2500
rect 21580 1205 21620 1220
rect 21579 1196 21621 1205
rect 21579 1156 21580 1196
rect 21620 1156 21621 1196
rect 21579 1147 21621 1156
rect 21580 1125 21620 1147
rect 21004 80 21044 895
rect 21100 533 21140 904
rect 21196 904 21332 944
rect 21388 1112 21428 1121
rect 21580 1076 21620 1085
rect 21099 524 21141 533
rect 21099 484 21100 524
rect 21140 484 21141 524
rect 21099 475 21141 484
rect 21196 80 21236 904
rect 21388 869 21428 1072
rect 21676 1028 21716 2500
rect 22252 2540 22292 3172
rect 22636 3212 22676 3221
rect 22636 2792 22676 3172
rect 22732 2969 22772 3424
rect 22923 3464 22965 3473
rect 22923 3424 22924 3464
rect 22964 3424 22965 3464
rect 22923 3415 22965 3424
rect 23116 3464 23156 3583
rect 22924 3330 22964 3415
rect 23020 3212 23060 3221
rect 22731 2960 22773 2969
rect 22731 2920 22732 2960
rect 22772 2920 22773 2960
rect 22731 2911 22773 2920
rect 22636 2752 22868 2792
rect 22252 2500 22484 2540
rect 21964 1364 22004 2500
rect 21964 1324 22100 1364
rect 21963 1196 22005 1205
rect 21963 1156 21964 1196
rect 22004 1156 22005 1196
rect 21963 1147 22005 1156
rect 21587 988 21716 1028
rect 21772 1112 21812 1121
rect 21484 944 21524 953
rect 21587 944 21627 988
rect 21772 944 21812 1072
rect 21964 1112 22004 1147
rect 21964 1061 22004 1072
rect 21387 860 21429 869
rect 21387 820 21388 860
rect 21428 820 21429 860
rect 21387 811 21429 820
rect 21387 524 21429 533
rect 21387 484 21388 524
rect 21428 484 21429 524
rect 21387 475 21429 484
rect 21388 80 21428 475
rect 21484 365 21524 904
rect 21580 904 21627 944
rect 21676 904 21812 944
rect 21868 944 21908 953
rect 22060 944 22100 1324
rect 22155 1112 22197 1121
rect 22155 1072 22156 1112
rect 22196 1072 22197 1112
rect 22155 1063 22197 1072
rect 22347 1112 22389 1121
rect 22347 1072 22348 1112
rect 22388 1072 22389 1112
rect 22347 1063 22389 1072
rect 22156 978 22196 1063
rect 22348 978 22388 1063
rect 21483 356 21525 365
rect 21483 316 21484 356
rect 21524 316 21525 356
rect 21483 307 21525 316
rect 21580 80 21620 904
rect 21676 197 21716 904
rect 21771 356 21813 365
rect 21771 316 21772 356
rect 21812 316 21813 356
rect 21771 307 21813 316
rect 21675 188 21717 197
rect 21675 148 21676 188
rect 21716 148 21717 188
rect 21675 139 21717 148
rect 21772 80 21812 307
rect 21868 281 21908 904
rect 21964 904 22100 944
rect 22251 944 22293 953
rect 22251 904 22252 944
rect 22292 904 22293 944
rect 21867 272 21909 281
rect 21867 232 21868 272
rect 21908 232 21909 272
rect 21867 223 21909 232
rect 21964 80 22004 904
rect 22251 895 22293 904
rect 22252 810 22292 895
rect 22444 776 22484 2500
rect 22540 1205 22580 1207
rect 22539 1196 22581 1205
rect 22539 1156 22540 1196
rect 22580 1156 22581 1196
rect 22539 1147 22581 1156
rect 22540 1112 22580 1147
rect 22540 1063 22580 1072
rect 22731 1112 22773 1121
rect 22731 1072 22732 1112
rect 22772 1072 22773 1112
rect 22731 1063 22773 1072
rect 22732 978 22772 1063
rect 22539 944 22581 953
rect 22539 904 22540 944
rect 22580 904 22581 944
rect 22539 895 22581 904
rect 22636 944 22676 953
rect 22348 736 22484 776
rect 22155 272 22197 281
rect 22155 232 22156 272
rect 22196 232 22197 272
rect 22155 223 22197 232
rect 22156 80 22196 223
rect 22348 80 22388 736
rect 22540 80 22580 895
rect 22636 533 22676 904
rect 22828 776 22868 2752
rect 23020 2540 23060 3172
rect 23116 2717 23156 3424
rect 23595 3464 23637 3473
rect 23595 3424 23596 3464
rect 23636 3424 23637 3464
rect 23595 3415 23637 3424
rect 23787 3464 23829 3473
rect 23787 3424 23788 3464
rect 23828 3424 23829 3464
rect 23787 3415 23829 3424
rect 23980 3464 24020 3473
rect 23596 3221 23636 3415
rect 23788 3330 23828 3415
rect 23980 3221 24020 3424
rect 24172 3464 24212 3473
rect 24172 3305 24212 3424
rect 24364 3464 24404 3473
rect 24171 3296 24213 3305
rect 24171 3256 24172 3296
rect 24212 3256 24213 3296
rect 24171 3247 24213 3256
rect 24364 3221 24404 3424
rect 24556 3464 24596 3473
rect 23595 3212 23637 3221
rect 23595 3172 23596 3212
rect 23636 3172 23637 3212
rect 23595 3163 23637 3172
rect 23692 3212 23732 3221
rect 23115 2708 23157 2717
rect 23115 2668 23116 2708
rect 23156 2668 23157 2708
rect 23115 2659 23157 2668
rect 23404 2633 23444 2718
rect 23403 2624 23445 2633
rect 23403 2584 23404 2624
rect 23444 2584 23445 2624
rect 23403 2575 23445 2584
rect 23596 2624 23636 3163
rect 23596 2575 23636 2584
rect 23500 2540 23540 2549
rect 23020 2500 23252 2540
rect 22924 1112 22964 1123
rect 22924 1037 22964 1072
rect 23115 1112 23157 1121
rect 23115 1072 23116 1112
rect 23156 1072 23157 1112
rect 23115 1063 23157 1072
rect 22923 1028 22965 1037
rect 22923 988 22924 1028
rect 22964 988 22965 1028
rect 22923 979 22965 988
rect 23116 978 23156 1063
rect 23019 944 23061 953
rect 23019 904 23020 944
rect 23060 904 23061 944
rect 23019 895 23061 904
rect 23020 810 23060 895
rect 23212 776 23252 2500
rect 23500 1364 23540 2500
rect 23692 1541 23732 3172
rect 23979 3212 24021 3221
rect 23979 3172 23980 3212
rect 24020 3172 24021 3212
rect 23979 3163 24021 3172
rect 24076 3212 24116 3221
rect 24076 2540 24116 3172
rect 24363 3212 24405 3221
rect 24363 3172 24364 3212
rect 24404 3172 24405 3212
rect 24363 3163 24405 3172
rect 24460 3212 24500 3221
rect 24460 2540 24500 3172
rect 24556 3053 24596 3424
rect 24652 3221 24692 4012
rect 24940 3977 24980 4096
rect 25036 4061 25076 4096
rect 25132 4136 25172 4171
rect 25132 4085 25172 4096
rect 25900 4136 25940 4255
rect 25900 4087 25940 4096
rect 26092 4136 26132 4147
rect 27916 4145 27956 4230
rect 26092 4061 26132 4096
rect 27915 4136 27957 4145
rect 27915 4096 27916 4136
rect 27956 4096 27957 4136
rect 27915 4087 27957 4096
rect 28012 4136 28052 4255
rect 32236 4145 32276 4230
rect 37228 4145 37268 4230
rect 28012 4087 28052 4096
rect 32140 4136 32180 4145
rect 25035 4052 25077 4061
rect 25035 4012 25036 4052
rect 25076 4012 25077 4052
rect 25035 4003 25077 4012
rect 26091 4052 26133 4061
rect 26091 4012 26092 4052
rect 26132 4012 26133 4052
rect 26091 4003 26133 4012
rect 31948 4052 31988 4061
rect 31988 4012 32084 4052
rect 31948 4003 31988 4012
rect 24844 3968 24884 3977
rect 24651 3212 24693 3221
rect 24651 3172 24652 3212
rect 24692 3172 24693 3212
rect 24651 3163 24693 3172
rect 24555 3044 24597 3053
rect 24555 3004 24556 3044
rect 24596 3004 24597 3044
rect 24555 2995 24597 3004
rect 24556 2885 24596 2995
rect 24555 2876 24597 2885
rect 24555 2836 24556 2876
rect 24596 2836 24597 2876
rect 24555 2827 24597 2836
rect 24076 2500 24404 2540
rect 24460 2500 24596 2540
rect 23691 1532 23733 1541
rect 23691 1492 23692 1532
rect 23732 1492 23733 1532
rect 23691 1483 23733 1492
rect 23500 1324 23636 1364
rect 23308 1205 23348 1207
rect 23307 1196 23349 1205
rect 23307 1156 23308 1196
rect 23348 1156 23349 1196
rect 23307 1147 23349 1156
rect 23308 1112 23348 1147
rect 23500 1121 23540 1206
rect 23308 1063 23348 1072
rect 23499 1112 23541 1121
rect 23499 1072 23500 1112
rect 23540 1072 23541 1112
rect 23499 1063 23541 1072
rect 23307 944 23349 953
rect 23307 904 23308 944
rect 23348 904 23349 944
rect 23307 895 23349 904
rect 23404 944 23444 953
rect 23596 944 23636 1324
rect 23692 1113 23732 1121
rect 23692 1112 23735 1113
rect 23732 1109 23735 1112
rect 23787 1112 23829 1121
rect 23787 1109 23788 1112
rect 23732 1072 23788 1109
rect 23828 1072 23829 1112
rect 23692 1069 23829 1072
rect 23692 1063 23732 1069
rect 23787 1063 23829 1069
rect 23884 1112 23924 1123
rect 24076 1112 24116 1121
rect 23884 1037 23924 1072
rect 23980 1072 24076 1112
rect 23883 1028 23925 1037
rect 23883 988 23884 1028
rect 23924 988 23925 1028
rect 23883 979 23925 988
rect 22732 736 22868 776
rect 23116 736 23252 776
rect 22635 524 22677 533
rect 22635 484 22636 524
rect 22676 484 22677 524
rect 22635 475 22677 484
rect 22732 80 22772 736
rect 22923 524 22965 533
rect 22923 484 22924 524
rect 22964 484 22965 524
rect 22923 475 22965 484
rect 22924 80 22964 475
rect 23116 80 23156 736
rect 23308 80 23348 895
rect 23404 281 23444 904
rect 23500 904 23636 944
rect 23787 944 23829 953
rect 23787 904 23788 944
rect 23828 904 23829 944
rect 23403 272 23445 281
rect 23403 232 23404 272
rect 23444 232 23445 272
rect 23403 223 23445 232
rect 23500 80 23540 904
rect 23787 895 23829 904
rect 23788 810 23828 895
rect 23883 524 23925 533
rect 23883 484 23884 524
rect 23924 484 23925 524
rect 23883 475 23925 484
rect 23691 272 23733 281
rect 23691 232 23692 272
rect 23732 232 23733 272
rect 23691 223 23733 232
rect 23692 80 23732 223
rect 23884 80 23924 475
rect 23980 449 24020 1072
rect 24076 1063 24116 1072
rect 24267 1112 24309 1121
rect 24267 1072 24268 1112
rect 24308 1072 24309 1112
rect 24267 1063 24309 1072
rect 24268 978 24308 1063
rect 24070 944 24112 953
rect 24171 944 24213 953
rect 24070 904 24071 944
rect 24111 904 24116 944
rect 24070 895 24116 904
rect 24171 904 24172 944
rect 24212 904 24213 944
rect 24171 895 24213 904
rect 23979 440 24021 449
rect 23979 400 23980 440
rect 24020 400 24021 440
rect 23979 391 24021 400
rect 24076 80 24116 895
rect 24172 810 24212 895
rect 24364 776 24404 2500
rect 24460 1205 24500 1207
rect 24459 1196 24501 1205
rect 24459 1156 24460 1196
rect 24500 1156 24501 1196
rect 24459 1147 24501 1156
rect 24460 1112 24500 1147
rect 24460 1063 24500 1072
rect 24459 944 24501 953
rect 24459 904 24460 944
rect 24500 904 24501 944
rect 24459 895 24501 904
rect 24268 736 24404 776
rect 24268 80 24308 736
rect 24460 80 24500 895
rect 24556 860 24596 2500
rect 24652 1952 24692 3163
rect 24844 2120 24884 3928
rect 24939 3968 24981 3977
rect 24939 3928 24940 3968
rect 24980 3928 24981 3968
rect 24939 3919 24981 3928
rect 25996 3968 26036 3977
rect 25323 3464 25365 3473
rect 25323 3424 25324 3464
rect 25364 3424 25365 3464
rect 25323 3415 25365 3424
rect 25515 3464 25557 3473
rect 25515 3424 25516 3464
rect 25556 3424 25557 3464
rect 25515 3415 25557 3424
rect 25708 3464 25748 3473
rect 25324 3330 25364 3415
rect 25516 3330 25556 3415
rect 25420 3212 25460 3221
rect 24844 2080 25076 2120
rect 24652 1903 24692 1912
rect 24843 1952 24885 1961
rect 24843 1912 24844 1952
rect 24884 1912 24885 1952
rect 24843 1903 24885 1912
rect 24844 1818 24884 1903
rect 24747 1700 24789 1709
rect 24747 1660 24748 1700
rect 24788 1660 24789 1700
rect 24747 1651 24789 1660
rect 24748 1566 24788 1651
rect 24652 1364 24692 1373
rect 24692 1324 24788 1364
rect 24652 1315 24692 1324
rect 24651 1196 24693 1205
rect 24651 1156 24652 1196
rect 24692 1156 24693 1196
rect 24651 1147 24693 1156
rect 24652 1112 24692 1147
rect 24652 1061 24692 1072
rect 24556 820 24692 860
rect 24652 80 24692 820
rect 24748 524 24788 1324
rect 24844 1121 24884 1206
rect 25036 1205 25076 2080
rect 25131 1700 25173 1709
rect 25131 1660 25132 1700
rect 25172 1660 25173 1700
rect 25131 1651 25173 1660
rect 25035 1196 25077 1205
rect 25035 1156 25036 1196
rect 25076 1156 25077 1196
rect 25035 1147 25077 1156
rect 24843 1112 24885 1121
rect 24843 1072 24844 1112
rect 24884 1072 24885 1112
rect 24843 1063 24885 1072
rect 25036 1112 25076 1147
rect 25036 1062 25076 1072
rect 24939 944 24981 953
rect 24939 904 24940 944
rect 24980 904 24981 944
rect 24939 895 24981 904
rect 24940 810 24980 895
rect 25132 860 25172 1651
rect 25227 944 25269 953
rect 25227 904 25228 944
rect 25268 904 25269 944
rect 25227 895 25269 904
rect 25036 820 25172 860
rect 24748 484 24884 524
rect 24844 80 24884 484
rect 25036 80 25076 820
rect 25228 80 25268 895
rect 25420 80 25460 3172
rect 25708 2465 25748 3424
rect 25899 3464 25941 3473
rect 25996 3464 26036 3928
rect 27724 3968 27764 3977
rect 27764 3928 28340 3968
rect 27724 3919 27764 3928
rect 27339 3800 27381 3809
rect 27339 3760 27340 3800
rect 27380 3760 27381 3800
rect 27339 3751 27381 3760
rect 26956 3557 26996 3588
rect 26955 3548 26997 3557
rect 26955 3508 26956 3548
rect 26996 3508 26997 3548
rect 26955 3499 26997 3508
rect 25899 3424 25900 3464
rect 25940 3424 26036 3464
rect 26092 3464 26132 3473
rect 25899 3415 25941 3424
rect 25900 3330 25940 3415
rect 25804 3212 25844 3221
rect 25707 2456 25749 2465
rect 25707 2416 25708 2456
rect 25748 2416 25749 2456
rect 25707 2407 25749 2416
rect 25515 1448 25557 1457
rect 25515 1408 25516 1448
rect 25556 1408 25557 1448
rect 25515 1399 25557 1408
rect 25516 1121 25556 1399
rect 25707 1280 25749 1289
rect 25707 1240 25708 1280
rect 25748 1240 25749 1280
rect 25707 1231 25749 1240
rect 25515 1112 25557 1121
rect 25515 1072 25516 1112
rect 25556 1072 25557 1112
rect 25515 1063 25557 1072
rect 25708 1112 25748 1231
rect 25708 1063 25748 1072
rect 25516 978 25556 1063
rect 25612 944 25652 953
rect 25612 533 25652 904
rect 25707 944 25749 953
rect 25707 904 25708 944
rect 25748 904 25749 944
rect 25707 895 25749 904
rect 25611 524 25653 533
rect 25611 484 25612 524
rect 25652 484 25653 524
rect 25611 475 25653 484
rect 25708 356 25748 895
rect 25612 316 25748 356
rect 25612 80 25652 316
rect 25804 80 25844 3172
rect 26092 3137 26132 3424
rect 26283 3464 26325 3473
rect 26283 3424 26284 3464
rect 26324 3424 26325 3464
rect 26283 3415 26325 3424
rect 26763 3464 26805 3473
rect 26763 3424 26764 3464
rect 26804 3424 26805 3464
rect 26763 3415 26805 3424
rect 26956 3464 26996 3499
rect 26188 3212 26228 3221
rect 26091 3128 26133 3137
rect 26091 3088 26092 3128
rect 26132 3088 26133 3128
rect 26091 3079 26133 3088
rect 26092 2213 26132 3079
rect 26091 2204 26133 2213
rect 26091 2164 26092 2204
rect 26132 2164 26133 2204
rect 26091 2155 26133 2164
rect 25900 1952 25940 1961
rect 25900 1289 25940 1912
rect 26092 1952 26132 1961
rect 26092 1877 26132 1912
rect 25996 1868 26036 1877
rect 25899 1280 25941 1289
rect 25899 1240 25900 1280
rect 25940 1240 25941 1280
rect 25899 1231 25941 1240
rect 25900 1112 25940 1123
rect 25996 1121 26036 1828
rect 26091 1868 26133 1877
rect 26091 1828 26092 1868
rect 26132 1828 26133 1868
rect 26091 1819 26133 1828
rect 26092 1373 26132 1819
rect 26091 1364 26133 1373
rect 26091 1324 26092 1364
rect 26132 1324 26133 1364
rect 26091 1315 26133 1324
rect 25900 1037 25940 1072
rect 25995 1112 26037 1121
rect 25995 1072 25996 1112
rect 26036 1072 26037 1112
rect 25995 1063 26037 1072
rect 26092 1112 26132 1123
rect 26092 1037 26132 1072
rect 25899 1028 25941 1037
rect 25899 988 25900 1028
rect 25940 988 25941 1028
rect 25899 979 25941 988
rect 26091 1028 26133 1037
rect 26091 988 26092 1028
rect 26132 988 26133 1028
rect 26091 979 26133 988
rect 25996 944 26036 953
rect 25996 701 26036 904
rect 25995 692 26037 701
rect 25995 652 25996 692
rect 26036 652 26037 692
rect 25995 643 26037 652
rect 25995 524 26037 533
rect 25995 484 25996 524
rect 26036 484 26037 524
rect 25995 475 26037 484
rect 25996 80 26036 475
rect 26188 80 26228 3172
rect 26284 2624 26324 3415
rect 26764 3330 26804 3415
rect 26860 3212 26900 3221
rect 26572 2633 26612 2718
rect 26380 2624 26420 2633
rect 26284 2584 26380 2624
rect 26380 2575 26420 2584
rect 26571 2624 26613 2633
rect 26571 2584 26572 2624
rect 26612 2584 26613 2624
rect 26571 2575 26613 2584
rect 26476 2540 26516 2549
rect 26860 2540 26900 3172
rect 26956 3053 26996 3424
rect 27147 3464 27189 3473
rect 27147 3424 27148 3464
rect 27188 3424 27189 3464
rect 27147 3415 27189 3424
rect 27340 3464 27380 3751
rect 27627 3716 27669 3725
rect 27627 3676 27628 3716
rect 27668 3676 27669 3716
rect 27627 3667 27669 3676
rect 27340 3415 27380 3424
rect 27628 3464 27668 3667
rect 27628 3415 27668 3424
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 27148 3330 27188 3415
rect 27244 3212 27284 3221
rect 27724 3212 27764 3221
rect 26955 3044 26997 3053
rect 26955 3004 26956 3044
rect 26996 3004 26997 3044
rect 26955 2995 26997 3004
rect 27244 2540 27284 3172
rect 27628 3172 27724 3212
rect 27628 2540 27668 3172
rect 27724 3163 27764 3172
rect 27820 2624 27860 3415
rect 28108 2633 28148 2718
rect 27916 2624 27956 2633
rect 27820 2584 27916 2624
rect 27916 2575 27956 2584
rect 28107 2624 28149 2633
rect 28107 2584 28108 2624
rect 28148 2584 28149 2624
rect 28107 2575 28149 2584
rect 28012 2540 28052 2549
rect 26860 2500 26996 2540
rect 27244 2500 27380 2540
rect 27628 2500 27764 2540
rect 26476 2120 26516 2500
rect 26476 2080 26612 2120
rect 26284 1112 26324 1121
rect 26284 785 26324 1072
rect 26475 1112 26517 1121
rect 26475 1072 26476 1112
rect 26516 1072 26517 1112
rect 26475 1063 26517 1072
rect 26380 953 26420 1038
rect 26476 978 26516 1063
rect 26379 944 26421 953
rect 26379 904 26380 944
rect 26420 904 26421 944
rect 26379 895 26421 904
rect 26283 776 26325 785
rect 26283 736 26284 776
rect 26324 736 26325 776
rect 26283 727 26325 736
rect 26379 692 26421 701
rect 26379 652 26380 692
rect 26420 652 26421 692
rect 26379 643 26421 652
rect 26380 80 26420 643
rect 26572 80 26612 2080
rect 26668 1205 26708 1207
rect 26667 1196 26709 1205
rect 26667 1156 26668 1196
rect 26708 1156 26709 1196
rect 26667 1147 26709 1156
rect 26668 1112 26708 1147
rect 26668 1063 26708 1072
rect 26859 1112 26901 1121
rect 26859 1072 26860 1112
rect 26900 1072 26901 1112
rect 26859 1063 26901 1072
rect 26860 978 26900 1063
rect 26667 944 26709 953
rect 26667 904 26668 944
rect 26708 904 26709 944
rect 26667 895 26709 904
rect 26764 944 26804 953
rect 26668 524 26708 895
rect 26764 701 26804 904
rect 26763 692 26805 701
rect 26763 652 26764 692
rect 26804 652 26805 692
rect 26763 643 26805 652
rect 26668 484 26804 524
rect 26764 80 26804 484
rect 26956 80 26996 2500
rect 27052 1112 27092 1121
rect 27052 617 27092 1072
rect 27243 1112 27285 1121
rect 27243 1072 27244 1112
rect 27284 1072 27285 1112
rect 27243 1063 27285 1072
rect 27148 953 27188 1038
rect 27244 978 27284 1063
rect 27147 944 27189 953
rect 27147 904 27148 944
rect 27188 904 27189 944
rect 27147 895 27189 904
rect 27147 692 27189 701
rect 27147 652 27148 692
rect 27188 652 27189 692
rect 27147 643 27189 652
rect 27051 608 27093 617
rect 27051 568 27052 608
rect 27092 568 27093 608
rect 27051 559 27093 568
rect 27052 281 27092 559
rect 27051 272 27093 281
rect 27051 232 27052 272
rect 27092 232 27093 272
rect 27051 223 27093 232
rect 27148 80 27188 643
rect 27340 80 27380 2500
rect 27435 1280 27477 1289
rect 27435 1240 27436 1280
rect 27476 1240 27477 1280
rect 27435 1231 27477 1240
rect 27436 1112 27476 1231
rect 27436 1063 27476 1072
rect 27627 1112 27669 1121
rect 27627 1072 27628 1112
rect 27668 1072 27669 1112
rect 27627 1063 27669 1072
rect 27628 978 27668 1063
rect 27435 944 27477 953
rect 27435 904 27436 944
rect 27476 904 27477 944
rect 27435 895 27477 904
rect 27532 944 27572 953
rect 27436 524 27476 895
rect 27532 701 27572 904
rect 27531 692 27573 701
rect 27531 652 27532 692
rect 27572 652 27573 692
rect 27531 643 27573 652
rect 27436 484 27572 524
rect 27532 80 27572 484
rect 27724 80 27764 2500
rect 28012 2120 28052 2500
rect 28012 2080 28148 2120
rect 27820 1112 27860 1121
rect 27820 869 27860 1072
rect 28011 1112 28053 1121
rect 28011 1072 28012 1112
rect 28052 1072 28053 1112
rect 28011 1063 28053 1072
rect 27916 953 27956 1038
rect 28012 978 28052 1063
rect 27915 944 27957 953
rect 27915 904 27916 944
rect 27956 904 27957 944
rect 27915 895 27957 904
rect 27819 860 27861 869
rect 27819 820 27820 860
rect 27860 820 27861 860
rect 27819 811 27861 820
rect 27820 533 27860 811
rect 27915 692 27957 701
rect 27915 652 27916 692
rect 27956 652 27957 692
rect 27915 643 27957 652
rect 27819 524 27861 533
rect 27819 484 27820 524
rect 27860 484 27861 524
rect 27819 475 27861 484
rect 27916 80 27956 643
rect 28108 80 28148 2080
rect 28204 1205 28244 1207
rect 28203 1196 28245 1205
rect 28203 1156 28204 1196
rect 28244 1156 28245 1196
rect 28203 1147 28245 1156
rect 28204 1112 28244 1147
rect 28300 1121 28340 3928
rect 31564 3592 31892 3632
rect 28396 3557 28436 3588
rect 28395 3548 28437 3557
rect 28395 3508 28396 3548
rect 28436 3508 28437 3548
rect 28395 3499 28437 3508
rect 28396 3464 28436 3499
rect 28396 3389 28436 3424
rect 28588 3464 28628 3475
rect 28588 3389 28628 3424
rect 28780 3464 28820 3473
rect 28395 3380 28437 3389
rect 28395 3340 28396 3380
rect 28436 3340 28437 3380
rect 28395 3331 28437 3340
rect 28587 3380 28629 3389
rect 28587 3340 28588 3380
rect 28628 3340 28629 3380
rect 28587 3331 28629 3340
rect 28492 3212 28532 3221
rect 28204 1063 28244 1072
rect 28299 1112 28341 1121
rect 28396 1112 28436 1121
rect 28299 1072 28300 1112
rect 28340 1072 28396 1112
rect 28299 1063 28341 1072
rect 28396 1063 28436 1072
rect 28203 944 28245 953
rect 28203 904 28204 944
rect 28244 904 28245 944
rect 28203 895 28245 904
rect 28300 944 28340 953
rect 28204 524 28244 895
rect 28300 701 28340 904
rect 28299 692 28341 701
rect 28299 652 28300 692
rect 28340 652 28341 692
rect 28299 643 28341 652
rect 28204 484 28340 524
rect 28300 80 28340 484
rect 28492 80 28532 3172
rect 28780 2969 28820 3424
rect 28972 3464 29012 3475
rect 28972 3389 29012 3424
rect 29164 3464 29204 3473
rect 28971 3380 29013 3389
rect 28971 3340 28972 3380
rect 29012 3340 29013 3380
rect 28971 3331 29013 3340
rect 28876 3212 28916 3221
rect 28779 2960 28821 2969
rect 28779 2920 28780 2960
rect 28820 2920 28821 2960
rect 28779 2911 28821 2920
rect 28588 1112 28628 1121
rect 28588 617 28628 1072
rect 28779 1112 28821 1121
rect 28779 1072 28780 1112
rect 28820 1072 28821 1112
rect 28779 1063 28821 1072
rect 28780 978 28820 1063
rect 28683 944 28725 953
rect 28683 904 28684 944
rect 28724 904 28725 944
rect 28683 895 28725 904
rect 28684 810 28724 895
rect 28683 692 28725 701
rect 28683 652 28684 692
rect 28724 652 28725 692
rect 28683 643 28725 652
rect 28587 608 28629 617
rect 28587 568 28588 608
rect 28628 568 28629 608
rect 28587 559 28629 568
rect 28684 80 28724 643
rect 28779 608 28821 617
rect 28779 568 28780 608
rect 28820 568 28821 608
rect 28779 559 28821 568
rect 28780 197 28820 559
rect 28779 188 28821 197
rect 28779 148 28780 188
rect 28820 148 28821 188
rect 28779 139 28821 148
rect 28876 80 28916 3172
rect 29164 2717 29204 3424
rect 29356 3464 29396 3475
rect 29356 3389 29396 3424
rect 29644 3464 29684 3473
rect 29644 3389 29684 3424
rect 29835 3464 29877 3473
rect 29835 3424 29836 3464
rect 29876 3424 29877 3464
rect 29835 3415 29877 3424
rect 30028 3464 30068 3475
rect 29355 3380 29397 3389
rect 29355 3340 29356 3380
rect 29396 3340 29397 3380
rect 29355 3331 29397 3340
rect 29643 3380 29685 3389
rect 29643 3340 29644 3380
rect 29684 3340 29685 3380
rect 29643 3331 29685 3340
rect 29260 3212 29300 3221
rect 29163 2708 29205 2717
rect 29163 2668 29164 2708
rect 29204 2668 29205 2708
rect 29163 2659 29205 2668
rect 28971 1532 29013 1541
rect 28971 1492 28972 1532
rect 29012 1492 29013 1532
rect 28971 1483 29013 1492
rect 28972 1121 29012 1483
rect 29164 1205 29204 1207
rect 29163 1196 29205 1205
rect 29163 1156 29164 1196
rect 29204 1156 29205 1196
rect 29163 1147 29205 1156
rect 28971 1112 29013 1121
rect 28971 1072 28972 1112
rect 29012 1072 29013 1112
rect 28971 1063 29013 1072
rect 29164 1112 29204 1147
rect 29164 1063 29204 1072
rect 28971 944 29013 953
rect 28971 904 28972 944
rect 29012 904 29013 944
rect 28971 895 29013 904
rect 29068 944 29108 953
rect 28972 356 29012 895
rect 29068 533 29108 904
rect 29067 524 29109 533
rect 29067 484 29068 524
rect 29108 484 29109 524
rect 29067 475 29109 484
rect 28972 316 29108 356
rect 29068 80 29108 316
rect 29260 80 29300 3172
rect 29644 3044 29684 3331
rect 29836 3330 29876 3415
rect 30028 3389 30068 3424
rect 30219 3464 30261 3473
rect 30219 3424 30220 3464
rect 30260 3424 30261 3464
rect 30219 3415 30261 3424
rect 30412 3464 30452 3475
rect 30027 3380 30069 3389
rect 30027 3340 30028 3380
rect 30068 3340 30069 3380
rect 30027 3331 30069 3340
rect 30220 3330 30260 3415
rect 30412 3389 30452 3424
rect 30604 3464 30644 3473
rect 31276 3464 31316 3473
rect 30644 3424 30740 3464
rect 30604 3415 30644 3424
rect 30411 3380 30453 3389
rect 30411 3340 30412 3380
rect 30452 3340 30453 3380
rect 30411 3331 30453 3340
rect 29740 3212 29780 3221
rect 30124 3212 30164 3221
rect 30508 3212 30548 3221
rect 29780 3172 30068 3212
rect 29740 3163 29780 3172
rect 29644 3004 29780 3044
rect 29740 2633 29780 3004
rect 29547 2624 29589 2633
rect 29547 2584 29548 2624
rect 29588 2584 29589 2624
rect 29547 2575 29589 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 29548 2490 29588 2575
rect 29644 2540 29684 2549
rect 29547 1196 29589 1205
rect 29547 1156 29548 1196
rect 29588 1156 29589 1196
rect 29547 1147 29589 1156
rect 29356 1112 29396 1121
rect 29356 617 29396 1072
rect 29548 1112 29588 1147
rect 29548 1061 29588 1072
rect 29452 944 29492 953
rect 29452 701 29492 904
rect 29451 692 29493 701
rect 29451 652 29452 692
rect 29492 652 29493 692
rect 29451 643 29493 652
rect 29355 608 29397 617
rect 29355 568 29356 608
rect 29396 568 29397 608
rect 29355 559 29397 568
rect 29356 197 29396 559
rect 29451 524 29493 533
rect 29451 484 29452 524
rect 29492 484 29493 524
rect 29451 475 29493 484
rect 29355 188 29397 197
rect 29355 148 29356 188
rect 29396 148 29397 188
rect 29355 139 29397 148
rect 29452 80 29492 475
rect 29644 80 29684 2500
rect 29740 2490 29780 2575
rect 29931 1196 29973 1205
rect 29931 1156 29932 1196
rect 29972 1156 29973 1196
rect 29931 1147 29973 1156
rect 29739 1112 29781 1121
rect 29739 1072 29740 1112
rect 29780 1072 29781 1112
rect 29739 1063 29781 1072
rect 29932 1112 29972 1147
rect 29740 978 29780 1063
rect 29932 1061 29972 1072
rect 29836 953 29876 1038
rect 29835 944 29877 953
rect 29835 904 29836 944
rect 29876 904 29877 944
rect 29835 895 29877 904
rect 29835 692 29877 701
rect 29835 652 29836 692
rect 29876 652 29877 692
rect 29835 643 29877 652
rect 29836 80 29876 643
rect 30028 80 30068 3172
rect 30164 3172 30260 3212
rect 30124 3163 30164 3172
rect 30220 1364 30260 3172
rect 30548 3172 30644 3212
rect 30508 3163 30548 3172
rect 30220 1324 30452 1364
rect 30124 1121 30164 1206
rect 30315 1196 30357 1205
rect 30315 1156 30316 1196
rect 30356 1156 30357 1196
rect 30315 1147 30357 1156
rect 30123 1112 30165 1121
rect 30123 1072 30124 1112
rect 30164 1072 30165 1112
rect 30123 1063 30165 1072
rect 30316 1112 30356 1147
rect 30316 1061 30356 1072
rect 30123 944 30165 953
rect 30123 904 30124 944
rect 30164 904 30165 944
rect 30123 895 30165 904
rect 30220 944 30260 953
rect 30124 524 30164 895
rect 30220 701 30260 904
rect 30219 692 30261 701
rect 30219 652 30220 692
rect 30260 652 30261 692
rect 30219 643 30261 652
rect 30124 484 30260 524
rect 30220 80 30260 484
rect 30412 80 30452 1324
rect 30508 1112 30548 1121
rect 30508 953 30548 1072
rect 30507 944 30549 953
rect 30507 904 30508 944
rect 30548 904 30549 944
rect 30604 944 30644 3172
rect 30700 2885 30740 3424
rect 31180 3424 31276 3464
rect 30699 2876 30741 2885
rect 30699 2836 30700 2876
rect 30740 2836 30741 2876
rect 30699 2827 30741 2836
rect 30699 2624 30741 2633
rect 30699 2584 30700 2624
rect 30740 2584 30741 2624
rect 30699 2575 30741 2584
rect 30891 2624 30933 2633
rect 30891 2584 30892 2624
rect 30932 2584 30933 2624
rect 30891 2575 30933 2584
rect 30700 2490 30740 2575
rect 30796 2540 30836 2549
rect 30700 1373 30740 1458
rect 30699 1364 30741 1373
rect 30699 1324 30700 1364
rect 30740 1324 30741 1364
rect 30796 1364 30836 2500
rect 30892 2490 30932 2575
rect 31180 2213 31220 3424
rect 31276 3415 31316 3424
rect 31467 3464 31509 3473
rect 31467 3424 31468 3464
rect 31508 3424 31509 3464
rect 31467 3415 31509 3424
rect 31468 3330 31508 3415
rect 31372 3212 31412 3221
rect 31276 3172 31372 3212
rect 31179 2204 31221 2213
rect 31179 2164 31180 2204
rect 31220 2164 31221 2204
rect 31179 2155 31221 2164
rect 31180 1709 31220 2155
rect 31179 1700 31221 1709
rect 31179 1660 31180 1700
rect 31220 1660 31221 1700
rect 31179 1651 31221 1660
rect 30796 1324 31220 1364
rect 30699 1315 30741 1324
rect 30700 1121 30740 1206
rect 30699 1112 30741 1121
rect 30699 1072 30700 1112
rect 30740 1072 30741 1112
rect 30699 1063 30741 1072
rect 30891 1112 30933 1121
rect 30891 1072 30892 1112
rect 30932 1072 30933 1112
rect 30891 1063 30933 1072
rect 31083 1112 31125 1121
rect 31083 1072 31084 1112
rect 31124 1072 31125 1112
rect 31083 1063 31125 1072
rect 30892 978 30932 1063
rect 31084 978 31124 1063
rect 30987 944 31029 953
rect 30604 904 30836 944
rect 30507 895 30549 904
rect 30603 692 30645 701
rect 30603 652 30604 692
rect 30644 652 30645 692
rect 30603 643 30645 652
rect 30604 80 30644 643
rect 30796 80 30836 904
rect 30987 904 30988 944
rect 31028 904 31029 944
rect 30987 895 31029 904
rect 30988 810 31028 895
rect 30987 608 31029 617
rect 30987 568 30988 608
rect 31028 568 31029 608
rect 30987 559 31029 568
rect 30988 80 31028 559
rect 31180 80 31220 1324
rect 31276 701 31316 3172
rect 31372 3163 31412 3172
rect 31564 3137 31604 3592
rect 31659 3464 31701 3473
rect 31659 3424 31660 3464
rect 31700 3424 31701 3464
rect 31659 3415 31701 3424
rect 31852 3464 31892 3592
rect 32044 3473 32084 4012
rect 32140 3893 32180 4096
rect 32235 4136 32277 4145
rect 32620 4136 32660 4145
rect 32235 4096 32236 4136
rect 32276 4096 32277 4136
rect 32235 4087 32277 4096
rect 32524 4096 32620 4136
rect 32524 3977 32564 4096
rect 32620 4087 32660 4096
rect 32811 4136 32853 4145
rect 32811 4096 32812 4136
rect 32852 4096 32853 4136
rect 32811 4087 32853 4096
rect 32908 4136 32948 4145
rect 32812 4002 32852 4087
rect 32235 3968 32277 3977
rect 32235 3928 32236 3968
rect 32276 3928 32277 3968
rect 32235 3919 32277 3928
rect 32523 3968 32565 3977
rect 32523 3928 32524 3968
rect 32564 3928 32565 3968
rect 32523 3919 32565 3928
rect 32620 3968 32660 3977
rect 32660 3928 32756 3968
rect 32620 3919 32660 3928
rect 32139 3884 32181 3893
rect 32139 3844 32140 3884
rect 32180 3844 32181 3884
rect 32139 3835 32181 3844
rect 32236 3834 32276 3919
rect 32235 3632 32277 3641
rect 32235 3592 32236 3632
rect 32276 3592 32277 3632
rect 32235 3583 32277 3592
rect 31852 3415 31892 3424
rect 32043 3464 32085 3473
rect 32043 3424 32044 3464
rect 32084 3424 32085 3464
rect 32043 3415 32085 3424
rect 32236 3464 32276 3583
rect 32236 3415 32276 3424
rect 32427 3464 32469 3473
rect 32427 3424 32428 3464
rect 32468 3424 32469 3464
rect 32427 3415 32469 3424
rect 32620 3464 32660 3473
rect 31563 3128 31605 3137
rect 31563 3088 31564 3128
rect 31604 3088 31605 3128
rect 31563 3079 31605 3088
rect 31564 2129 31604 3079
rect 31660 3044 31700 3415
rect 32044 3330 32084 3415
rect 32428 3330 32468 3415
rect 31756 3221 31796 3306
rect 31755 3212 31797 3221
rect 31755 3172 31756 3212
rect 31796 3172 31797 3212
rect 31755 3163 31797 3172
rect 32140 3212 32180 3221
rect 32524 3212 32564 3221
rect 32180 3172 32468 3212
rect 32140 3163 32180 3172
rect 31660 3004 31892 3044
rect 31659 2624 31701 2633
rect 31659 2584 31660 2624
rect 31700 2584 31701 2624
rect 31659 2575 31701 2584
rect 31852 2624 31892 3004
rect 31852 2575 31892 2584
rect 31660 2490 31700 2575
rect 31756 2540 31796 2549
rect 31563 2120 31605 2129
rect 31563 2080 31564 2120
rect 31604 2080 31605 2120
rect 31563 2071 31605 2080
rect 31756 1784 31796 2500
rect 31948 1961 31988 2046
rect 31947 1952 31989 1961
rect 32140 1952 32180 1963
rect 31947 1912 31948 1952
rect 31988 1912 32084 1952
rect 31947 1903 31989 1912
rect 31564 1744 31796 1784
rect 31467 1616 31509 1625
rect 31467 1576 31468 1616
rect 31508 1576 31509 1616
rect 31467 1567 31509 1576
rect 31468 1121 31508 1567
rect 31467 1112 31509 1121
rect 31467 1072 31468 1112
rect 31508 1072 31509 1112
rect 31467 1063 31509 1072
rect 31468 978 31508 1063
rect 31371 944 31413 953
rect 31371 904 31372 944
rect 31412 904 31413 944
rect 31371 895 31413 904
rect 31275 692 31317 701
rect 31275 652 31276 692
rect 31316 652 31317 692
rect 31275 643 31317 652
rect 31372 80 31412 895
rect 31564 80 31604 1744
rect 31948 1700 31988 1709
rect 31756 1660 31948 1700
rect 31660 1289 31700 1374
rect 31659 1280 31701 1289
rect 31659 1240 31660 1280
rect 31700 1240 31701 1280
rect 31659 1231 31701 1240
rect 31659 1112 31701 1121
rect 31659 1072 31660 1112
rect 31700 1072 31701 1112
rect 31659 1063 31701 1072
rect 31660 978 31700 1063
rect 31756 80 31796 1660
rect 31948 1651 31988 1660
rect 31851 1364 31893 1373
rect 31851 1324 31852 1364
rect 31892 1324 31893 1364
rect 31851 1315 31893 1324
rect 31852 1205 31892 1315
rect 31851 1196 31893 1205
rect 31851 1156 31852 1196
rect 31892 1156 31893 1196
rect 31851 1147 31893 1156
rect 31852 1112 31892 1147
rect 32044 1121 32084 1912
rect 32140 1877 32180 1912
rect 32139 1868 32181 1877
rect 32139 1828 32140 1868
rect 32180 1828 32181 1868
rect 32139 1819 32181 1828
rect 32139 1280 32181 1289
rect 32139 1240 32140 1280
rect 32180 1240 32181 1280
rect 32428 1280 32468 3172
rect 32524 1457 32564 3172
rect 32620 3053 32660 3424
rect 32619 3044 32661 3053
rect 32619 3004 32620 3044
rect 32660 3004 32661 3044
rect 32619 2995 32661 3004
rect 32620 1793 32660 2995
rect 32716 1961 32756 3928
rect 32908 3893 32948 4096
rect 37227 4136 37269 4145
rect 37227 4096 37228 4136
rect 37268 4096 37269 4136
rect 37227 4087 37269 4096
rect 37324 4136 37364 4339
rect 37707 4220 37749 4229
rect 37707 4180 37708 4220
rect 37748 4180 37749 4220
rect 37707 4171 37749 4180
rect 37996 4180 38132 4220
rect 37324 4087 37364 4096
rect 37708 4136 37748 4171
rect 37708 4085 37748 4096
rect 37803 4136 37845 4145
rect 37996 4136 38036 4180
rect 37803 4096 37804 4136
rect 37844 4096 37940 4136
rect 37803 4087 37845 4096
rect 37516 4052 37556 4061
rect 37227 3968 37269 3977
rect 37227 3928 37228 3968
rect 37268 3928 37269 3968
rect 37227 3919 37269 3928
rect 32907 3884 32949 3893
rect 32907 3844 32908 3884
rect 32948 3844 32949 3884
rect 32907 3835 32949 3844
rect 37228 3834 37268 3919
rect 33003 3800 33045 3809
rect 33003 3760 33004 3800
rect 33044 3760 33045 3800
rect 33003 3751 33045 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 35691 3800 35733 3809
rect 35691 3760 35692 3800
rect 35732 3760 35733 3800
rect 35691 3751 35733 3760
rect 33004 3641 33044 3751
rect 33387 3716 33429 3725
rect 33387 3676 33388 3716
rect 33428 3676 33429 3716
rect 33387 3667 33429 3676
rect 33003 3632 33045 3641
rect 33003 3592 33004 3632
rect 33044 3592 33045 3632
rect 33003 3583 33045 3592
rect 32811 3464 32853 3473
rect 32811 3424 32812 3464
rect 32852 3424 32853 3464
rect 32811 3415 32853 3424
rect 33004 3464 33044 3583
rect 33004 3415 33044 3424
rect 33195 3464 33237 3473
rect 33195 3424 33196 3464
rect 33236 3424 33237 3464
rect 33195 3415 33237 3424
rect 33388 3464 33428 3667
rect 33676 3592 33908 3632
rect 33676 3548 33716 3592
rect 33676 3499 33716 3508
rect 33388 3415 33428 3424
rect 33579 3464 33621 3473
rect 33579 3424 33580 3464
rect 33620 3424 33621 3464
rect 33579 3415 33621 3424
rect 33772 3464 33812 3473
rect 32812 3330 32852 3415
rect 33196 3330 33236 3415
rect 33580 3330 33620 3415
rect 32908 3212 32948 3221
rect 33292 3212 33332 3221
rect 32715 1952 32757 1961
rect 32715 1912 32716 1952
rect 32756 1912 32757 1952
rect 32715 1903 32757 1912
rect 32619 1784 32661 1793
rect 32619 1744 32620 1784
rect 32660 1744 32661 1784
rect 32619 1735 32661 1744
rect 32523 1448 32565 1457
rect 32523 1408 32524 1448
rect 32564 1408 32565 1448
rect 32523 1399 32565 1408
rect 32619 1280 32661 1289
rect 32428 1240 32564 1280
rect 32139 1231 32181 1240
rect 31852 1062 31892 1072
rect 32043 1112 32085 1121
rect 32043 1072 32044 1112
rect 32084 1072 32085 1112
rect 32043 1063 32085 1072
rect 32044 978 32084 1063
rect 31948 944 31988 953
rect 31948 860 31988 904
rect 31948 820 32084 860
rect 31947 692 31989 701
rect 31947 652 31948 692
rect 31988 652 31989 692
rect 31947 643 31989 652
rect 31948 80 31988 643
rect 32044 449 32084 820
rect 32043 440 32085 449
rect 32043 400 32044 440
rect 32084 400 32085 440
rect 32043 391 32085 400
rect 32140 80 32180 1231
rect 32236 1205 32276 1220
rect 32235 1196 32277 1205
rect 32235 1156 32236 1196
rect 32276 1156 32277 1196
rect 32235 1147 32277 1156
rect 32236 1125 32276 1147
rect 32236 1076 32276 1085
rect 32427 1112 32469 1121
rect 32427 1072 32428 1112
rect 32468 1072 32469 1112
rect 32427 1063 32469 1072
rect 32428 978 32468 1063
rect 32235 944 32277 953
rect 32235 904 32236 944
rect 32276 904 32277 944
rect 32235 895 32277 904
rect 32332 944 32372 953
rect 32524 944 32564 1240
rect 32619 1240 32620 1280
rect 32660 1240 32661 1280
rect 32619 1231 32661 1240
rect 32620 1112 32660 1231
rect 32620 1063 32660 1072
rect 32811 1112 32853 1121
rect 32811 1072 32812 1112
rect 32852 1072 32853 1112
rect 32811 1063 32853 1072
rect 32812 978 32852 1063
rect 32715 944 32757 953
rect 32524 904 32660 944
rect 32236 356 32276 895
rect 32332 533 32372 904
rect 32620 692 32660 904
rect 32715 904 32716 944
rect 32756 904 32757 944
rect 32715 895 32757 904
rect 32716 810 32756 895
rect 32908 701 32948 3172
rect 33196 3172 33292 3212
rect 33196 1448 33236 3172
rect 33292 3163 33332 3172
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 33772 2633 33812 3424
rect 33771 2624 33813 2633
rect 33771 2584 33772 2624
rect 33812 2584 33813 2624
rect 33771 2575 33813 2584
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 33196 1408 33243 1448
rect 33203 1364 33243 1408
rect 33203 1324 33716 1364
rect 33196 1121 33236 1206
rect 33195 1112 33237 1121
rect 33004 1101 33044 1110
rect 33195 1072 33196 1112
rect 33236 1072 33237 1112
rect 33195 1063 33237 1072
rect 33388 1112 33428 1123
rect 33004 1028 33044 1061
rect 33388 1037 33428 1072
rect 33579 1112 33621 1121
rect 33579 1072 33580 1112
rect 33620 1072 33621 1112
rect 33579 1063 33621 1072
rect 33003 988 33044 1028
rect 33387 1028 33429 1037
rect 33387 988 33388 1028
rect 33428 988 33429 1028
rect 33003 860 33043 988
rect 33387 979 33429 988
rect 33580 978 33620 1063
rect 33100 944 33140 953
rect 33291 944 33333 953
rect 33140 904 33236 944
rect 33100 895 33140 904
rect 33003 820 33044 860
rect 32907 692 32949 701
rect 32620 652 32756 692
rect 32331 524 32373 533
rect 32331 484 32332 524
rect 32372 484 32373 524
rect 32331 475 32373 484
rect 32523 440 32565 449
rect 32523 400 32524 440
rect 32564 400 32565 440
rect 32523 391 32565 400
rect 32236 316 32372 356
rect 32332 80 32372 316
rect 32524 80 32564 391
rect 32716 80 32756 652
rect 32907 652 32908 692
rect 32948 652 32949 692
rect 32907 643 32949 652
rect 32907 524 32949 533
rect 32907 484 32908 524
rect 32948 484 32949 524
rect 32907 475 32949 484
rect 32908 80 32948 475
rect 33004 281 33044 820
rect 33099 608 33141 617
rect 33099 568 33100 608
rect 33140 568 33141 608
rect 33099 559 33141 568
rect 33003 272 33045 281
rect 33003 232 33004 272
rect 33044 232 33045 272
rect 33003 223 33045 232
rect 33100 80 33140 559
rect 33196 533 33236 904
rect 33291 904 33292 944
rect 33332 904 33333 944
rect 33291 895 33333 904
rect 33484 944 33524 953
rect 33195 524 33237 533
rect 33195 484 33196 524
rect 33236 484 33237 524
rect 33195 475 33237 484
rect 33292 80 33332 895
rect 33484 860 33524 904
rect 33484 820 33620 860
rect 33483 692 33525 701
rect 33483 652 33484 692
rect 33524 652 33525 692
rect 33483 643 33525 652
rect 33484 80 33524 643
rect 33580 449 33620 820
rect 33676 692 33716 1324
rect 33868 1289 33908 3592
rect 34155 3548 34197 3557
rect 34155 3508 34156 3548
rect 34196 3508 34197 3548
rect 34155 3499 34197 3508
rect 33963 3464 34005 3473
rect 33963 3424 33964 3464
rect 34004 3424 34005 3464
rect 33963 3415 34005 3424
rect 34156 3464 34196 3499
rect 33964 3330 34004 3415
rect 34156 3413 34196 3424
rect 34347 3464 34389 3473
rect 34347 3424 34348 3464
rect 34388 3424 34389 3464
rect 34347 3415 34389 3424
rect 34540 3464 34580 3473
rect 34348 3330 34388 3415
rect 34060 3212 34100 3221
rect 34443 3212 34485 3221
rect 34100 3172 34292 3212
rect 34060 3163 34100 3172
rect 34252 2540 34292 3172
rect 34443 3172 34444 3212
rect 34484 3172 34485 3212
rect 34443 3163 34485 3172
rect 34444 3078 34484 3163
rect 34540 2969 34580 3424
rect 34731 3464 34773 3473
rect 34731 3424 34732 3464
rect 34772 3424 34773 3464
rect 34731 3415 34773 3424
rect 34924 3464 34964 3473
rect 34732 3330 34772 3415
rect 34828 3212 34868 3221
rect 34539 2960 34581 2969
rect 34539 2920 34540 2960
rect 34580 2920 34581 2960
rect 34539 2911 34581 2920
rect 34060 2500 34292 2540
rect 33867 1280 33909 1289
rect 33867 1240 33868 1280
rect 33908 1240 33909 1280
rect 33867 1231 33909 1240
rect 33772 1112 33812 1121
rect 33772 869 33812 1072
rect 33963 1112 34005 1121
rect 33963 1072 33964 1112
rect 34004 1072 34005 1112
rect 33963 1063 34005 1072
rect 33964 978 34004 1063
rect 34060 1028 34100 2500
rect 34828 2465 34868 3172
rect 34924 2717 34964 3424
rect 35115 3464 35157 3473
rect 35115 3424 35116 3464
rect 35156 3424 35157 3464
rect 35115 3415 35157 3424
rect 35308 3464 35348 3473
rect 35116 3330 35156 3415
rect 35212 3212 35252 3221
rect 35212 2876 35252 3172
rect 35308 3053 35348 3424
rect 35499 3464 35541 3473
rect 35499 3424 35500 3464
rect 35540 3424 35541 3464
rect 35499 3415 35541 3424
rect 35692 3464 35732 3751
rect 37516 3473 37556 4012
rect 37804 4002 37844 4087
rect 37707 3968 37749 3977
rect 37707 3928 37708 3968
rect 37748 3928 37749 3968
rect 37707 3919 37749 3928
rect 37708 3800 37748 3919
rect 37708 3760 37844 3800
rect 35692 3415 35732 3424
rect 35883 3464 35925 3473
rect 35883 3424 35884 3464
rect 35924 3424 35925 3464
rect 35883 3415 35925 3424
rect 36076 3464 36116 3473
rect 35500 3330 35540 3415
rect 35884 3330 35924 3415
rect 36076 3389 36116 3424
rect 36267 3464 36309 3473
rect 36267 3424 36268 3464
rect 36308 3424 36309 3464
rect 36267 3415 36309 3424
rect 36460 3464 36500 3473
rect 36075 3380 36117 3389
rect 36075 3340 36076 3380
rect 36116 3340 36117 3380
rect 36075 3331 36117 3340
rect 35596 3212 35636 3221
rect 35980 3212 36020 3221
rect 35636 3172 35924 3212
rect 35596 3163 35636 3172
rect 35307 3044 35349 3053
rect 35307 3004 35308 3044
rect 35348 3004 35349 3044
rect 35307 2995 35349 3004
rect 35212 2836 35732 2876
rect 34923 2708 34965 2717
rect 34923 2668 34924 2708
rect 34964 2668 34965 2708
rect 34923 2659 34965 2668
rect 35692 2540 35732 2836
rect 35596 2500 35732 2540
rect 34827 2456 34869 2465
rect 34827 2416 34828 2456
rect 34868 2416 34869 2456
rect 34827 2407 34869 2416
rect 35307 2456 35349 2465
rect 35307 2416 35308 2456
rect 35348 2416 35349 2456
rect 35307 2407 35349 2416
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 35308 1457 35348 2407
rect 34923 1448 34965 1457
rect 34923 1408 34924 1448
rect 34964 1408 34965 1448
rect 34923 1399 34965 1408
rect 35307 1448 35349 1457
rect 35307 1408 35308 1448
rect 35348 1408 35349 1448
rect 35307 1399 35349 1408
rect 34443 1280 34485 1289
rect 34443 1240 34444 1280
rect 34484 1240 34485 1280
rect 34443 1231 34485 1240
rect 34156 1205 34196 1220
rect 34155 1196 34197 1205
rect 34155 1156 34156 1196
rect 34196 1156 34197 1196
rect 34155 1147 34197 1156
rect 34156 1125 34196 1147
rect 34156 1076 34196 1085
rect 34251 1113 34293 1121
rect 34348 1113 34388 1121
rect 34251 1112 34388 1113
rect 34251 1072 34252 1112
rect 34292 1073 34348 1112
rect 34292 1072 34293 1073
rect 34251 1063 34293 1072
rect 34348 1063 34388 1072
rect 34060 988 34196 1028
rect 33868 944 33908 953
rect 33771 860 33813 869
rect 33771 820 33772 860
rect 33812 820 33813 860
rect 33771 811 33813 820
rect 33676 652 33812 692
rect 33675 524 33717 533
rect 33675 484 33676 524
rect 33716 484 33717 524
rect 33675 475 33717 484
rect 33579 440 33621 449
rect 33579 400 33580 440
rect 33620 400 33621 440
rect 33579 391 33621 400
rect 33676 80 33716 475
rect 33772 356 33812 652
rect 33868 533 33908 904
rect 34156 617 34196 988
rect 34252 944 34292 953
rect 34155 608 34197 617
rect 34155 568 34156 608
rect 34196 568 34197 608
rect 34155 559 34197 568
rect 33867 524 33909 533
rect 33867 484 33868 524
rect 33908 484 33909 524
rect 33867 475 33909 484
rect 34252 449 34292 904
rect 34444 692 34484 1231
rect 34731 1196 34773 1205
rect 34731 1156 34732 1196
rect 34772 1156 34773 1196
rect 34731 1147 34773 1156
rect 34539 1112 34581 1121
rect 34539 1072 34540 1112
rect 34580 1072 34581 1112
rect 34539 1063 34581 1072
rect 34732 1112 34772 1147
rect 34540 978 34580 1063
rect 34732 1061 34772 1072
rect 34924 1112 34964 1399
rect 35116 1205 35156 1220
rect 35115 1196 35157 1205
rect 35115 1156 35116 1196
rect 35156 1156 35157 1196
rect 35115 1147 35157 1156
rect 35499 1196 35541 1205
rect 35499 1156 35500 1196
rect 35540 1156 35541 1196
rect 35499 1147 35541 1156
rect 35116 1125 35156 1147
rect 35116 1076 35156 1085
rect 35308 1113 35348 1121
rect 35403 1113 35445 1121
rect 35308 1112 35445 1113
rect 34924 1063 34964 1072
rect 35348 1073 35404 1112
rect 35348 1072 35355 1073
rect 35403 1072 35404 1073
rect 35444 1072 35445 1112
rect 35308 1063 35348 1072
rect 35403 1063 35445 1072
rect 35500 1112 35540 1147
rect 35500 1061 35540 1072
rect 34636 953 34676 1038
rect 35020 1028 35060 1037
rect 35060 988 35163 1028
rect 35020 979 35060 988
rect 34635 944 34677 953
rect 34635 904 34636 944
rect 34676 904 34677 944
rect 34635 895 34677 904
rect 35123 860 35163 988
rect 35211 944 35253 953
rect 35211 904 35212 944
rect 35252 904 35253 944
rect 35211 895 35253 904
rect 35403 944 35445 953
rect 35403 904 35404 944
rect 35444 904 35445 944
rect 35403 895 35445 904
rect 35116 820 35163 860
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 34348 652 34484 692
rect 34059 440 34101 449
rect 34059 400 34060 440
rect 34100 400 34101 440
rect 34059 391 34101 400
rect 34251 440 34293 449
rect 34251 400 34252 440
rect 34292 400 34293 440
rect 34251 391 34293 400
rect 33772 316 33908 356
rect 33868 80 33908 316
rect 34060 80 34100 391
rect 34348 272 34388 652
rect 34635 608 34677 617
rect 34635 568 34636 608
rect 34676 568 34677 608
rect 34635 559 34677 568
rect 34443 524 34485 533
rect 34443 484 34444 524
rect 34484 484 34485 524
rect 34443 475 34485 484
rect 34252 232 34388 272
rect 34252 80 34292 232
rect 34444 80 34484 475
rect 34636 80 34676 559
rect 34731 524 34773 533
rect 34731 484 34732 524
rect 34772 484 34773 524
rect 34731 475 34773 484
rect 34732 197 34772 475
rect 34827 440 34869 449
rect 34827 400 34828 440
rect 34868 400 34869 440
rect 34827 391 34869 400
rect 35019 440 35061 449
rect 35019 400 35020 440
rect 35060 400 35061 440
rect 35019 391 35061 400
rect 34731 188 34773 197
rect 34731 148 34732 188
rect 34772 148 34773 188
rect 34731 139 34773 148
rect 34828 80 34868 391
rect 35020 80 35060 391
rect 35116 197 35156 820
rect 35115 188 35157 197
rect 35115 148 35116 188
rect 35156 148 35157 188
rect 35115 139 35157 148
rect 35212 80 35252 895
rect 35404 810 35444 895
rect 35403 440 35445 449
rect 35403 400 35404 440
rect 35444 400 35445 440
rect 35403 391 35445 400
rect 35404 80 35444 391
rect 35596 356 35636 2500
rect 35691 2204 35733 2213
rect 35691 2164 35692 2204
rect 35732 2164 35733 2204
rect 35691 2155 35733 2164
rect 35692 1709 35732 2155
rect 35691 1700 35733 1709
rect 35691 1660 35692 1700
rect 35732 1660 35733 1700
rect 35691 1651 35733 1660
rect 35884 1448 35924 3172
rect 35980 1541 36020 3172
rect 36076 3053 36116 3331
rect 36268 3330 36308 3415
rect 36364 3212 36404 3221
rect 36075 3044 36117 3053
rect 36075 3004 36076 3044
rect 36116 3004 36117 3044
rect 36075 2995 36117 3004
rect 35979 1532 36021 1541
rect 35979 1492 35980 1532
rect 36020 1492 36021 1532
rect 35979 1483 36021 1492
rect 36364 1457 36404 3172
rect 36460 2885 36500 3424
rect 36651 3464 36693 3473
rect 36651 3424 36652 3464
rect 36692 3424 36693 3464
rect 36651 3415 36693 3424
rect 36843 3464 36885 3473
rect 36843 3424 36844 3464
rect 36884 3424 36885 3464
rect 36843 3415 36885 3424
rect 37515 3464 37557 3473
rect 37515 3424 37516 3464
rect 37556 3424 37557 3464
rect 37515 3415 37557 3424
rect 37707 3464 37749 3473
rect 37707 3424 37708 3464
rect 37748 3424 37749 3464
rect 37707 3415 37749 3424
rect 37804 3464 37844 3760
rect 37900 3464 37940 4096
rect 37996 4087 38036 4096
rect 38092 4061 38132 4180
rect 38091 4052 38133 4061
rect 38091 4012 38092 4052
rect 38132 4012 38133 4052
rect 38091 4003 38133 4012
rect 37996 3968 38036 3977
rect 37996 3809 38036 3928
rect 37995 3800 38037 3809
rect 37995 3760 37996 3800
rect 38036 3760 38037 3800
rect 37995 3751 38037 3760
rect 37996 3464 38036 3473
rect 37900 3424 37996 3464
rect 37804 3415 37844 3424
rect 37996 3415 38036 3424
rect 38092 3464 38132 3473
rect 38188 3464 38228 4339
rect 38380 4145 38420 4230
rect 38475 4220 38517 4229
rect 38475 4180 38476 4220
rect 38516 4180 38517 4220
rect 38475 4171 38517 4180
rect 38379 4136 38421 4145
rect 38379 4096 38380 4136
rect 38420 4096 38421 4136
rect 38379 4087 38421 4096
rect 38476 4136 38516 4171
rect 38476 4085 38516 4096
rect 38956 4061 38996 4423
rect 38955 4052 38997 4061
rect 38955 4012 38956 4052
rect 38996 4012 38997 4052
rect 38955 4003 38997 4012
rect 38379 3968 38421 3977
rect 38379 3928 38380 3968
rect 38420 3928 38421 3968
rect 38379 3919 38421 3928
rect 38380 3834 38420 3919
rect 38283 3716 38325 3725
rect 38283 3676 38284 3716
rect 38324 3676 38325 3716
rect 38283 3667 38325 3676
rect 38132 3424 38228 3464
rect 38284 3464 38324 3667
rect 40972 3641 41012 4684
rect 41164 4675 41204 4684
rect 41260 4556 41300 5440
rect 41451 5480 41493 5489
rect 41451 5440 41452 5480
rect 41492 5440 41493 5480
rect 41451 5431 41493 5440
rect 41452 5144 41492 5431
rect 41548 5237 41588 5524
rect 41547 5228 41589 5237
rect 41547 5188 41548 5228
rect 41588 5188 41589 5228
rect 41547 5179 41589 5188
rect 41452 5095 41492 5104
rect 41547 5060 41589 5069
rect 41547 5020 41548 5060
rect 41588 5020 41589 5060
rect 41547 5011 41589 5020
rect 41355 4976 41397 4985
rect 41355 4936 41356 4976
rect 41396 4936 41397 4976
rect 41355 4927 41397 4936
rect 41452 4976 41492 4985
rect 41356 4842 41396 4927
rect 41260 4516 41396 4556
rect 41259 4388 41301 4397
rect 41259 4348 41260 4388
rect 41300 4348 41301 4388
rect 41259 4339 41301 4348
rect 41260 4136 41300 4339
rect 41356 4136 41396 4516
rect 41452 4313 41492 4936
rect 41451 4304 41493 4313
rect 41451 4264 41452 4304
rect 41492 4264 41493 4304
rect 41451 4255 41493 4264
rect 41548 4178 41588 5011
rect 41644 4985 41684 6280
rect 41740 6271 41780 6280
rect 46732 6320 46772 6607
rect 47596 6488 47636 6607
rect 47596 6439 47636 6448
rect 47883 6488 47925 6497
rect 47883 6448 47884 6488
rect 47924 6448 47925 6488
rect 47883 6439 47925 6448
rect 48460 6488 48500 6607
rect 48556 6497 48596 6616
rect 49035 6656 49077 6665
rect 49035 6616 49036 6656
rect 49076 6616 49077 6656
rect 49035 6607 49077 6616
rect 48460 6439 48500 6448
rect 48555 6488 48597 6497
rect 48555 6448 48556 6488
rect 48596 6448 48597 6488
rect 48555 6439 48597 6448
rect 48747 6488 48789 6497
rect 48747 6448 48748 6488
rect 48788 6448 48789 6488
rect 48747 6439 48789 6448
rect 49036 6488 49076 6607
rect 49420 6497 49460 9940
rect 49804 9932 49844 9940
rect 49976 9932 50056 10000
rect 49804 9920 50056 9932
rect 60920 9920 61000 10000
rect 71864 9920 71944 10000
rect 82808 9920 82888 10000
rect 93752 9920 93832 10000
rect 49804 9892 50036 9920
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 49228 6488 49268 6497
rect 49076 6448 49228 6488
rect 49036 6439 49076 6448
rect 49228 6439 49268 6448
rect 49419 6488 49461 6497
rect 49419 6448 49420 6488
rect 49460 6448 49461 6488
rect 49419 6439 49461 6448
rect 47884 6354 47924 6439
rect 48748 6354 48788 6439
rect 48844 6404 48884 6413
rect 49324 6404 49364 6413
rect 48884 6364 48980 6404
rect 48844 6355 48884 6364
rect 46732 6271 46772 6280
rect 46827 6320 46869 6329
rect 46827 6280 46828 6320
rect 46868 6280 46869 6320
rect 46827 6271 46869 6280
rect 47596 6320 47636 6329
rect 44524 6236 44564 6245
rect 46060 6236 46100 6245
rect 44332 5657 44372 5742
rect 44524 5657 44564 6196
rect 45964 6196 46060 6236
rect 46100 6196 46292 6236
rect 41740 5648 41780 5657
rect 41740 5069 41780 5608
rect 41836 5648 41876 5657
rect 44236 5648 44276 5657
rect 41876 5608 41972 5648
rect 41836 5599 41876 5608
rect 41835 5480 41877 5489
rect 41835 5440 41836 5480
rect 41876 5440 41877 5480
rect 41835 5431 41877 5440
rect 41739 5060 41781 5069
rect 41739 5020 41740 5060
rect 41780 5020 41781 5060
rect 41739 5011 41781 5020
rect 41643 4976 41685 4985
rect 41643 4936 41644 4976
rect 41684 4936 41685 4976
rect 41643 4927 41685 4936
rect 41836 4892 41876 5431
rect 41740 4852 41876 4892
rect 41740 4397 41780 4852
rect 41836 4724 41876 4733
rect 41739 4388 41781 4397
rect 41451 4136 41493 4145
rect 41356 4096 41452 4136
rect 41492 4096 41493 4136
rect 41548 4129 41588 4138
rect 41644 4348 41740 4388
rect 41780 4348 41781 4388
rect 41260 4087 41300 4096
rect 41451 4087 41493 4096
rect 41452 4002 41492 4087
rect 41644 3977 41684 4348
rect 41739 4339 41781 4348
rect 41740 4052 41780 4061
rect 41259 3968 41301 3977
rect 41259 3928 41260 3968
rect 41300 3928 41301 3968
rect 41259 3919 41301 3928
rect 41643 3968 41685 3977
rect 41643 3928 41644 3968
rect 41684 3928 41685 3968
rect 41643 3919 41685 3928
rect 41260 3834 41300 3919
rect 41740 3725 41780 4012
rect 41739 3716 41781 3725
rect 41739 3676 41740 3716
rect 41780 3676 41781 3716
rect 41739 3667 41781 3676
rect 38379 3632 38421 3641
rect 38379 3592 38380 3632
rect 38420 3592 38421 3632
rect 38379 3583 38421 3592
rect 38571 3632 38613 3641
rect 38571 3592 38572 3632
rect 38612 3592 38613 3632
rect 38571 3583 38613 3592
rect 40971 3632 41013 3641
rect 40971 3592 40972 3632
rect 41012 3592 41013 3632
rect 38092 3415 38132 3424
rect 36652 3330 36692 3415
rect 36844 3330 36884 3415
rect 36748 3212 36788 3221
rect 36788 3172 37268 3212
rect 36748 3163 36788 3172
rect 36459 2876 36501 2885
rect 36459 2836 36460 2876
rect 36500 2836 36501 2876
rect 36459 2827 36501 2836
rect 36460 2297 36500 2827
rect 36459 2288 36501 2297
rect 36459 2248 36460 2288
rect 36500 2248 36501 2288
rect 36459 2239 36501 2248
rect 36747 1532 36789 1541
rect 36747 1492 36748 1532
rect 36788 1492 36789 1532
rect 36747 1483 36789 1492
rect 36363 1448 36405 1457
rect 35884 1408 35931 1448
rect 35891 1364 35931 1408
rect 36363 1408 36364 1448
rect 36404 1408 36405 1448
rect 36363 1399 36405 1408
rect 35891 1324 36020 1364
rect 35883 1196 35925 1205
rect 35883 1156 35884 1196
rect 35924 1156 35925 1196
rect 35883 1147 35925 1156
rect 35692 1112 35732 1121
rect 35692 869 35732 1072
rect 35884 1112 35924 1147
rect 35980 1121 36020 1324
rect 36267 1196 36309 1205
rect 36267 1156 36268 1196
rect 36308 1156 36309 1196
rect 36267 1147 36309 1156
rect 35884 1061 35924 1072
rect 35979 1112 36021 1121
rect 35979 1072 35980 1112
rect 36020 1072 36021 1112
rect 35979 1063 36021 1072
rect 36076 1112 36116 1121
rect 35788 944 35828 953
rect 35691 860 35733 869
rect 35691 820 35692 860
rect 35732 820 35733 860
rect 35691 811 35733 820
rect 35788 533 35828 904
rect 35979 944 36021 953
rect 35979 904 35980 944
rect 36020 904 36021 944
rect 35979 895 36021 904
rect 35787 524 35829 533
rect 35787 484 35788 524
rect 35828 484 35829 524
rect 35787 475 35829 484
rect 35596 316 35828 356
rect 35595 188 35637 197
rect 35595 148 35596 188
rect 35636 148 35637 188
rect 35595 139 35637 148
rect 35596 80 35636 139
rect 35788 80 35828 316
rect 35980 80 36020 895
rect 36076 365 36116 1072
rect 36268 1112 36308 1147
rect 36652 1121 36692 1206
rect 36268 1061 36308 1072
rect 36363 1112 36405 1121
rect 36363 1072 36364 1112
rect 36404 1072 36405 1112
rect 36363 1063 36405 1072
rect 36460 1112 36500 1121
rect 36171 944 36213 953
rect 36171 904 36172 944
rect 36212 904 36213 944
rect 36171 895 36213 904
rect 36172 810 36212 895
rect 36364 692 36404 1063
rect 36460 869 36500 1072
rect 36651 1112 36693 1121
rect 36651 1072 36652 1112
rect 36692 1072 36693 1112
rect 36651 1063 36693 1072
rect 36556 944 36596 953
rect 36748 944 36788 1483
rect 37131 1448 37173 1457
rect 37131 1408 37132 1448
rect 37172 1408 37173 1448
rect 37131 1399 37173 1408
rect 36843 1112 36885 1121
rect 36843 1072 36844 1112
rect 36884 1072 36885 1112
rect 36843 1063 36885 1072
rect 37035 1112 37077 1121
rect 37035 1072 37036 1112
rect 37076 1072 37077 1112
rect 37035 1063 37077 1072
rect 36844 978 36884 1063
rect 37036 978 37076 1063
rect 36459 860 36501 869
rect 36459 820 36460 860
rect 36500 820 36501 860
rect 36459 811 36501 820
rect 36172 652 36404 692
rect 36075 356 36117 365
rect 36075 316 36076 356
rect 36116 316 36117 356
rect 36075 307 36117 316
rect 36172 80 36212 652
rect 36556 533 36596 904
rect 36652 904 36788 944
rect 36940 944 36980 953
rect 36363 524 36405 533
rect 36363 484 36364 524
rect 36404 484 36405 524
rect 36363 475 36405 484
rect 36555 524 36597 533
rect 36555 484 36556 524
rect 36596 484 36597 524
rect 36555 475 36597 484
rect 36364 80 36404 475
rect 36652 356 36692 904
rect 36843 860 36885 869
rect 36843 820 36844 860
rect 36884 820 36885 860
rect 36843 811 36885 820
rect 36844 524 36884 811
rect 36556 316 36692 356
rect 36748 484 36884 524
rect 36556 80 36596 316
rect 36748 80 36788 484
rect 36940 449 36980 904
rect 37132 692 37172 1399
rect 37228 944 37268 3172
rect 37708 3044 37748 3415
rect 38284 3380 38324 3424
rect 38380 3389 38420 3583
rect 38475 3464 38517 3473
rect 38475 3424 38476 3464
rect 38516 3424 38517 3464
rect 38475 3415 38517 3424
rect 38188 3340 38324 3380
rect 38379 3380 38421 3389
rect 38379 3340 38380 3380
rect 38420 3340 38421 3380
rect 38188 3296 38228 3340
rect 38379 3331 38421 3340
rect 38476 3330 38516 3415
rect 38092 3256 38228 3296
rect 37804 3212 37844 3221
rect 37844 3172 37940 3212
rect 37804 3163 37844 3172
rect 37708 3004 37844 3044
rect 37612 2624 37652 2635
rect 37804 2633 37844 3004
rect 37612 2381 37652 2584
rect 37803 2624 37845 2633
rect 37803 2584 37804 2624
rect 37844 2584 37845 2624
rect 37803 2575 37845 2584
rect 37708 2540 37748 2549
rect 37611 2372 37653 2381
rect 37611 2332 37612 2372
rect 37652 2332 37653 2372
rect 37611 2323 37653 2332
rect 37612 1961 37652 2323
rect 37611 1952 37653 1961
rect 37611 1912 37612 1952
rect 37652 1912 37653 1952
rect 37611 1903 37653 1912
rect 37708 1280 37748 2500
rect 37803 1616 37845 1625
rect 37803 1576 37804 1616
rect 37844 1576 37845 1616
rect 37803 1567 37845 1576
rect 37612 1240 37748 1280
rect 37324 1121 37364 1206
rect 37323 1112 37365 1121
rect 37323 1072 37324 1112
rect 37364 1072 37365 1112
rect 37323 1063 37365 1072
rect 37515 1112 37557 1121
rect 37515 1072 37516 1112
rect 37556 1072 37557 1112
rect 37515 1063 37557 1072
rect 37516 978 37556 1063
rect 37419 944 37461 953
rect 37228 904 37364 944
rect 37036 652 37172 692
rect 36939 440 36981 449
rect 36939 400 36940 440
rect 36980 400 36981 440
rect 36939 391 36981 400
rect 37036 272 37076 652
rect 37131 524 37173 533
rect 37131 484 37132 524
rect 37172 484 37173 524
rect 37131 475 37173 484
rect 36940 232 37076 272
rect 36940 80 36980 232
rect 37132 80 37172 475
rect 37324 80 37364 904
rect 37419 904 37420 944
rect 37460 904 37461 944
rect 37612 944 37652 1240
rect 37804 1196 37844 1567
rect 37708 1156 37844 1196
rect 37708 1112 37748 1156
rect 37900 1121 37940 3172
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 37708 1063 37748 1072
rect 37899 1112 37941 1121
rect 37899 1072 37900 1112
rect 37940 1072 37941 1112
rect 37899 1063 37941 1072
rect 37804 944 37844 953
rect 37612 904 37748 944
rect 37419 895 37461 904
rect 37420 810 37460 895
rect 37515 440 37557 449
rect 37515 400 37516 440
rect 37556 400 37557 440
rect 37515 391 37557 400
rect 37516 80 37556 391
rect 37708 80 37748 904
rect 37804 533 37844 904
rect 37899 944 37941 953
rect 37899 904 37900 944
rect 37940 904 37941 944
rect 37996 944 38036 2827
rect 38092 2213 38132 3256
rect 38380 3212 38420 3221
rect 38380 3128 38420 3172
rect 38284 3088 38420 3128
rect 38284 2885 38324 3088
rect 38572 3044 38612 3583
rect 40492 3557 40532 3588
rect 40971 3583 41013 3592
rect 40491 3548 40533 3557
rect 40491 3508 40492 3548
rect 40532 3508 40533 3548
rect 40491 3499 40533 3508
rect 41355 3548 41397 3557
rect 41355 3508 41356 3548
rect 41396 3508 41397 3548
rect 41355 3499 41397 3508
rect 38859 3464 38901 3473
rect 38859 3424 38860 3464
rect 38900 3424 38901 3464
rect 38859 3415 38901 3424
rect 39052 3464 39092 3475
rect 38860 3330 38900 3415
rect 39052 3389 39092 3424
rect 39243 3464 39285 3473
rect 39243 3424 39244 3464
rect 39284 3424 39285 3464
rect 39243 3415 39285 3424
rect 39436 3464 39476 3473
rect 39051 3380 39093 3389
rect 39051 3340 39052 3380
rect 39092 3340 39093 3380
rect 39051 3331 39093 3340
rect 38380 3004 38612 3044
rect 38956 3212 38996 3221
rect 38283 2876 38325 2885
rect 38283 2836 38284 2876
rect 38324 2836 38325 2876
rect 38283 2827 38325 2836
rect 38188 2611 38228 2635
rect 38188 2549 38228 2571
rect 38380 2624 38420 3004
rect 38572 2633 38612 2718
rect 38764 2633 38804 2718
rect 38187 2540 38229 2549
rect 38187 2500 38188 2540
rect 38228 2500 38229 2540
rect 38187 2491 38229 2500
rect 38284 2540 38324 2549
rect 38091 2204 38133 2213
rect 38091 2164 38092 2204
rect 38132 2164 38133 2204
rect 38091 2155 38133 2164
rect 38091 1364 38133 1373
rect 38091 1324 38092 1364
rect 38132 1324 38133 1364
rect 38091 1315 38133 1324
rect 38092 1112 38132 1315
rect 38284 1280 38324 2500
rect 38380 2129 38420 2584
rect 38571 2624 38613 2633
rect 38571 2584 38572 2624
rect 38612 2584 38613 2624
rect 38571 2575 38613 2584
rect 38763 2624 38805 2633
rect 38763 2584 38764 2624
rect 38804 2584 38805 2624
rect 38763 2575 38805 2584
rect 38668 2540 38708 2549
rect 38379 2120 38421 2129
rect 38379 2080 38380 2120
rect 38420 2080 38421 2120
rect 38379 2071 38421 2080
rect 38668 1364 38708 2500
rect 38668 1324 38804 1364
rect 38284 1240 38420 1280
rect 38092 1063 38132 1072
rect 38283 1112 38325 1121
rect 38283 1072 38284 1112
rect 38324 1072 38325 1112
rect 38283 1063 38325 1072
rect 38284 978 38324 1063
rect 38187 944 38229 953
rect 37996 904 38132 944
rect 37899 895 37941 904
rect 37803 524 37845 533
rect 37803 484 37804 524
rect 37844 484 37845 524
rect 37803 475 37845 484
rect 37900 80 37940 895
rect 38092 80 38132 904
rect 38187 904 38188 944
rect 38228 904 38229 944
rect 38187 895 38229 904
rect 38188 810 38228 895
rect 38380 860 38420 1240
rect 38476 1205 38516 1207
rect 38475 1196 38517 1205
rect 38475 1156 38476 1196
rect 38516 1156 38517 1196
rect 38475 1147 38517 1156
rect 38476 1112 38516 1147
rect 38668 1121 38708 1206
rect 38476 1063 38516 1072
rect 38667 1112 38709 1121
rect 38667 1072 38668 1112
rect 38708 1072 38709 1112
rect 38667 1063 38709 1072
rect 38572 944 38612 953
rect 38380 820 38516 860
rect 38283 524 38325 533
rect 38283 484 38284 524
rect 38324 484 38325 524
rect 38283 475 38325 484
rect 38284 80 38324 475
rect 38476 80 38516 820
rect 38572 533 38612 904
rect 38667 944 38709 953
rect 38667 904 38668 944
rect 38708 904 38709 944
rect 38764 944 38804 1324
rect 38956 1280 38996 3172
rect 39052 1793 39092 3331
rect 39244 3330 39284 3415
rect 39436 3305 39476 3424
rect 39627 3464 39669 3473
rect 39627 3424 39628 3464
rect 39668 3424 39669 3464
rect 39627 3415 39669 3424
rect 39820 3464 39860 3473
rect 39628 3330 39668 3415
rect 39435 3296 39477 3305
rect 39435 3256 39436 3296
rect 39476 3256 39477 3296
rect 39435 3247 39477 3256
rect 39340 3212 39380 3221
rect 39340 2540 39380 3172
rect 39436 3137 39476 3247
rect 39820 3221 39860 3424
rect 40011 3464 40053 3473
rect 40011 3424 40012 3464
rect 40052 3424 40053 3464
rect 40011 3415 40053 3424
rect 40299 3464 40341 3473
rect 40299 3424 40300 3464
rect 40340 3424 40341 3464
rect 40299 3415 40341 3424
rect 40492 3464 40532 3499
rect 39724 3212 39764 3221
rect 39435 3128 39477 3137
rect 39435 3088 39436 3128
rect 39476 3088 39477 3128
rect 39435 3079 39477 3088
rect 39724 2540 39764 3172
rect 39819 3212 39861 3221
rect 39819 3172 39820 3212
rect 39860 3172 39861 3212
rect 39819 3163 39861 3172
rect 40012 2624 40052 3415
rect 40300 3330 40340 3415
rect 40492 3305 40532 3424
rect 40779 3464 40821 3473
rect 40779 3424 40780 3464
rect 40820 3424 40821 3464
rect 40779 3415 40821 3424
rect 40972 3464 41012 3473
rect 40780 3330 40820 3415
rect 40491 3296 40533 3305
rect 40491 3256 40492 3296
rect 40532 3256 40533 3296
rect 40491 3247 40533 3256
rect 40396 3212 40436 3221
rect 40204 2633 40244 2718
rect 40012 2575 40052 2584
rect 40203 2624 40245 2633
rect 40203 2584 40204 2624
rect 40244 2584 40245 2624
rect 40203 2575 40245 2584
rect 40108 2540 40148 2549
rect 39340 2500 39572 2540
rect 39724 2500 39956 2540
rect 39051 1784 39093 1793
rect 39051 1744 39052 1784
rect 39092 1744 39093 1784
rect 39051 1735 39093 1744
rect 38956 1240 39188 1280
rect 38859 1196 38901 1205
rect 38859 1156 38860 1196
rect 38900 1156 38901 1196
rect 38859 1147 38901 1156
rect 38860 1112 38900 1147
rect 38860 1061 38900 1072
rect 39051 1112 39093 1121
rect 39051 1072 39052 1112
rect 39092 1072 39093 1112
rect 39051 1063 39093 1072
rect 39052 978 39092 1063
rect 38955 944 38997 953
rect 38764 904 38900 944
rect 38667 895 38709 904
rect 38571 524 38613 533
rect 38571 484 38572 524
rect 38612 484 38613 524
rect 38571 475 38613 484
rect 38668 80 38708 895
rect 38860 80 38900 904
rect 38955 904 38956 944
rect 38996 904 38997 944
rect 39148 944 39188 1240
rect 39243 1196 39285 1205
rect 39243 1156 39244 1196
rect 39284 1156 39285 1196
rect 39243 1147 39285 1156
rect 39244 1112 39284 1147
rect 39436 1121 39476 1206
rect 39244 1061 39284 1072
rect 39435 1112 39477 1121
rect 39435 1072 39436 1112
rect 39476 1072 39477 1112
rect 39435 1063 39477 1072
rect 39340 944 39380 953
rect 39148 904 39284 944
rect 38955 895 38997 904
rect 38956 810 38996 895
rect 39051 524 39093 533
rect 39051 484 39052 524
rect 39092 484 39093 524
rect 39051 475 39093 484
rect 39052 80 39092 475
rect 39244 80 39284 904
rect 39340 449 39380 904
rect 39435 944 39477 953
rect 39435 904 39436 944
rect 39476 904 39477 944
rect 39532 944 39572 2500
rect 39627 1280 39669 1289
rect 39627 1240 39628 1280
rect 39668 1240 39669 1280
rect 39627 1231 39669 1240
rect 39628 1112 39668 1231
rect 39628 1063 39668 1072
rect 39819 1112 39861 1121
rect 39819 1072 39820 1112
rect 39860 1072 39861 1112
rect 39819 1063 39861 1072
rect 39820 978 39860 1063
rect 39723 944 39765 953
rect 39532 904 39668 944
rect 39435 895 39477 904
rect 39339 440 39381 449
rect 39339 400 39340 440
rect 39380 400 39381 440
rect 39339 391 39381 400
rect 39436 80 39476 895
rect 39628 80 39668 904
rect 39723 904 39724 944
rect 39764 904 39765 944
rect 39916 944 39956 2500
rect 40396 2540 40436 3172
rect 40876 3212 40916 3221
rect 40876 2540 40916 3172
rect 40972 2969 41012 3424
rect 41163 3464 41205 3473
rect 41163 3424 41164 3464
rect 41204 3424 41205 3464
rect 41163 3415 41205 3424
rect 41356 3464 41396 3499
rect 41164 3330 41204 3415
rect 41260 3212 41300 3221
rect 40971 2960 41013 2969
rect 40971 2920 40972 2960
rect 41012 2920 41013 2960
rect 40971 2911 41013 2920
rect 40972 2801 41012 2911
rect 40971 2792 41013 2801
rect 40971 2752 40972 2792
rect 41012 2752 41013 2792
rect 40971 2743 41013 2752
rect 40396 2500 40724 2540
rect 40876 2500 41108 2540
rect 40108 1364 40148 2500
rect 40108 1324 40340 1364
rect 40011 1196 40053 1205
rect 40011 1156 40012 1196
rect 40052 1156 40053 1196
rect 40011 1147 40053 1156
rect 40012 1112 40052 1147
rect 40204 1121 40244 1206
rect 40012 1061 40052 1072
rect 40203 1112 40245 1121
rect 40203 1072 40204 1112
rect 40244 1072 40245 1112
rect 40203 1063 40245 1072
rect 40108 944 40148 953
rect 39916 904 40052 944
rect 39723 895 39765 904
rect 39724 810 39764 895
rect 39819 440 39861 449
rect 39819 400 39820 440
rect 39860 400 39861 440
rect 39819 391 39861 400
rect 39820 80 39860 391
rect 40012 80 40052 904
rect 40108 533 40148 904
rect 40203 944 40245 953
rect 40203 904 40204 944
rect 40244 904 40245 944
rect 40300 944 40340 1324
rect 40395 1196 40437 1205
rect 40395 1156 40396 1196
rect 40436 1156 40437 1196
rect 40395 1147 40437 1156
rect 40396 1112 40436 1147
rect 40396 1061 40436 1072
rect 40587 1112 40629 1121
rect 40587 1072 40588 1112
rect 40628 1072 40629 1112
rect 40587 1063 40629 1072
rect 40588 978 40628 1063
rect 40491 944 40533 953
rect 40300 904 40436 944
rect 40203 895 40245 904
rect 40107 524 40149 533
rect 40107 484 40108 524
rect 40148 484 40149 524
rect 40107 475 40149 484
rect 40204 80 40244 895
rect 40396 80 40436 904
rect 40491 904 40492 944
rect 40532 904 40533 944
rect 40684 944 40724 2500
rect 40780 1121 40820 1206
rect 40972 1205 41012 1207
rect 40971 1196 41013 1205
rect 40971 1156 40972 1196
rect 41012 1156 41013 1196
rect 40971 1147 41013 1156
rect 40779 1112 40821 1121
rect 40779 1072 40780 1112
rect 40820 1072 40821 1112
rect 40779 1063 40821 1072
rect 40972 1112 41012 1147
rect 40972 1063 41012 1072
rect 40876 944 40916 953
rect 40684 904 40820 944
rect 40491 895 40533 904
rect 40492 810 40532 895
rect 40587 524 40629 533
rect 40587 484 40588 524
rect 40628 484 40629 524
rect 40587 475 40629 484
rect 40588 80 40628 475
rect 40780 80 40820 904
rect 40876 533 40916 904
rect 40971 944 41013 953
rect 40971 904 40972 944
rect 41012 904 41013 944
rect 41068 944 41108 2500
rect 41260 1700 41300 3172
rect 41356 2717 41396 3424
rect 41643 3464 41685 3473
rect 41643 3424 41644 3464
rect 41684 3424 41685 3464
rect 41643 3415 41685 3424
rect 41644 2717 41684 3415
rect 41836 3221 41876 4684
rect 41932 4397 41972 5608
rect 44044 5564 44084 5573
rect 42123 5480 42165 5489
rect 42123 5440 42124 5480
rect 42164 5440 42165 5480
rect 42123 5431 42165 5440
rect 42124 5144 42164 5431
rect 42124 5095 42164 5104
rect 42027 5060 42069 5069
rect 42027 5020 42028 5060
rect 42068 5020 42069 5060
rect 42027 5011 42069 5020
rect 42699 5060 42741 5069
rect 42699 5020 42700 5060
rect 42740 5020 42741 5060
rect 42699 5011 42741 5020
rect 42028 4976 42068 5011
rect 42028 4925 42068 4936
rect 42123 4976 42165 4985
rect 42123 4936 42124 4976
rect 42164 4936 42165 4976
rect 42123 4927 42165 4936
rect 41931 4388 41973 4397
rect 41931 4348 41932 4388
rect 41972 4348 41973 4388
rect 41931 4339 41973 4348
rect 41932 4145 41972 4339
rect 42124 4313 42164 4927
rect 42123 4304 42165 4313
rect 42123 4264 42124 4304
rect 42164 4264 42165 4304
rect 42123 4255 42165 4264
rect 42603 4304 42645 4313
rect 42603 4264 42604 4304
rect 42644 4264 42645 4304
rect 42603 4255 42645 4264
rect 42027 4220 42069 4229
rect 42027 4180 42028 4220
rect 42068 4180 42069 4220
rect 42027 4171 42069 4180
rect 42316 4180 42452 4220
rect 41931 4136 41973 4145
rect 41931 4096 41932 4136
rect 41972 4096 41973 4136
rect 41931 4087 41973 4096
rect 42028 4136 42068 4171
rect 41932 4002 41972 4087
rect 42028 4085 42068 4096
rect 42316 3977 42356 4180
rect 42412 4136 42452 4180
rect 42412 4087 42452 4096
rect 42604 4136 42644 4255
rect 42604 4087 42644 4096
rect 42700 4136 42740 5011
rect 43947 4556 43989 4565
rect 43947 4516 43948 4556
rect 43988 4516 43989 4556
rect 43947 4507 43989 4516
rect 42795 4388 42837 4397
rect 42795 4348 42796 4388
rect 42836 4348 42837 4388
rect 42795 4339 42837 4348
rect 43084 4388 43124 4397
rect 43124 4348 43412 4388
rect 43084 4339 43124 4348
rect 42700 4087 42740 4096
rect 42507 4052 42549 4061
rect 42507 4012 42508 4052
rect 42548 4012 42549 4052
rect 42507 4003 42549 4012
rect 42027 3968 42069 3977
rect 42027 3928 42028 3968
rect 42068 3928 42069 3968
rect 42027 3919 42069 3928
rect 42315 3968 42357 3977
rect 42315 3928 42316 3968
rect 42356 3928 42357 3968
rect 42315 3919 42357 3928
rect 42412 3968 42452 3977
rect 42028 3834 42068 3919
rect 41931 3464 41973 3473
rect 41931 3424 41932 3464
rect 41972 3424 41973 3464
rect 41931 3415 41973 3424
rect 42124 3464 42164 3473
rect 41932 3330 41972 3415
rect 42124 3389 42164 3424
rect 42316 3464 42356 3919
rect 42316 3415 42356 3424
rect 42123 3380 42165 3389
rect 42123 3340 42124 3380
rect 42164 3340 42165 3380
rect 42123 3331 42165 3340
rect 41835 3212 41877 3221
rect 41835 3172 41836 3212
rect 41876 3172 41877 3212
rect 41835 3163 41877 3172
rect 42027 3212 42069 3221
rect 42027 3172 42028 3212
rect 42068 3172 42069 3212
rect 42027 3163 42069 3172
rect 41836 2969 41876 3163
rect 42028 3078 42068 3163
rect 42124 3137 42164 3331
rect 42316 3212 42356 3221
rect 42123 3128 42165 3137
rect 42123 3088 42124 3128
rect 42164 3088 42165 3128
rect 42123 3079 42165 3088
rect 41835 2960 41877 2969
rect 41835 2920 41836 2960
rect 41876 2920 41877 2960
rect 41835 2911 41877 2920
rect 41355 2708 41397 2717
rect 41355 2668 41356 2708
rect 41396 2668 41397 2708
rect 41355 2659 41397 2668
rect 41643 2708 41685 2717
rect 41643 2668 41644 2708
rect 41684 2668 41685 2708
rect 41643 2659 41685 2668
rect 41644 2624 41684 2659
rect 41836 2633 41876 2718
rect 42027 2708 42069 2717
rect 42027 2668 42028 2708
rect 42068 2668 42069 2708
rect 42027 2659 42069 2668
rect 41644 2574 41684 2584
rect 41835 2624 41877 2633
rect 41835 2584 41836 2624
rect 41876 2584 41877 2624
rect 41835 2575 41877 2584
rect 42028 2624 42068 2659
rect 42220 2633 42260 2718
rect 42028 2573 42068 2584
rect 42219 2624 42261 2633
rect 42219 2584 42220 2624
rect 42260 2584 42261 2624
rect 42219 2575 42261 2584
rect 42316 2549 42356 3172
rect 41739 2540 41781 2549
rect 41739 2500 41740 2540
rect 41780 2500 41781 2540
rect 41739 2491 41781 2500
rect 42124 2540 42164 2549
rect 41740 2406 41780 2491
rect 42027 2456 42069 2465
rect 42027 2416 42028 2456
rect 42068 2416 42069 2456
rect 42027 2407 42069 2416
rect 41260 1660 41492 1700
rect 41164 1121 41204 1206
rect 41163 1112 41205 1121
rect 41163 1072 41164 1112
rect 41204 1072 41205 1112
rect 41163 1063 41205 1072
rect 41355 1112 41397 1121
rect 41355 1072 41356 1112
rect 41396 1072 41397 1112
rect 41355 1063 41397 1072
rect 41356 978 41396 1063
rect 41259 944 41301 953
rect 41068 904 41204 944
rect 40971 895 41013 904
rect 40875 524 40917 533
rect 40875 484 40876 524
rect 40916 484 40917 524
rect 40875 475 40917 484
rect 40972 80 41012 895
rect 41164 80 41204 904
rect 41259 904 41260 944
rect 41300 904 41301 944
rect 41259 895 41301 904
rect 41260 810 41300 895
rect 41452 860 41492 1660
rect 42028 1289 42068 2407
rect 42124 1364 42164 2500
rect 42315 2540 42357 2549
rect 42315 2500 42316 2540
rect 42356 2500 42357 2540
rect 42315 2491 42357 2500
rect 42412 2465 42452 3928
rect 42508 3464 42548 4003
rect 42796 3884 42836 4339
rect 43179 4220 43221 4229
rect 43179 4180 43180 4220
rect 43220 4180 43221 4220
rect 43179 4171 43221 4180
rect 42892 4136 42932 4145
rect 42892 3977 42932 4096
rect 43084 4136 43124 4147
rect 43084 4061 43124 4096
rect 43180 4136 43220 4171
rect 43180 4085 43220 4096
rect 43083 4052 43125 4061
rect 43083 4012 43084 4052
rect 43124 4012 43125 4052
rect 43083 4003 43125 4012
rect 42891 3968 42933 3977
rect 42891 3928 42892 3968
rect 42932 3928 42933 3968
rect 42891 3919 42933 3928
rect 42508 3415 42548 3424
rect 42604 3844 42836 3884
rect 42604 3464 42644 3844
rect 42604 3415 42644 3424
rect 42796 3464 42836 3473
rect 42603 3212 42645 3221
rect 42603 3172 42604 3212
rect 42644 3172 42645 3212
rect 42603 3163 42645 3172
rect 42411 2456 42453 2465
rect 42411 2416 42412 2456
rect 42452 2416 42453 2456
rect 42411 2407 42453 2416
rect 42124 1324 42260 1364
rect 42027 1280 42069 1289
rect 42027 1240 42028 1280
rect 42068 1240 42069 1280
rect 42027 1231 42069 1240
rect 41740 1121 41780 1206
rect 41547 1112 41589 1121
rect 41547 1072 41548 1112
rect 41588 1072 41589 1112
rect 41547 1063 41589 1072
rect 41739 1112 41781 1121
rect 41739 1072 41740 1112
rect 41780 1072 41781 1112
rect 41739 1063 41781 1072
rect 41943 1101 41983 1123
rect 42028 1121 42068 1231
rect 42123 1196 42165 1205
rect 42123 1156 42124 1196
rect 42164 1156 42165 1196
rect 42123 1147 42165 1156
rect 41548 978 41588 1063
rect 42027 1112 42069 1121
rect 42027 1072 42028 1112
rect 42068 1072 42069 1112
rect 42027 1063 42069 1072
rect 42124 1112 42164 1147
rect 42124 1061 42164 1072
rect 41943 1037 41983 1061
rect 41942 1028 41984 1037
rect 41942 988 41943 1028
rect 41983 988 41984 1028
rect 41942 979 41984 988
rect 41644 944 41684 953
rect 41452 820 41588 860
rect 41355 524 41397 533
rect 41355 484 41356 524
rect 41396 484 41397 524
rect 41355 475 41397 484
rect 41356 80 41396 475
rect 41548 80 41588 820
rect 41644 449 41684 904
rect 41739 944 41781 953
rect 41739 904 41740 944
rect 41780 904 41781 944
rect 41739 895 41781 904
rect 42027 944 42069 953
rect 42027 904 42028 944
rect 42068 904 42069 944
rect 42220 944 42260 1324
rect 42315 1280 42357 1289
rect 42315 1240 42316 1280
rect 42356 1240 42357 1280
rect 42315 1231 42357 1240
rect 42316 1121 42356 1231
rect 42508 1205 42548 1207
rect 42507 1196 42549 1205
rect 42507 1156 42508 1196
rect 42548 1156 42549 1196
rect 42507 1147 42549 1156
rect 42315 1112 42357 1121
rect 42315 1072 42316 1112
rect 42356 1072 42357 1112
rect 42315 1063 42357 1072
rect 42508 1112 42548 1147
rect 42508 1063 42548 1072
rect 42412 944 42452 953
rect 42220 904 42351 944
rect 42027 895 42069 904
rect 41643 440 41685 449
rect 41643 400 41644 440
rect 41684 400 41685 440
rect 41643 391 41685 400
rect 41740 80 41780 895
rect 42028 810 42068 895
rect 42311 776 42351 904
rect 42311 736 42356 776
rect 41931 608 41973 617
rect 41931 568 41932 608
rect 41972 568 41973 608
rect 41931 559 41973 568
rect 41932 80 41972 559
rect 42123 440 42165 449
rect 42123 400 42124 440
rect 42164 400 42165 440
rect 42123 391 42165 400
rect 42124 80 42164 391
rect 42316 80 42356 736
rect 42412 449 42452 904
rect 42507 944 42549 953
rect 42507 904 42508 944
rect 42548 904 42549 944
rect 42604 944 42644 3163
rect 42796 2717 42836 3424
rect 42988 3464 43028 3473
rect 43028 3424 43220 3464
rect 42988 3415 43028 3424
rect 43180 3221 43220 3424
rect 42892 3212 42932 3221
rect 43179 3212 43221 3221
rect 42932 3172 43124 3212
rect 42892 3163 42932 3172
rect 42795 2708 42837 2717
rect 42795 2668 42796 2708
rect 42836 2668 42837 2708
rect 42795 2659 42837 2668
rect 42796 2624 42836 2659
rect 42988 2633 43028 2718
rect 42796 2573 42836 2584
rect 42987 2624 43029 2633
rect 42987 2584 42988 2624
rect 43028 2584 43029 2624
rect 42987 2575 43029 2584
rect 42892 2540 42932 2549
rect 42892 2045 42932 2500
rect 42891 2036 42933 2045
rect 42891 1996 42892 2036
rect 42932 1996 42933 2036
rect 42891 1987 42933 1996
rect 43084 1364 43124 3172
rect 43179 3172 43180 3212
rect 43220 3172 43221 3212
rect 43179 3163 43221 3172
rect 43180 2297 43220 3163
rect 43179 2288 43221 2297
rect 43179 2248 43180 2288
rect 43220 2248 43221 2288
rect 43179 2239 43221 2248
rect 43372 1373 43412 4348
rect 43563 3800 43605 3809
rect 43563 3760 43564 3800
rect 43604 3760 43605 3800
rect 43563 3751 43605 3760
rect 43467 2036 43509 2045
rect 43467 1996 43468 2036
rect 43508 1996 43509 2036
rect 43467 1987 43509 1996
rect 42988 1324 43124 1364
rect 43371 1364 43413 1373
rect 43371 1324 43372 1364
rect 43412 1324 43413 1364
rect 42699 1196 42741 1205
rect 42699 1156 42700 1196
rect 42740 1156 42741 1196
rect 42699 1147 42741 1156
rect 42700 1112 42740 1147
rect 42700 1061 42740 1072
rect 42891 1112 42933 1121
rect 42891 1072 42892 1112
rect 42932 1072 42933 1112
rect 42891 1063 42933 1072
rect 42892 978 42932 1063
rect 42795 944 42837 953
rect 42604 904 42740 944
rect 42507 895 42549 904
rect 42411 440 42453 449
rect 42411 400 42412 440
rect 42452 400 42453 440
rect 42411 391 42453 400
rect 42508 80 42548 895
rect 42700 80 42740 904
rect 42795 904 42796 944
rect 42836 904 42837 944
rect 42988 944 43028 1324
rect 43371 1315 43413 1324
rect 43084 1121 43124 1206
rect 43276 1121 43316 1206
rect 43372 1205 43412 1315
rect 43371 1196 43413 1205
rect 43371 1156 43372 1196
rect 43412 1156 43413 1196
rect 43371 1147 43413 1156
rect 43083 1112 43125 1121
rect 43083 1072 43084 1112
rect 43124 1072 43125 1112
rect 43083 1063 43125 1072
rect 43275 1112 43317 1121
rect 43275 1072 43276 1112
rect 43316 1072 43317 1112
rect 43275 1063 43317 1072
rect 43180 944 43220 953
rect 42988 904 43124 944
rect 42795 895 42837 904
rect 42796 810 42836 895
rect 42891 440 42933 449
rect 42891 400 42892 440
rect 42932 400 42933 440
rect 42891 391 42933 400
rect 42892 80 42932 391
rect 43084 80 43124 904
rect 43180 365 43220 904
rect 43275 944 43317 953
rect 43275 904 43276 944
rect 43316 904 43317 944
rect 43275 895 43317 904
rect 43179 356 43221 365
rect 43179 316 43180 356
rect 43220 316 43221 356
rect 43179 307 43221 316
rect 43276 80 43316 895
rect 43468 80 43508 1987
rect 43564 1280 43604 3751
rect 43948 3557 43988 4507
rect 43947 3548 43989 3557
rect 43947 3508 43948 3548
rect 43988 3508 43989 3548
rect 43947 3499 43989 3508
rect 43948 2624 43988 3499
rect 44044 2885 44084 5524
rect 44236 4229 44276 5608
rect 44331 5648 44373 5657
rect 44331 5608 44332 5648
rect 44372 5608 44373 5648
rect 44331 5599 44373 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44908 5648 44948 5659
rect 45004 5657 45044 5742
rect 44908 5573 44948 5608
rect 45003 5648 45045 5657
rect 45003 5608 45004 5648
rect 45044 5608 45140 5648
rect 45003 5599 45045 5608
rect 44619 5564 44661 5573
rect 44619 5524 44620 5564
rect 44660 5524 44661 5564
rect 44619 5515 44661 5524
rect 44716 5564 44756 5573
rect 44332 5480 44372 5489
rect 44332 5153 44372 5440
rect 44331 5144 44373 5153
rect 44331 5104 44332 5144
rect 44372 5104 44373 5144
rect 44331 5095 44373 5104
rect 44235 4220 44277 4229
rect 44235 4180 44236 4220
rect 44276 4180 44277 4220
rect 44235 4171 44277 4180
rect 44332 4145 44372 5095
rect 44620 5069 44660 5515
rect 44619 5060 44661 5069
rect 44619 5020 44620 5060
rect 44660 5020 44661 5060
rect 44619 5011 44661 5020
rect 44620 4178 44660 5011
rect 44331 4136 44373 4145
rect 44331 4096 44332 4136
rect 44372 4096 44373 4136
rect 44331 4087 44373 4096
rect 44428 4136 44564 4151
rect 44428 4111 44524 4136
rect 44428 4061 44468 4111
rect 44620 4129 44660 4138
rect 44524 4087 44564 4096
rect 44427 4052 44469 4061
rect 44716 4052 44756 5524
rect 44907 5564 44949 5573
rect 44907 5524 44908 5564
rect 44948 5524 44949 5564
rect 44907 5515 44949 5524
rect 45004 5480 45044 5489
rect 45004 5153 45044 5440
rect 44811 5144 44853 5153
rect 44811 5104 44812 5144
rect 44852 5104 44853 5144
rect 44811 5095 44853 5104
rect 45003 5144 45045 5153
rect 45003 5104 45004 5144
rect 45044 5104 45045 5144
rect 45003 5095 45045 5104
rect 44812 4136 44852 5095
rect 45100 4976 45140 5608
rect 45868 5153 45908 5238
rect 45867 5144 45909 5153
rect 45867 5104 45868 5144
rect 45908 5104 45909 5144
rect 45867 5095 45909 5104
rect 44812 4087 44852 4096
rect 45004 4936 45140 4976
rect 45868 4976 45908 4987
rect 45964 4985 46004 6196
rect 46060 6187 46100 6196
rect 46060 5648 46100 5657
rect 46252 5648 46292 6196
rect 46828 6186 46868 6271
rect 46100 5608 46196 5648
rect 46060 5599 46100 5608
rect 46060 5480 46100 5489
rect 45004 4136 45044 4936
rect 45868 4901 45908 4936
rect 45963 4976 46005 4985
rect 45963 4936 45964 4976
rect 46004 4936 46005 4976
rect 45963 4927 46005 4936
rect 45867 4892 45909 4901
rect 45867 4852 45868 4892
rect 45908 4852 45909 4892
rect 45867 4843 45909 4852
rect 45964 4842 46004 4927
rect 46060 4388 46100 5440
rect 46156 5153 46196 5608
rect 46252 5599 46292 5608
rect 46348 5648 46388 5659
rect 46348 5573 46388 5608
rect 47596 5573 47636 6280
rect 48268 6320 48308 6329
rect 46347 5564 46389 5573
rect 46347 5524 46348 5564
rect 46388 5524 46389 5564
rect 46347 5515 46389 5524
rect 46539 5564 46581 5573
rect 46539 5524 46540 5564
rect 46580 5524 46581 5564
rect 46539 5515 46581 5524
rect 47595 5564 47637 5573
rect 47595 5524 47596 5564
rect 47636 5524 47637 5564
rect 47595 5515 47637 5524
rect 46155 5144 46197 5153
rect 46155 5104 46156 5144
rect 46196 5104 46197 5144
rect 46155 5095 46197 5104
rect 46540 4976 46580 5515
rect 46636 5153 46676 5238
rect 48076 5153 48116 5238
rect 46635 5144 46677 5153
rect 48075 5144 48117 5153
rect 46635 5104 46636 5144
rect 46676 5104 46677 5144
rect 46635 5095 46677 5104
rect 47980 5104 48076 5144
rect 48116 5104 48117 5144
rect 46540 4927 46580 4936
rect 46635 4976 46677 4985
rect 46635 4936 46636 4976
rect 46676 4936 46677 4976
rect 46635 4927 46677 4936
rect 46251 4892 46293 4901
rect 46251 4852 46252 4892
rect 46292 4852 46293 4892
rect 46251 4843 46293 4852
rect 45868 4348 46100 4388
rect 46156 4724 46196 4733
rect 45099 4220 45141 4229
rect 45099 4180 45100 4220
rect 45140 4180 45141 4220
rect 45099 4171 45141 4180
rect 45004 4061 45044 4096
rect 45100 4136 45140 4171
rect 45100 4085 45140 4096
rect 44427 4012 44428 4052
rect 44468 4012 44469 4052
rect 44427 4003 44469 4012
rect 44620 4012 44756 4052
rect 45003 4052 45045 4061
rect 45003 4012 45004 4052
rect 45044 4012 45045 4052
rect 44332 3968 44372 3977
rect 44235 3716 44277 3725
rect 44235 3676 44236 3716
rect 44276 3676 44277 3716
rect 44235 3667 44277 3676
rect 44043 2876 44085 2885
rect 44043 2836 44044 2876
rect 44084 2836 44085 2876
rect 44043 2827 44085 2836
rect 44044 2624 44084 2633
rect 43948 2584 44044 2624
rect 43948 2540 43988 2584
rect 44044 2575 44084 2584
rect 44236 2624 44276 3667
rect 43660 2500 43988 2540
rect 44140 2540 44180 2549
rect 43660 1952 43700 2500
rect 43660 1903 43700 1912
rect 43851 1952 43893 1961
rect 43851 1912 43852 1952
rect 43892 1912 43893 1952
rect 43851 1903 43893 1912
rect 43852 1818 43892 1903
rect 43756 1700 43796 1709
rect 43796 1660 43892 1700
rect 43756 1651 43796 1660
rect 43564 1240 43796 1280
rect 43756 1121 43796 1240
rect 43563 1112 43605 1121
rect 43563 1072 43564 1112
rect 43604 1072 43605 1112
rect 43563 1063 43605 1072
rect 43755 1112 43797 1121
rect 43755 1072 43756 1112
rect 43796 1072 43797 1112
rect 43755 1063 43797 1072
rect 43564 978 43604 1063
rect 43756 978 43796 1063
rect 43660 944 43700 953
rect 43660 533 43700 904
rect 43659 524 43701 533
rect 43659 484 43660 524
rect 43700 484 43701 524
rect 43659 475 43701 484
rect 43659 356 43701 365
rect 43659 316 43660 356
rect 43700 316 43701 356
rect 43659 307 43701 316
rect 43660 80 43700 307
rect 43852 80 43892 1660
rect 44140 1280 44180 2500
rect 44236 2465 44276 2584
rect 44235 2456 44277 2465
rect 44235 2416 44236 2456
rect 44276 2416 44277 2456
rect 44235 2407 44277 2416
rect 44332 1457 44372 3928
rect 44620 3809 44660 4012
rect 45003 4003 45045 4012
rect 44812 3968 44852 3977
rect 44716 3928 44812 3968
rect 44619 3800 44661 3809
rect 44619 3760 44620 3800
rect 44660 3760 44661 3800
rect 44619 3751 44661 3760
rect 44619 3632 44661 3641
rect 44619 3592 44620 3632
rect 44660 3592 44661 3632
rect 44619 3583 44661 3592
rect 44427 3548 44469 3557
rect 44427 3508 44428 3548
rect 44468 3508 44469 3548
rect 44427 3499 44469 3508
rect 44428 3464 44468 3499
rect 44428 3413 44468 3424
rect 44620 3464 44660 3583
rect 44524 3212 44564 3221
rect 44524 2540 44564 3172
rect 44620 3137 44660 3424
rect 44619 3128 44661 3137
rect 44619 3088 44620 3128
rect 44660 3088 44661 3128
rect 44619 3079 44661 3088
rect 44524 2500 44660 2540
rect 44331 1448 44373 1457
rect 44331 1408 44332 1448
rect 44372 1408 44373 1448
rect 44331 1399 44373 1408
rect 44140 1240 44276 1280
rect 43948 1112 43988 1121
rect 43948 617 43988 1072
rect 44139 1112 44181 1121
rect 44139 1072 44140 1112
rect 44180 1072 44181 1112
rect 44139 1063 44181 1072
rect 44140 978 44180 1063
rect 44044 944 44084 953
rect 44044 692 44084 904
rect 44139 692 44181 701
rect 44044 652 44140 692
rect 44180 652 44181 692
rect 44139 643 44181 652
rect 43947 608 43989 617
rect 43947 568 43948 608
rect 43988 568 43989 608
rect 43947 559 43989 568
rect 44043 524 44085 533
rect 44043 484 44044 524
rect 44084 484 44085 524
rect 44043 475 44085 484
rect 44044 80 44084 475
rect 44236 80 44276 1240
rect 44343 1205 44383 1220
rect 44342 1196 44384 1205
rect 44342 1156 44343 1196
rect 44383 1156 44384 1196
rect 44342 1147 44384 1156
rect 44343 1125 44383 1147
rect 44343 1076 44383 1085
rect 44427 1113 44469 1121
rect 44524 1113 44564 1121
rect 44427 1112 44564 1113
rect 44427 1072 44428 1112
rect 44468 1073 44524 1112
rect 44468 1072 44469 1073
rect 44427 1063 44469 1072
rect 44524 1063 44564 1072
rect 44428 944 44468 953
rect 44468 904 44564 944
rect 44428 895 44468 904
rect 44331 776 44373 785
rect 44331 736 44332 776
rect 44372 736 44373 776
rect 44331 727 44373 736
rect 44332 449 44372 727
rect 44427 692 44469 701
rect 44427 652 44428 692
rect 44468 652 44469 692
rect 44427 643 44469 652
rect 44331 440 44373 449
rect 44331 400 44332 440
rect 44372 400 44373 440
rect 44331 391 44373 400
rect 44428 80 44468 643
rect 44524 281 44564 904
rect 44523 272 44565 281
rect 44523 232 44524 272
rect 44564 232 44565 272
rect 44523 223 44565 232
rect 44620 80 44660 2500
rect 44716 1112 44756 3928
rect 44812 3919 44852 3928
rect 44811 3548 44853 3557
rect 44811 3508 44812 3548
rect 44852 3508 44853 3548
rect 44811 3499 44853 3508
rect 45195 3548 45237 3557
rect 45195 3508 45196 3548
rect 45236 3508 45237 3548
rect 45195 3499 45237 3508
rect 45579 3548 45621 3557
rect 45579 3508 45580 3548
rect 45620 3508 45621 3548
rect 45579 3499 45621 3508
rect 44812 2624 44852 3499
rect 45196 3464 45236 3499
rect 45196 3413 45236 3424
rect 45387 3464 45429 3473
rect 45580 3464 45620 3499
rect 45387 3424 45388 3464
rect 45428 3424 45524 3464
rect 45387 3415 45429 3424
rect 45388 3330 45428 3415
rect 45292 3212 45332 3221
rect 45003 2876 45045 2885
rect 45003 2836 45004 2876
rect 45044 2836 45045 2876
rect 45003 2827 45045 2836
rect 44812 2575 44852 2584
rect 45004 2624 45044 2827
rect 45004 2575 45044 2584
rect 44908 2540 44948 2549
rect 44908 1280 44948 2500
rect 45292 1280 45332 3172
rect 45484 2213 45524 3424
rect 45580 3413 45620 3424
rect 45772 3464 45812 3473
rect 45676 3212 45716 3221
rect 45483 2204 45525 2213
rect 45483 2164 45484 2204
rect 45524 2164 45525 2204
rect 45483 2155 45525 2164
rect 45676 1616 45716 3172
rect 45772 3053 45812 3424
rect 45771 3044 45813 3053
rect 45771 3004 45772 3044
rect 45812 3004 45813 3044
rect 45771 2995 45813 3004
rect 45772 2129 45812 2995
rect 45868 2540 45908 4348
rect 46060 4145 46100 4230
rect 46059 4136 46101 4145
rect 46059 4096 46060 4136
rect 46100 4096 46101 4136
rect 46059 4087 46101 4096
rect 46060 3968 46100 3977
rect 46060 3809 46100 3928
rect 46059 3800 46101 3809
rect 46059 3760 46060 3800
rect 46100 3760 46101 3800
rect 46059 3751 46101 3760
rect 46156 3632 46196 4684
rect 46252 4229 46292 4843
rect 46348 4724 46388 4733
rect 46388 4684 46484 4724
rect 46348 4675 46388 4684
rect 46251 4220 46293 4229
rect 46251 4180 46252 4220
rect 46292 4180 46293 4220
rect 46251 4171 46293 4180
rect 46252 4136 46292 4171
rect 46252 4086 46292 4096
rect 46347 4136 46389 4145
rect 46347 4096 46348 4136
rect 46388 4096 46389 4136
rect 46347 4087 46389 4096
rect 46348 4002 46388 4087
rect 46156 3592 46292 3632
rect 45963 3548 46005 3557
rect 45963 3508 45964 3548
rect 46004 3508 46005 3548
rect 45963 3499 46005 3508
rect 45964 3464 46004 3499
rect 45964 3413 46004 3424
rect 46156 3464 46196 3473
rect 46060 3212 46100 3221
rect 46060 2540 46100 3172
rect 46156 3053 46196 3424
rect 46155 3044 46197 3053
rect 46155 3004 46156 3044
rect 46196 3004 46197 3044
rect 46155 2995 46197 3004
rect 45868 2500 46004 2540
rect 46060 2500 46196 2540
rect 45771 2120 45813 2129
rect 45771 2080 45772 2120
rect 45812 2080 45813 2120
rect 45771 2071 45813 2080
rect 45676 1576 45812 1616
rect 44908 1240 45044 1280
rect 45292 1240 45428 1280
rect 44716 533 44756 1072
rect 44907 1112 44949 1121
rect 44907 1072 44908 1112
rect 44948 1072 44949 1112
rect 44907 1063 44949 1072
rect 44908 978 44948 1063
rect 44812 944 44852 953
rect 44812 701 44852 904
rect 44811 692 44853 701
rect 44811 652 44812 692
rect 44852 652 44853 692
rect 44811 643 44853 652
rect 44715 524 44757 533
rect 44715 484 44716 524
rect 44756 484 44757 524
rect 44715 475 44757 484
rect 44811 272 44853 281
rect 44811 232 44812 272
rect 44852 232 44853 272
rect 44811 223 44853 232
rect 44812 80 44852 223
rect 45004 80 45044 1240
rect 45100 1205 45140 1236
rect 45099 1196 45141 1205
rect 45099 1156 45100 1196
rect 45140 1156 45141 1196
rect 45099 1147 45141 1156
rect 45100 1112 45140 1147
rect 45100 785 45140 1072
rect 45291 1112 45333 1121
rect 45291 1072 45292 1112
rect 45332 1072 45333 1112
rect 45291 1063 45333 1072
rect 45292 978 45332 1063
rect 45196 944 45236 953
rect 45196 860 45236 904
rect 45196 820 45332 860
rect 45099 776 45141 785
rect 45099 736 45100 776
rect 45140 736 45141 776
rect 45099 727 45141 736
rect 45195 692 45237 701
rect 45195 652 45196 692
rect 45236 652 45237 692
rect 45195 643 45237 652
rect 45196 80 45236 643
rect 45292 617 45332 820
rect 45291 608 45333 617
rect 45291 568 45292 608
rect 45332 568 45333 608
rect 45291 559 45333 568
rect 45388 80 45428 1240
rect 45676 1121 45716 1206
rect 45484 1112 45524 1121
rect 45484 953 45524 1072
rect 45675 1112 45717 1121
rect 45675 1072 45676 1112
rect 45716 1072 45717 1112
rect 45675 1063 45717 1072
rect 45483 944 45525 953
rect 45483 904 45484 944
rect 45524 904 45525 944
rect 45483 895 45525 904
rect 45580 944 45620 953
rect 45580 701 45620 904
rect 45579 692 45621 701
rect 45579 652 45580 692
rect 45620 652 45621 692
rect 45579 643 45621 652
rect 45483 608 45525 617
rect 45483 568 45484 608
rect 45524 568 45525 608
rect 45483 559 45525 568
rect 45484 440 45524 559
rect 45484 400 45620 440
rect 45580 80 45620 400
rect 45772 80 45812 1576
rect 45867 1364 45909 1373
rect 45867 1324 45868 1364
rect 45908 1324 45909 1364
rect 45867 1315 45909 1324
rect 45868 1112 45908 1315
rect 45964 1205 46004 2500
rect 45963 1196 46005 1205
rect 45963 1156 45964 1196
rect 46004 1156 46005 1196
rect 45963 1147 46005 1156
rect 45868 1037 45908 1072
rect 46059 1112 46101 1121
rect 46059 1072 46060 1112
rect 46100 1072 46101 1112
rect 46059 1063 46101 1072
rect 45867 1028 45909 1037
rect 45867 988 45868 1028
rect 45908 988 45909 1028
rect 45867 979 45909 988
rect 45868 948 45908 979
rect 45964 953 46004 1038
rect 46060 978 46100 1063
rect 45963 944 46005 953
rect 45963 904 45964 944
rect 46004 904 46005 944
rect 45963 895 46005 904
rect 45963 692 46005 701
rect 45963 652 45964 692
rect 46004 652 46005 692
rect 45963 643 46005 652
rect 45964 80 46004 643
rect 46156 80 46196 2500
rect 46252 1961 46292 3592
rect 46347 3548 46389 3557
rect 46347 3508 46348 3548
rect 46388 3508 46389 3548
rect 46347 3499 46389 3508
rect 46348 2624 46388 3499
rect 46444 3473 46484 4684
rect 46636 4229 46676 4927
rect 47787 4304 47829 4313
rect 47787 4264 47788 4304
rect 47828 4264 47829 4304
rect 47787 4255 47829 4264
rect 46635 4220 46677 4229
rect 46635 4180 46636 4220
rect 46676 4180 46677 4220
rect 46635 4171 46677 4180
rect 47788 3977 47828 4255
rect 47980 4136 48020 5104
rect 48075 5095 48117 5104
rect 48076 4976 48116 4985
rect 48076 4397 48116 4936
rect 48171 4976 48213 4985
rect 48171 4936 48172 4976
rect 48212 4936 48213 4976
rect 48171 4927 48213 4936
rect 48172 4842 48212 4927
rect 48268 4901 48308 6280
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 48940 5396 48980 6364
rect 49324 5648 49364 6364
rect 49420 6354 49460 6439
rect 56427 6320 56469 6329
rect 56427 6280 56428 6320
rect 56468 6280 56469 6320
rect 56427 6271 56469 6280
rect 53452 5900 53492 5909
rect 53492 5860 53972 5900
rect 53452 5851 53492 5860
rect 51820 5776 52148 5816
rect 49515 5648 49557 5657
rect 49324 5608 49516 5648
rect 49556 5608 49557 5648
rect 49515 5599 49557 5608
rect 50476 5648 50516 5657
rect 48748 5356 48980 5396
rect 48748 4985 48788 5356
rect 48844 5153 48884 5238
rect 48843 5144 48885 5153
rect 48843 5104 48844 5144
rect 48884 5104 48885 5144
rect 48843 5095 48885 5104
rect 49323 5144 49365 5153
rect 49323 5104 49324 5144
rect 49364 5104 49365 5144
rect 49323 5095 49365 5104
rect 48747 4976 48789 4985
rect 48747 4936 48748 4976
rect 48788 4936 48789 4976
rect 48747 4927 48789 4936
rect 48844 4976 48884 4985
rect 48267 4892 48309 4901
rect 48267 4852 48268 4892
rect 48308 4852 48309 4892
rect 48267 4843 48309 4852
rect 48556 4817 48596 4902
rect 48748 4842 48788 4927
rect 48844 4817 48884 4936
rect 49035 4976 49077 4985
rect 49035 4936 49036 4976
rect 49076 4936 49077 4976
rect 49035 4927 49077 4936
rect 49324 4976 49364 5095
rect 48555 4808 48597 4817
rect 48555 4768 48556 4808
rect 48596 4768 48597 4808
rect 48555 4759 48597 4768
rect 48843 4808 48885 4817
rect 48843 4768 48844 4808
rect 48884 4768 48885 4808
rect 48843 4759 48885 4768
rect 48364 4724 48404 4733
rect 48268 4684 48364 4724
rect 48075 4388 48117 4397
rect 48075 4348 48076 4388
rect 48116 4348 48117 4388
rect 48075 4339 48117 4348
rect 48171 4304 48213 4313
rect 48171 4264 48172 4304
rect 48212 4264 48213 4304
rect 48171 4255 48213 4264
rect 48172 4136 48212 4255
rect 47980 4096 48172 4136
rect 48172 4087 48212 4096
rect 47787 3968 47829 3977
rect 47787 3928 47788 3968
rect 47828 3928 47829 3968
rect 47787 3919 47829 3928
rect 48172 3968 48212 3977
rect 47595 3716 47637 3725
rect 47595 3676 47596 3716
rect 47636 3676 47637 3716
rect 47595 3667 47637 3676
rect 47211 3548 47253 3557
rect 47211 3508 47212 3548
rect 47252 3508 47253 3548
rect 47211 3499 47253 3508
rect 46443 3464 46485 3473
rect 46443 3424 46444 3464
rect 46484 3424 46485 3464
rect 46443 3415 46485 3424
rect 46828 3464 46868 3473
rect 46828 3305 46868 3424
rect 47019 3464 47061 3473
rect 47019 3424 47020 3464
rect 47060 3424 47061 3464
rect 47019 3415 47061 3424
rect 47212 3464 47252 3499
rect 47020 3330 47060 3415
rect 46827 3296 46869 3305
rect 46827 3256 46828 3296
rect 46868 3256 46869 3296
rect 46827 3247 46869 3256
rect 46924 3212 46964 3221
rect 46540 2633 46580 2718
rect 46348 2575 46388 2584
rect 46539 2624 46581 2633
rect 46539 2584 46540 2624
rect 46580 2584 46581 2624
rect 46539 2575 46581 2584
rect 46444 2540 46484 2549
rect 46251 1952 46293 1961
rect 46251 1912 46252 1952
rect 46292 1912 46293 1952
rect 46251 1903 46293 1912
rect 46444 1280 46484 2500
rect 46444 1240 46580 1280
rect 46252 1205 46292 1207
rect 46251 1196 46293 1205
rect 46251 1156 46252 1196
rect 46292 1156 46293 1196
rect 46251 1147 46293 1156
rect 46252 1112 46292 1147
rect 46252 1063 46292 1072
rect 46443 1112 46485 1121
rect 46443 1072 46444 1112
rect 46484 1072 46485 1112
rect 46443 1063 46485 1072
rect 46444 978 46484 1063
rect 46251 944 46293 953
rect 46251 904 46252 944
rect 46292 904 46293 944
rect 46251 895 46293 904
rect 46348 944 46388 953
rect 46252 524 46292 895
rect 46348 701 46388 904
rect 46347 692 46389 701
rect 46347 652 46348 692
rect 46388 652 46389 692
rect 46347 643 46389 652
rect 46252 484 46388 524
rect 46348 80 46388 484
rect 46540 80 46580 1240
rect 46636 1205 46676 1236
rect 46635 1196 46677 1205
rect 46635 1156 46636 1196
rect 46676 1156 46677 1196
rect 46635 1147 46677 1156
rect 46636 1112 46676 1147
rect 46636 1037 46676 1072
rect 46827 1112 46869 1121
rect 46827 1072 46828 1112
rect 46868 1072 46869 1112
rect 46827 1063 46869 1072
rect 46635 1028 46677 1037
rect 46635 988 46636 1028
rect 46676 988 46677 1028
rect 46635 979 46677 988
rect 46732 953 46772 1038
rect 46828 978 46868 1063
rect 46731 944 46773 953
rect 46731 904 46732 944
rect 46772 904 46773 944
rect 46731 895 46773 904
rect 46731 692 46773 701
rect 46731 652 46732 692
rect 46772 652 46773 692
rect 46731 643 46773 652
rect 46732 80 46772 643
rect 46924 80 46964 3172
rect 47212 2801 47252 3424
rect 47403 3464 47445 3473
rect 47403 3424 47404 3464
rect 47444 3424 47445 3464
rect 47403 3415 47445 3424
rect 47596 3464 47636 3667
rect 47596 3415 47636 3424
rect 47787 3464 47829 3473
rect 47787 3424 47788 3464
rect 47828 3424 47829 3464
rect 47787 3415 47829 3424
rect 47404 3330 47444 3415
rect 47308 3212 47348 3221
rect 47211 2792 47253 2801
rect 47211 2752 47212 2792
rect 47252 2752 47253 2792
rect 47211 2743 47253 2752
rect 47020 1121 47060 1206
rect 47019 1112 47061 1121
rect 47019 1072 47020 1112
rect 47060 1072 47061 1112
rect 47019 1063 47061 1072
rect 47212 1112 47252 1123
rect 47212 1037 47252 1072
rect 47211 1028 47253 1037
rect 47211 988 47212 1028
rect 47252 988 47253 1028
rect 47211 979 47253 988
rect 47019 944 47061 953
rect 47019 904 47020 944
rect 47060 904 47061 944
rect 47019 895 47061 904
rect 47116 944 47156 953
rect 47020 524 47060 895
rect 47116 701 47156 904
rect 47115 692 47157 701
rect 47115 652 47116 692
rect 47156 652 47157 692
rect 47115 643 47157 652
rect 47020 484 47156 524
rect 47116 80 47156 484
rect 47308 80 47348 3172
rect 47692 3212 47732 3221
rect 47404 1112 47444 1121
rect 47404 869 47444 1072
rect 47596 1112 47636 1123
rect 47500 953 47540 1038
rect 47596 1037 47636 1072
rect 47595 1028 47637 1037
rect 47595 988 47596 1028
rect 47636 988 47637 1028
rect 47595 979 47637 988
rect 47499 944 47541 953
rect 47499 904 47500 944
rect 47540 904 47541 944
rect 47499 895 47541 904
rect 47403 860 47445 869
rect 47403 820 47404 860
rect 47444 820 47445 860
rect 47403 811 47445 820
rect 47499 692 47541 701
rect 47499 652 47500 692
rect 47540 652 47541 692
rect 47499 643 47541 652
rect 47500 80 47540 643
rect 47692 80 47732 3172
rect 47788 2801 47828 3415
rect 48075 3380 48117 3389
rect 48075 3340 48076 3380
rect 48116 3340 48117 3380
rect 48075 3331 48117 3340
rect 48076 2885 48116 3331
rect 48075 2876 48117 2885
rect 48075 2836 48076 2876
rect 48116 2836 48117 2876
rect 48075 2827 48117 2836
rect 47787 2792 47829 2801
rect 47787 2752 47788 2792
rect 47828 2752 47829 2792
rect 47787 2743 47829 2752
rect 47788 2624 47828 2743
rect 48075 2708 48117 2717
rect 48075 2668 48076 2708
rect 48116 2668 48117 2708
rect 48075 2659 48117 2668
rect 47884 2624 47924 2633
rect 47788 2584 47884 2624
rect 47884 2575 47924 2584
rect 48076 2624 48116 2659
rect 48076 2573 48116 2584
rect 47980 2540 48020 2549
rect 47980 1280 48020 2500
rect 48172 1532 48212 3928
rect 48268 3557 48308 4684
rect 48364 4675 48404 4684
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 49036 4313 49076 4927
rect 49324 4817 49364 4936
rect 49516 4976 49556 5599
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 49612 5069 49652 5100
rect 49611 5060 49653 5069
rect 49611 5020 49612 5060
rect 49652 5020 49653 5060
rect 49611 5011 49653 5020
rect 49516 4927 49556 4936
rect 49612 4976 49652 5011
rect 50380 4985 50420 5070
rect 49323 4808 49365 4817
rect 49323 4768 49324 4808
rect 49364 4768 49365 4808
rect 49323 4759 49365 4768
rect 49516 4724 49556 4733
rect 48651 4304 48693 4313
rect 48651 4264 48652 4304
rect 48692 4264 48693 4304
rect 48651 4255 48693 4264
rect 49035 4304 49077 4313
rect 49035 4264 49036 4304
rect 49076 4264 49077 4304
rect 49035 4255 49077 4264
rect 48364 4145 48404 4230
rect 48363 4136 48405 4145
rect 48363 4096 48364 4136
rect 48404 4096 48405 4136
rect 48363 4087 48405 4096
rect 48460 4136 48500 4145
rect 48555 4136 48597 4145
rect 48500 4096 48556 4136
rect 48596 4096 48597 4136
rect 48460 4087 48500 4096
rect 48555 4087 48597 4096
rect 48652 4136 48692 4255
rect 48843 4220 48885 4229
rect 48843 4180 48844 4220
rect 48884 4180 48885 4220
rect 48843 4171 48885 4180
rect 48652 4087 48692 4096
rect 48844 4136 48884 4171
rect 48844 4085 48884 4096
rect 48939 4136 48981 4145
rect 49036 4136 49076 4255
rect 48939 4096 48940 4136
rect 48980 4096 49076 4136
rect 48939 4087 48981 4096
rect 48747 4052 48789 4061
rect 48747 4012 48748 4052
rect 48788 4012 48789 4052
rect 48747 4003 48789 4012
rect 48652 3968 48692 3977
rect 48364 3928 48652 3968
rect 48267 3548 48309 3557
rect 48267 3508 48268 3548
rect 48308 3508 48309 3548
rect 48267 3499 48309 3508
rect 48267 2792 48309 2801
rect 48267 2752 48268 2792
rect 48308 2752 48309 2792
rect 48267 2743 48309 2752
rect 48268 2624 48308 2743
rect 48364 2717 48404 3928
rect 48652 3919 48692 3928
rect 48748 3557 48788 4003
rect 48940 4002 48980 4087
rect 49131 3632 49173 3641
rect 49131 3592 49132 3632
rect 49172 3592 49173 3632
rect 49131 3583 49173 3592
rect 48747 3548 48789 3557
rect 48747 3508 48748 3548
rect 48788 3508 48789 3548
rect 48747 3499 48789 3508
rect 48940 3464 48980 3473
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 48843 2876 48885 2885
rect 48843 2836 48844 2876
rect 48884 2836 48885 2876
rect 48843 2827 48885 2836
rect 48651 2792 48693 2801
rect 48651 2752 48652 2792
rect 48692 2752 48693 2792
rect 48651 2743 48693 2752
rect 48363 2708 48405 2717
rect 48363 2668 48364 2708
rect 48404 2668 48405 2708
rect 48363 2659 48405 2668
rect 48460 2633 48500 2718
rect 48268 2575 48308 2584
rect 48459 2624 48501 2633
rect 48459 2584 48460 2624
rect 48500 2584 48501 2624
rect 48459 2575 48501 2584
rect 48652 2624 48692 2743
rect 48652 2575 48692 2584
rect 48844 2624 48884 2827
rect 48940 2801 48980 3424
rect 49132 3464 49172 3583
rect 49132 3221 49172 3424
rect 49036 3212 49076 3221
rect 48939 2792 48981 2801
rect 48939 2752 48940 2792
rect 48980 2752 48981 2792
rect 48939 2743 48981 2752
rect 48844 2575 48884 2584
rect 48364 2540 48404 2549
rect 48172 1492 48308 1532
rect 47980 1240 48116 1280
rect 47788 1121 47828 1206
rect 47787 1112 47829 1121
rect 47787 1072 47788 1112
rect 47828 1072 47829 1112
rect 47787 1063 47829 1072
rect 47980 1112 48020 1123
rect 47980 1037 48020 1072
rect 47979 1028 48021 1037
rect 47979 988 47980 1028
rect 48020 988 48021 1028
rect 47979 979 48021 988
rect 47787 944 47829 953
rect 47787 904 47788 944
rect 47828 904 47829 944
rect 47787 895 47829 904
rect 47884 944 47924 953
rect 47788 524 47828 895
rect 47884 701 47924 904
rect 47883 692 47925 701
rect 47883 652 47884 692
rect 47924 652 47925 692
rect 47883 643 47925 652
rect 47788 484 47924 524
rect 47884 80 47924 484
rect 48076 80 48116 1240
rect 48268 1205 48308 1492
rect 48364 1280 48404 2500
rect 48748 2540 48788 2549
rect 48748 1700 48788 2500
rect 49036 1700 49076 3172
rect 49131 3212 49173 3221
rect 49131 3172 49132 3212
rect 49172 3172 49173 3212
rect 49131 3163 49173 3172
rect 49131 2792 49173 2801
rect 49131 2752 49132 2792
rect 49172 2752 49173 2792
rect 49131 2743 49173 2752
rect 49132 2624 49172 2743
rect 49324 2633 49364 2718
rect 49132 2575 49172 2584
rect 49323 2624 49365 2633
rect 49323 2584 49324 2624
rect 49364 2584 49365 2624
rect 49323 2575 49365 2584
rect 49228 2540 49268 2549
rect 49228 1784 49268 2500
rect 49516 1868 49556 4684
rect 49612 4229 49652 4936
rect 50379 4976 50421 4985
rect 50379 4936 50380 4976
rect 50420 4936 50421 4976
rect 50379 4927 50421 4936
rect 50476 4901 50516 5608
rect 50668 5648 50708 5657
rect 50572 5564 50612 5573
rect 50572 4976 50612 5524
rect 50668 5153 50708 5608
rect 51243 5312 51285 5321
rect 51243 5272 51244 5312
rect 51284 5272 51285 5312
rect 51243 5263 51285 5272
rect 50667 5144 50709 5153
rect 50667 5104 50668 5144
rect 50708 5104 50709 5144
rect 50667 5095 50709 5104
rect 50860 5069 50900 5082
rect 50859 5060 50901 5069
rect 50859 5020 50860 5060
rect 50900 5020 50901 5060
rect 50859 5011 50901 5020
rect 50860 4987 50900 5011
rect 50668 4976 50708 4985
rect 50572 4936 50668 4976
rect 50860 4938 50900 4947
rect 50475 4892 50517 4901
rect 50475 4852 50476 4892
rect 50516 4852 50517 4892
rect 50475 4843 50517 4852
rect 50380 4808 50420 4819
rect 50380 4733 50420 4768
rect 50188 4724 50228 4733
rect 50092 4684 50188 4724
rect 49611 4220 49653 4229
rect 49611 4180 49612 4220
rect 49652 4180 49653 4220
rect 49611 4171 49653 4180
rect 50092 3968 50132 4684
rect 50188 4675 50228 4684
rect 50379 4724 50421 4733
rect 50379 4684 50380 4724
rect 50420 4684 50421 4724
rect 50379 4675 50421 4684
rect 50187 4556 50229 4565
rect 50187 4516 50188 4556
rect 50228 4516 50229 4556
rect 50187 4507 50229 4516
rect 50188 4145 50228 4507
rect 50187 4136 50229 4145
rect 50187 4096 50188 4136
rect 50228 4096 50229 4136
rect 50187 4087 50229 4096
rect 50380 4136 50420 4145
rect 50476 4136 50516 4843
rect 50668 4733 50708 4936
rect 50764 4892 50804 4901
rect 50667 4724 50709 4733
rect 50667 4684 50668 4724
rect 50708 4684 50709 4724
rect 50667 4675 50709 4684
rect 50667 4388 50709 4397
rect 50667 4348 50668 4388
rect 50708 4348 50709 4388
rect 50667 4339 50709 4348
rect 50668 4220 50708 4339
rect 50764 4304 50804 4852
rect 51244 4817 51284 5263
rect 51531 4976 51573 4985
rect 51531 4936 51532 4976
rect 51572 4936 51573 4976
rect 51531 4927 51573 4936
rect 51532 4817 51572 4927
rect 51243 4808 51285 4817
rect 51243 4768 51244 4808
rect 51284 4768 51285 4808
rect 51243 4759 51285 4768
rect 51531 4808 51573 4817
rect 51531 4768 51532 4808
rect 51572 4768 51573 4808
rect 51531 4759 51573 4768
rect 50764 4264 50900 4304
rect 50668 4180 50804 4220
rect 50572 4145 50612 4164
rect 50571 4136 50613 4145
rect 50420 4096 50572 4136
rect 50612 4096 50613 4136
rect 50380 4087 50420 4096
rect 50571 4087 50613 4096
rect 50764 4136 50804 4180
rect 50764 4087 50804 4096
rect 50284 4052 50324 4061
rect 50092 3928 50228 3968
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 50091 3464 50133 3473
rect 50091 3424 50092 3464
rect 50132 3424 50133 3464
rect 50091 3415 50133 3424
rect 50092 3330 50132 3415
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 49516 1828 49748 1868
rect 49228 1744 49652 1784
rect 48748 1660 48980 1700
rect 49036 1660 49268 1700
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 48555 1280 48597 1289
rect 48940 1280 48980 1660
rect 48364 1240 48500 1280
rect 48166 1196 48208 1205
rect 48267 1196 48309 1205
rect 48166 1156 48167 1196
rect 48207 1156 48212 1196
rect 48166 1147 48212 1156
rect 48267 1156 48268 1196
rect 48308 1156 48309 1196
rect 48267 1147 48309 1156
rect 48172 1112 48212 1147
rect 48172 1063 48212 1072
rect 48364 1112 48404 1123
rect 48268 953 48308 1038
rect 48364 1037 48404 1072
rect 48363 1028 48405 1037
rect 48363 988 48364 1028
rect 48404 988 48405 1028
rect 48363 979 48405 988
rect 48267 944 48309 953
rect 48267 904 48268 944
rect 48308 904 48309 944
rect 48267 895 48309 904
rect 48267 692 48309 701
rect 48267 652 48268 692
rect 48308 652 48309 692
rect 48267 643 48309 652
rect 48268 80 48308 643
rect 48460 80 48500 1240
rect 48555 1240 48556 1280
rect 48596 1240 48597 1280
rect 48555 1231 48597 1240
rect 48844 1240 48980 1280
rect 48556 1112 48596 1231
rect 48748 1205 48788 1236
rect 48747 1196 48789 1205
rect 48747 1156 48748 1196
rect 48788 1156 48789 1196
rect 48747 1147 48789 1156
rect 48556 1063 48596 1072
rect 48748 1112 48788 1147
rect 48748 1037 48788 1072
rect 48747 1028 48789 1037
rect 48747 988 48748 1028
rect 48788 988 48789 1028
rect 48747 979 48789 988
rect 48555 944 48597 953
rect 48555 904 48556 944
rect 48596 904 48597 944
rect 48555 895 48597 904
rect 48652 944 48692 953
rect 48556 524 48596 895
rect 48652 701 48692 904
rect 48651 692 48693 701
rect 48651 652 48652 692
rect 48692 652 48693 692
rect 48651 643 48693 652
rect 48556 484 48692 524
rect 48652 80 48692 484
rect 48844 80 48884 1240
rect 49131 1196 49173 1205
rect 49131 1156 49132 1196
rect 49172 1156 49173 1196
rect 49131 1147 49173 1156
rect 48939 1112 48981 1121
rect 48939 1072 48940 1112
rect 48980 1072 48981 1112
rect 48939 1063 48981 1072
rect 49132 1112 49172 1147
rect 48940 978 48980 1063
rect 49132 1061 49172 1072
rect 49036 944 49076 953
rect 49076 904 49172 944
rect 49036 895 49076 904
rect 49035 692 49077 701
rect 49035 652 49036 692
rect 49076 652 49077 692
rect 49035 643 49077 652
rect 49036 80 49076 643
rect 49132 197 49172 904
rect 49131 188 49173 197
rect 49131 148 49132 188
rect 49172 148 49173 188
rect 49131 139 49173 148
rect 49228 80 49268 1660
rect 49515 1280 49557 1289
rect 49515 1240 49516 1280
rect 49556 1240 49557 1280
rect 49515 1231 49557 1240
rect 49323 1196 49365 1205
rect 49323 1156 49324 1196
rect 49364 1156 49365 1196
rect 49323 1147 49365 1156
rect 49324 1112 49364 1147
rect 49324 1061 49364 1072
rect 49516 1112 49556 1231
rect 49516 1063 49556 1072
rect 49420 944 49460 953
rect 49420 533 49460 904
rect 49419 524 49461 533
rect 49419 484 49420 524
rect 49460 484 49461 524
rect 49419 475 49461 484
rect 49419 188 49461 197
rect 49419 148 49420 188
rect 49460 148 49461 188
rect 49419 139 49461 148
rect 49420 80 49460 139
rect 49612 80 49652 1744
rect 49708 1205 49748 1828
rect 49803 1364 49845 1373
rect 49803 1324 49804 1364
rect 49844 1324 49845 1364
rect 49803 1315 49845 1324
rect 49707 1196 49749 1205
rect 49707 1156 49708 1196
rect 49748 1156 49749 1196
rect 49707 1147 49749 1156
rect 49804 1037 49844 1315
rect 49803 1028 49845 1037
rect 49803 988 49804 1028
rect 49844 988 49845 1028
rect 49803 979 49845 988
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 50188 608 50228 3928
rect 50284 3632 50324 4012
rect 50572 4002 50612 4087
rect 50668 4052 50708 4061
rect 50668 3968 50708 4012
rect 50668 3928 50804 3968
rect 50284 3592 50420 3632
rect 50284 3464 50324 3475
rect 50284 3389 50324 3424
rect 50283 3380 50325 3389
rect 50283 3340 50284 3380
rect 50324 3340 50325 3380
rect 50283 3331 50325 3340
rect 50284 3212 50324 3221
rect 50284 1625 50324 3172
rect 50380 3053 50420 3592
rect 50668 3473 50708 3558
rect 50667 3464 50709 3473
rect 50667 3424 50668 3464
rect 50708 3424 50709 3464
rect 50667 3415 50709 3424
rect 50764 3305 50804 3928
rect 50668 3296 50708 3305
rect 50763 3296 50805 3305
rect 50708 3256 50764 3296
rect 50804 3256 50805 3296
rect 50668 3247 50708 3256
rect 50763 3247 50805 3256
rect 50764 3228 50804 3247
rect 50476 3212 50516 3221
rect 50379 3044 50421 3053
rect 50379 3004 50380 3044
rect 50420 3004 50421 3044
rect 50379 2995 50421 3004
rect 50283 1616 50325 1625
rect 50283 1576 50284 1616
rect 50324 1576 50325 1616
rect 50283 1567 50325 1576
rect 50476 1364 50516 3172
rect 50571 3044 50613 3053
rect 50571 3004 50572 3044
rect 50612 3004 50613 3044
rect 50571 2995 50613 3004
rect 50284 1324 50516 1364
rect 50284 944 50324 1324
rect 50572 1289 50612 2995
rect 50667 1616 50709 1625
rect 50667 1576 50668 1616
rect 50708 1576 50709 1616
rect 50667 1567 50709 1576
rect 50571 1280 50613 1289
rect 50571 1240 50572 1280
rect 50612 1240 50613 1280
rect 50571 1231 50613 1240
rect 50379 1196 50421 1205
rect 50379 1156 50380 1196
rect 50420 1156 50421 1196
rect 50379 1147 50421 1156
rect 50380 1112 50420 1147
rect 50380 1061 50420 1072
rect 50572 1112 50612 1231
rect 50572 1063 50612 1072
rect 50475 944 50517 953
rect 50284 904 50420 944
rect 50283 776 50325 785
rect 50283 736 50284 776
rect 50324 736 50325 776
rect 50283 727 50325 736
rect 49996 568 50228 608
rect 49803 524 49845 533
rect 49803 484 49804 524
rect 49844 484 49845 524
rect 49803 475 49845 484
rect 49804 80 49844 475
rect 49996 80 50036 568
rect 50284 440 50324 727
rect 50188 400 50324 440
rect 50188 80 50228 400
rect 50380 80 50420 904
rect 50475 904 50476 944
rect 50516 904 50517 944
rect 50475 895 50517 904
rect 50476 810 50516 895
rect 50668 860 50708 1567
rect 50572 820 50708 860
rect 50764 944 50804 953
rect 50572 80 50612 820
rect 50764 80 50804 904
rect 50860 785 50900 4264
rect 50955 4136 50997 4145
rect 50955 4096 50956 4136
rect 50996 4096 50997 4136
rect 50955 4087 50997 4096
rect 51244 4136 51284 4759
rect 51435 4388 51477 4397
rect 51435 4348 51436 4388
rect 51476 4348 51477 4388
rect 51435 4339 51477 4348
rect 51436 4145 51476 4339
rect 51532 4313 51572 4759
rect 51820 4565 51860 5776
rect 51916 5648 51956 5659
rect 51916 5573 51956 5608
rect 52108 5648 52148 5776
rect 52588 5692 53012 5732
rect 52108 5599 52148 5608
rect 52492 5648 52532 5657
rect 51915 5564 51957 5573
rect 51915 5524 51916 5564
rect 51956 5524 51957 5564
rect 51915 5515 51957 5524
rect 52012 5564 52052 5573
rect 52012 5069 52052 5524
rect 52300 5564 52340 5573
rect 52300 5480 52340 5524
rect 52108 5440 52340 5480
rect 52011 5060 52053 5069
rect 52011 5020 52012 5060
rect 52052 5020 52053 5060
rect 52011 5011 52053 5020
rect 52108 4892 52148 5440
rect 52492 5228 52532 5608
rect 52588 5648 52628 5692
rect 52588 5599 52628 5608
rect 52779 5564 52821 5573
rect 52779 5524 52780 5564
rect 52820 5524 52821 5564
rect 52779 5515 52821 5524
rect 52588 5480 52628 5489
rect 52588 5321 52628 5440
rect 52587 5312 52629 5321
rect 52587 5272 52588 5312
rect 52628 5272 52629 5312
rect 52587 5263 52629 5272
rect 52204 5188 52532 5228
rect 52204 4985 52244 5188
rect 52299 5060 52341 5069
rect 52299 5020 52300 5060
rect 52340 5020 52341 5060
rect 52299 5011 52341 5020
rect 52203 4976 52245 4985
rect 52203 4936 52204 4976
rect 52244 4936 52245 4976
rect 52203 4927 52245 4936
rect 52012 4852 52148 4892
rect 51819 4556 51861 4565
rect 51819 4516 51820 4556
rect 51860 4516 51861 4556
rect 51819 4507 51861 4516
rect 51531 4304 51573 4313
rect 51531 4264 51532 4304
rect 51572 4264 51573 4304
rect 51531 4255 51573 4264
rect 51244 4087 51284 4096
rect 51435 4136 51477 4145
rect 51435 4096 51436 4136
rect 51476 4096 51477 4136
rect 51435 4087 51477 4096
rect 51532 4136 51572 4255
rect 51532 4087 51572 4096
rect 50956 3464 50996 4087
rect 51436 4002 51476 4087
rect 51243 3968 51285 3977
rect 51243 3928 51244 3968
rect 51284 3928 51285 3968
rect 51243 3919 51285 3928
rect 51147 3548 51189 3557
rect 51147 3508 51148 3548
rect 51188 3508 51189 3548
rect 51147 3499 51189 3508
rect 50956 3415 50996 3424
rect 51148 3464 51188 3499
rect 51148 3413 51188 3424
rect 51052 3212 51092 3221
rect 51052 2045 51092 3172
rect 51244 2120 51284 3919
rect 52012 3473 52052 4852
rect 52300 4808 52340 5011
rect 52396 4985 52436 5070
rect 52683 5060 52725 5069
rect 52683 5020 52684 5060
rect 52724 5020 52725 5060
rect 52683 5011 52725 5020
rect 52685 4987 52725 5011
rect 52395 4976 52437 4985
rect 52395 4936 52396 4976
rect 52436 4936 52437 4976
rect 52395 4927 52437 4936
rect 52685 4926 52725 4947
rect 52396 4808 52436 4817
rect 52300 4768 52396 4808
rect 52396 4759 52436 4768
rect 52204 4724 52244 4733
rect 52684 4724 52724 4733
rect 52108 4684 52204 4724
rect 52011 3464 52053 3473
rect 52011 3424 52012 3464
rect 52052 3424 52053 3464
rect 52011 3415 52053 3424
rect 52012 3221 52052 3415
rect 52011 3212 52053 3221
rect 52011 3172 52012 3212
rect 52052 3172 52053 3212
rect 52011 3163 52053 3172
rect 51819 2288 51861 2297
rect 51819 2248 51820 2288
rect 51860 2248 51861 2288
rect 51819 2239 51861 2248
rect 51148 2080 51284 2120
rect 51051 2036 51093 2045
rect 51051 1996 51052 2036
rect 51092 1996 51093 2036
rect 51051 1987 51093 1996
rect 50956 1289 50996 1374
rect 51051 1364 51093 1373
rect 51051 1324 51052 1364
rect 51092 1324 51093 1364
rect 51051 1315 51093 1324
rect 50955 1280 50997 1289
rect 50955 1240 50956 1280
rect 50996 1240 50997 1280
rect 50955 1231 50997 1240
rect 50956 1112 50996 1121
rect 51052 1112 51092 1315
rect 51148 1121 51188 2080
rect 51435 2036 51477 2045
rect 51435 1996 51436 2036
rect 51476 1996 51477 2036
rect 51435 1987 51477 1996
rect 51243 1952 51285 1961
rect 51243 1912 51244 1952
rect 51284 1912 51285 1952
rect 51243 1903 51285 1912
rect 51436 1952 51476 1987
rect 51724 1961 51764 1980
rect 51244 1818 51284 1903
rect 51436 1877 51476 1912
rect 51723 1952 51765 1961
rect 51820 1952 51860 2239
rect 52108 2120 52148 4684
rect 52204 4675 52244 4684
rect 52588 4684 52684 4724
rect 52588 4397 52628 4684
rect 52684 4675 52724 4684
rect 52203 4388 52245 4397
rect 52300 4388 52340 4397
rect 52203 4348 52204 4388
rect 52244 4348 52300 4388
rect 52203 4339 52245 4348
rect 52300 4339 52340 4348
rect 52587 4388 52629 4397
rect 52587 4348 52588 4388
rect 52628 4348 52629 4388
rect 52587 4339 52629 4348
rect 52780 4304 52820 5515
rect 52876 4976 52916 4987
rect 52972 4985 53012 5692
rect 53740 5657 53780 5742
rect 53644 5648 53684 5657
rect 53548 5608 53644 5648
rect 53548 4985 53588 5608
rect 53644 5599 53684 5608
rect 53739 5648 53781 5657
rect 53739 5608 53740 5648
rect 53780 5608 53781 5648
rect 53739 5599 53781 5608
rect 53740 5480 53780 5489
rect 53740 5321 53780 5440
rect 53739 5312 53781 5321
rect 53739 5272 53740 5312
rect 53780 5272 53781 5312
rect 53739 5263 53781 5272
rect 52876 4901 52916 4936
rect 52971 4976 53013 4985
rect 52971 4936 52972 4976
rect 53012 4936 53013 4976
rect 52971 4927 53013 4936
rect 53547 4976 53589 4985
rect 53547 4936 53548 4976
rect 53588 4936 53589 4976
rect 53547 4927 53589 4936
rect 53740 4976 53780 4985
rect 52875 4892 52917 4901
rect 52875 4852 52876 4892
rect 52916 4852 52917 4892
rect 52875 4843 52917 4852
rect 52972 4313 53012 4927
rect 53548 4842 53588 4927
rect 53740 4817 53780 4936
rect 53835 4892 53877 4901
rect 53835 4852 53836 4892
rect 53876 4852 53877 4892
rect 53835 4843 53877 4852
rect 53451 4808 53493 4817
rect 53451 4768 53452 4808
rect 53492 4768 53493 4808
rect 53451 4759 53493 4768
rect 53739 4808 53781 4817
rect 53739 4768 53740 4808
rect 53780 4768 53781 4808
rect 53739 4759 53781 4768
rect 53356 4313 53396 4398
rect 52971 4304 53013 4313
rect 52684 4264 52916 4304
rect 52203 4220 52245 4229
rect 52684 4220 52724 4264
rect 52203 4180 52204 4220
rect 52244 4180 52245 4220
rect 52203 4171 52245 4180
rect 52588 4180 52724 4220
rect 52204 4136 52244 4171
rect 52396 4151 52436 4160
rect 52588 4151 52628 4180
rect 52436 4111 52588 4136
rect 52396 4096 52628 4111
rect 52779 4136 52821 4145
rect 52779 4096 52780 4136
rect 52820 4096 52821 4136
rect 52204 4085 52244 4096
rect 52779 4087 52821 4096
rect 52684 4052 52724 4061
rect 52492 4012 52684 4052
rect 52492 3296 52532 4012
rect 52684 4003 52724 4012
rect 52780 4002 52820 4087
rect 52876 3884 52916 4264
rect 52971 4264 52972 4304
rect 53012 4264 53013 4304
rect 52971 4255 53013 4264
rect 53355 4304 53397 4313
rect 53355 4264 53356 4304
rect 53396 4264 53397 4304
rect 53355 4255 53397 4264
rect 53355 4136 53397 4145
rect 53355 4096 53356 4136
rect 53396 4096 53397 4136
rect 53355 4087 53397 4096
rect 53356 4002 53396 4087
rect 52588 3844 52916 3884
rect 53164 3968 53204 3977
rect 52588 3464 52628 3844
rect 52779 3548 52821 3557
rect 52779 3508 52780 3548
rect 52820 3508 52821 3548
rect 52779 3499 52821 3508
rect 52588 3415 52628 3424
rect 52780 3464 52820 3499
rect 52780 3413 52820 3424
rect 52684 3296 52724 3305
rect 52492 3256 52628 3296
rect 52299 2288 52341 2297
rect 52299 2248 52300 2288
rect 52340 2248 52341 2288
rect 52299 2239 52341 2248
rect 52108 2080 52244 2120
rect 51723 1912 51724 1952
rect 51764 1912 51820 1952
rect 51723 1903 51765 1912
rect 51820 1903 51860 1912
rect 51915 1952 51957 1961
rect 51915 1912 51916 1952
rect 51956 1912 51957 1952
rect 51915 1903 51957 1912
rect 52107 1952 52149 1961
rect 52107 1912 52108 1952
rect 52148 1912 52149 1952
rect 52107 1903 52149 1912
rect 51340 1868 51380 1877
rect 51340 1280 51380 1828
rect 51435 1868 51477 1877
rect 51435 1828 51436 1868
rect 51476 1828 51477 1868
rect 51435 1819 51477 1828
rect 51244 1240 51380 1280
rect 51436 1254 51476 1819
rect 51820 1784 51860 1793
rect 51916 1784 51956 1903
rect 52108 1818 52148 1903
rect 51860 1744 51956 1784
rect 52204 1784 52244 2080
rect 52300 1952 52340 2239
rect 52300 1903 52340 1912
rect 52204 1744 52340 1784
rect 51820 1735 51860 1744
rect 51628 1700 51668 1709
rect 52108 1700 52148 1709
rect 50996 1072 51092 1112
rect 51147 1112 51189 1121
rect 51147 1072 51148 1112
rect 51188 1072 51189 1112
rect 51244 1112 51284 1240
rect 51436 1205 51476 1214
rect 51532 1660 51628 1700
rect 51435 1112 51477 1121
rect 51244 1072 51380 1112
rect 50956 1063 50996 1072
rect 51147 1063 51189 1072
rect 50955 944 50997 953
rect 51244 944 51284 953
rect 50955 904 50956 944
rect 50996 904 50997 944
rect 50955 895 50997 904
rect 51148 904 51244 944
rect 50859 776 50901 785
rect 50859 736 50860 776
rect 50900 736 50901 776
rect 50859 727 50901 736
rect 50956 80 50996 895
rect 51148 80 51188 904
rect 51244 895 51284 904
rect 51340 80 51380 1072
rect 51435 1072 51436 1112
rect 51476 1072 51477 1112
rect 51435 1063 51477 1072
rect 51436 978 51476 1063
rect 51532 80 51572 1660
rect 51628 1651 51668 1660
rect 51916 1660 52108 1700
rect 51916 1028 51956 1660
rect 52108 1651 52148 1660
rect 52204 1289 52244 1374
rect 52203 1280 52245 1289
rect 52203 1240 52204 1280
rect 52244 1240 52245 1280
rect 52203 1231 52245 1240
rect 52203 1112 52245 1121
rect 52203 1072 52204 1112
rect 52244 1072 52245 1112
rect 52203 1063 52245 1072
rect 51724 988 51956 1028
rect 51724 80 51764 988
rect 52204 978 52244 1063
rect 52012 944 52052 953
rect 51916 904 52012 944
rect 51916 80 51956 904
rect 52012 895 52052 904
rect 52107 944 52149 953
rect 52107 904 52108 944
rect 52148 904 52149 944
rect 52107 895 52149 904
rect 52108 80 52148 895
rect 52300 80 52340 1744
rect 52588 1289 52628 3256
rect 52684 2540 52724 3256
rect 52684 2500 52820 2540
rect 52780 1784 52820 2500
rect 52875 2288 52917 2297
rect 52875 2248 52876 2288
rect 52916 2248 52917 2288
rect 52875 2239 52917 2248
rect 52876 1952 52916 2239
rect 53164 2120 53204 3928
rect 53452 3809 53492 4759
rect 53644 4724 53684 4733
rect 53644 4313 53684 4684
rect 53836 4649 53876 4843
rect 53835 4640 53877 4649
rect 53835 4600 53836 4640
rect 53876 4600 53877 4640
rect 53835 4591 53877 4600
rect 53643 4304 53685 4313
rect 53643 4264 53644 4304
rect 53684 4264 53685 4304
rect 53643 4255 53685 4264
rect 53644 4136 53684 4255
rect 53836 4145 53876 4591
rect 53644 4087 53684 4096
rect 53835 4136 53877 4145
rect 53835 4096 53836 4136
rect 53876 4096 53877 4136
rect 53835 4087 53877 4096
rect 53836 4002 53876 4087
rect 53740 3968 53780 3977
rect 53451 3800 53493 3809
rect 53451 3760 53452 3800
rect 53492 3760 53493 3800
rect 53451 3751 53493 3760
rect 53259 3548 53301 3557
rect 53259 3508 53260 3548
rect 53300 3508 53301 3548
rect 53259 3499 53301 3508
rect 53260 3464 53300 3499
rect 53260 3413 53300 3424
rect 53452 3464 53492 3751
rect 53452 3415 53492 3424
rect 53355 3212 53397 3221
rect 53355 3172 53356 3212
rect 53396 3172 53397 3212
rect 53355 3163 53397 3172
rect 53356 3078 53396 3163
rect 53740 2540 53780 3928
rect 53932 3389 53972 5860
rect 54316 5648 54356 5657
rect 54316 4985 54356 5608
rect 54507 5648 54549 5657
rect 54507 5608 54508 5648
rect 54548 5608 54549 5648
rect 54507 5599 54549 5608
rect 55468 5648 55508 5657
rect 54412 5564 54452 5573
rect 54315 4976 54357 4985
rect 54315 4936 54316 4976
rect 54356 4936 54357 4976
rect 54315 4927 54357 4936
rect 54412 4901 54452 5524
rect 54508 5514 54548 5599
rect 55276 5564 55316 5573
rect 55316 5524 55412 5564
rect 55276 5515 55316 5524
rect 55083 5312 55125 5321
rect 55083 5272 55084 5312
rect 55124 5272 55125 5312
rect 55083 5263 55125 5272
rect 54796 5020 54932 5060
rect 54411 4892 54453 4901
rect 54411 4852 54412 4892
rect 54452 4852 54453 4892
rect 54411 4843 54453 4852
rect 54700 4724 54740 4733
rect 54604 4684 54700 4724
rect 53931 3380 53973 3389
rect 53931 3340 53932 3380
rect 53972 3340 53973 3380
rect 53931 3331 53973 3340
rect 54219 3212 54261 3221
rect 54219 3172 54220 3212
rect 54260 3172 54261 3212
rect 54219 3163 54261 3172
rect 53548 2500 53780 2540
rect 53355 2288 53397 2297
rect 53355 2248 53356 2288
rect 53396 2248 53397 2288
rect 53355 2239 53397 2248
rect 53164 2080 53300 2120
rect 52876 1903 52916 1912
rect 52971 1952 53013 1961
rect 52971 1912 52972 1952
rect 53012 1912 53013 1952
rect 52971 1903 53013 1912
rect 53163 1952 53205 1961
rect 53163 1912 53164 1952
rect 53204 1912 53205 1952
rect 53163 1903 53205 1912
rect 52876 1784 52916 1793
rect 52972 1784 53012 1903
rect 53164 1818 53204 1903
rect 52780 1744 52876 1784
rect 52916 1744 53012 1784
rect 52876 1735 52916 1744
rect 52684 1700 52724 1709
rect 53164 1700 53204 1709
rect 52724 1660 52820 1700
rect 52684 1651 52724 1660
rect 52587 1280 52629 1289
rect 52587 1240 52588 1280
rect 52628 1240 52629 1280
rect 52587 1231 52629 1240
rect 52492 1112 52532 1121
rect 52588 1112 52628 1231
rect 52532 1072 52628 1112
rect 52683 1112 52725 1121
rect 52683 1072 52684 1112
rect 52724 1072 52725 1112
rect 52492 1063 52532 1072
rect 52683 1063 52725 1072
rect 52684 978 52724 1063
rect 52587 944 52629 953
rect 52587 904 52588 944
rect 52628 904 52629 944
rect 52587 895 52629 904
rect 52588 810 52628 895
rect 52780 860 52820 1660
rect 52972 1660 53164 1700
rect 52972 1280 53012 1660
rect 53164 1651 53204 1660
rect 53260 1532 53300 2080
rect 53356 1952 53396 2239
rect 53356 1903 53396 1912
rect 52684 820 52820 860
rect 52876 1240 53012 1280
rect 53068 1492 53300 1532
rect 52491 776 52533 785
rect 52491 736 52492 776
rect 52532 736 52533 776
rect 52491 727 52533 736
rect 52492 80 52532 727
rect 52684 80 52724 820
rect 52876 80 52916 1240
rect 53068 80 53108 1492
rect 53548 1448 53588 2500
rect 54027 1700 54069 1709
rect 54027 1660 54028 1700
rect 54068 1660 54069 1700
rect 54027 1651 54069 1660
rect 53739 1616 53781 1625
rect 53739 1576 53740 1616
rect 53780 1576 53781 1616
rect 53739 1567 53781 1576
rect 53260 1408 53588 1448
rect 53260 80 53300 1408
rect 53547 1112 53589 1121
rect 53547 1072 53548 1112
rect 53588 1072 53589 1112
rect 53547 1063 53589 1072
rect 53740 1112 53780 1567
rect 53740 1063 53780 1072
rect 53548 978 53588 1063
rect 53451 944 53493 953
rect 53451 904 53452 944
rect 53492 904 53493 944
rect 53451 895 53493 904
rect 53644 944 53684 953
rect 53452 80 53492 895
rect 53547 524 53589 533
rect 53547 484 53548 524
rect 53588 484 53589 524
rect 53547 475 53589 484
rect 53548 197 53588 475
rect 53547 188 53589 197
rect 53547 148 53548 188
rect 53588 148 53589 188
rect 53547 139 53589 148
rect 53644 80 53684 904
rect 53931 944 53973 953
rect 53931 904 53932 944
rect 53972 904 53973 944
rect 53931 895 53973 904
rect 53932 810 53972 895
rect 53835 524 53877 533
rect 53835 484 53836 524
rect 53876 484 53877 524
rect 53835 475 53877 484
rect 53836 80 53876 475
rect 54028 80 54068 1651
rect 54123 1616 54165 1625
rect 54123 1576 54124 1616
rect 54164 1576 54165 1616
rect 54123 1567 54165 1576
rect 54124 1280 54164 1567
rect 54220 1373 54260 3163
rect 54507 3044 54549 3053
rect 54507 3004 54508 3044
rect 54548 3004 54549 3044
rect 54507 2995 54549 3004
rect 54315 2288 54357 2297
rect 54315 2248 54316 2288
rect 54356 2248 54357 2288
rect 54315 2239 54357 2248
rect 54316 1952 54356 2239
rect 54316 1903 54356 1912
rect 54508 1952 54548 2995
rect 54508 1868 54548 1912
rect 54412 1828 54548 1868
rect 54412 1457 54452 1828
rect 54507 1700 54549 1709
rect 54507 1660 54508 1700
rect 54548 1660 54549 1700
rect 54507 1651 54549 1660
rect 54508 1566 54548 1651
rect 54411 1448 54453 1457
rect 54411 1408 54412 1448
rect 54452 1408 54453 1448
rect 54604 1448 54644 4684
rect 54700 4675 54740 4684
rect 54796 4649 54836 5020
rect 54892 4976 54932 5020
rect 54892 4927 54932 4936
rect 54891 4808 54933 4817
rect 54891 4768 54892 4808
rect 54932 4768 54933 4808
rect 54891 4759 54933 4768
rect 54892 4674 54932 4759
rect 54795 4640 54837 4649
rect 54795 4600 54796 4640
rect 54836 4600 54837 4640
rect 54795 4591 54837 4600
rect 54796 4304 54836 4591
rect 54700 4264 54836 4304
rect 54700 2624 54740 4264
rect 54891 4220 54933 4229
rect 54891 4180 54892 4220
rect 54932 4180 54933 4220
rect 54891 4171 54933 4180
rect 54795 4136 54837 4145
rect 54795 4096 54796 4136
rect 54836 4096 54837 4136
rect 54795 4087 54837 4096
rect 54700 2297 54740 2584
rect 54699 2288 54741 2297
rect 54699 2248 54700 2288
rect 54740 2248 54741 2288
rect 54699 2239 54741 2248
rect 54604 1408 54740 1448
rect 54411 1399 54453 1408
rect 54219 1364 54261 1373
rect 54219 1324 54220 1364
rect 54260 1324 54261 1364
rect 54219 1315 54261 1324
rect 54124 1231 54164 1240
rect 54220 1254 54260 1315
rect 54604 1280 54644 1289
rect 54220 1240 54604 1254
rect 54220 1214 54644 1240
rect 54604 1124 54644 1133
rect 54123 1112 54165 1121
rect 54123 1072 54124 1112
rect 54164 1072 54165 1112
rect 54123 1063 54165 1072
rect 54507 1112 54549 1121
rect 54507 1072 54508 1112
rect 54548 1084 54604 1112
rect 54548 1072 54644 1084
rect 54507 1063 54549 1072
rect 54124 978 54164 1063
rect 54700 1028 54740 1408
rect 54604 988 54740 1028
rect 54412 944 54452 953
rect 54220 904 54412 944
rect 54220 80 54260 904
rect 54412 895 54452 904
rect 54411 356 54453 365
rect 54411 316 54412 356
rect 54452 316 54453 356
rect 54411 307 54453 316
rect 54412 80 54452 307
rect 54604 80 54644 988
rect 54796 80 54836 4087
rect 54892 3893 54932 4171
rect 55084 4136 55124 5263
rect 55372 5153 55412 5524
rect 55371 5144 55413 5153
rect 55371 5104 55372 5144
rect 55412 5104 55413 5144
rect 55371 5095 55413 5104
rect 55180 4976 55220 4987
rect 55180 4901 55220 4936
rect 55372 4976 55412 4985
rect 55179 4892 55221 4901
rect 55179 4852 55180 4892
rect 55220 4852 55221 4892
rect 55179 4843 55221 4852
rect 55180 4724 55220 4733
rect 55180 4145 55220 4684
rect 55372 4649 55412 4936
rect 55371 4640 55413 4649
rect 55371 4600 55372 4640
rect 55412 4600 55413 4640
rect 55371 4591 55413 4600
rect 55275 4556 55317 4565
rect 55275 4516 55276 4556
rect 55316 4516 55317 4556
rect 55275 4507 55317 4516
rect 55084 4087 55124 4096
rect 55179 4136 55221 4145
rect 55179 4096 55180 4136
rect 55220 4096 55221 4136
rect 55179 4087 55221 4096
rect 55276 4136 55316 4507
rect 55372 4136 55412 4145
rect 55468 4136 55508 5608
rect 55564 5648 55604 5657
rect 56331 5648 56373 5657
rect 55604 5608 55700 5648
rect 55564 5599 55604 5608
rect 55564 5480 55604 5489
rect 55564 5321 55604 5440
rect 55563 5312 55605 5321
rect 55563 5272 55564 5312
rect 55604 5272 55605 5312
rect 55563 5263 55605 5272
rect 55660 4565 55700 5608
rect 56331 5608 56332 5648
rect 56372 5608 56373 5648
rect 56331 5599 56373 5608
rect 56428 5648 56468 6271
rect 56620 5648 56660 5657
rect 56428 5608 56620 5648
rect 56332 5514 56372 5599
rect 56140 5480 56180 5489
rect 55852 5440 56140 5480
rect 55659 4556 55701 4565
rect 55659 4516 55660 4556
rect 55700 4516 55701 4556
rect 55659 4507 55701 4516
rect 55084 3968 55124 3977
rect 55124 3928 55220 3968
rect 55084 3919 55124 3928
rect 54891 3884 54933 3893
rect 54891 3844 54892 3884
rect 54932 3844 54933 3884
rect 54891 3835 54933 3844
rect 54892 3464 54932 3835
rect 55083 3800 55125 3809
rect 55083 3760 55084 3800
rect 55124 3760 55125 3800
rect 55083 3751 55125 3760
rect 54892 3415 54932 3424
rect 55084 3464 55124 3751
rect 55084 3415 55124 3424
rect 54987 3212 55029 3221
rect 54987 3172 54988 3212
rect 55028 3172 55029 3212
rect 54987 3163 55029 3172
rect 54988 3078 55028 3163
rect 55180 2969 55220 3928
rect 55276 3464 55316 4096
rect 55369 4096 55372 4136
rect 55412 4096 55508 4136
rect 55369 4087 55412 4096
rect 55369 3968 55409 4087
rect 55369 3928 55412 3968
rect 55372 3809 55412 3928
rect 55371 3800 55413 3809
rect 55659 3800 55701 3809
rect 55371 3760 55372 3800
rect 55412 3760 55508 3800
rect 55371 3751 55413 3760
rect 55276 3415 55316 3424
rect 55468 3464 55508 3760
rect 55659 3760 55660 3800
rect 55700 3760 55701 3800
rect 55659 3751 55701 3760
rect 55563 3716 55605 3725
rect 55563 3676 55564 3716
rect 55604 3676 55605 3716
rect 55563 3667 55605 3676
rect 55468 3415 55508 3424
rect 55372 3212 55412 3221
rect 55372 3053 55412 3172
rect 55371 3044 55413 3053
rect 55371 3004 55372 3044
rect 55412 3004 55413 3044
rect 55371 2995 55413 3004
rect 55179 2960 55221 2969
rect 55179 2920 55180 2960
rect 55220 2920 55221 2960
rect 55179 2911 55221 2920
rect 55276 2801 55316 2861
rect 55564 2801 55604 3667
rect 54892 2792 54932 2801
rect 55275 2792 55317 2801
rect 54932 2752 55220 2792
rect 54892 2743 54932 2752
rect 54891 2616 54933 2625
rect 54891 2573 54892 2616
rect 54932 2573 54933 2616
rect 54891 2567 54933 2573
rect 54892 2481 54932 2567
rect 55084 2456 55124 2465
rect 54988 2416 55084 2456
rect 54892 944 54932 953
rect 54892 533 54932 904
rect 54891 524 54933 533
rect 54891 484 54892 524
rect 54932 484 54933 524
rect 54891 475 54933 484
rect 54988 80 55028 2416
rect 55084 2407 55124 2416
rect 55083 1448 55125 1457
rect 55083 1408 55084 1448
rect 55124 1408 55125 1448
rect 55083 1399 55125 1408
rect 55084 1280 55124 1399
rect 55084 1231 55124 1240
rect 55083 1112 55125 1121
rect 55083 1072 55084 1112
rect 55124 1072 55125 1112
rect 55083 1063 55125 1072
rect 55084 978 55124 1063
rect 55180 80 55220 2752
rect 55275 2743 55276 2792
rect 55316 2743 55317 2792
rect 55563 2792 55605 2801
rect 55563 2752 55564 2792
rect 55604 2752 55605 2792
rect 55563 2743 55605 2752
rect 55276 2717 55316 2726
rect 55372 2633 55412 2644
rect 55276 2621 55316 2625
rect 55371 2624 55413 2633
rect 55371 2621 55372 2624
rect 55276 2616 55372 2621
rect 55316 2584 55372 2616
rect 55412 2584 55413 2624
rect 55316 2581 55413 2584
rect 55276 2297 55316 2576
rect 55371 2575 55413 2581
rect 55564 2456 55604 2465
rect 55275 2288 55317 2297
rect 55275 2248 55276 2288
rect 55316 2248 55317 2288
rect 55275 2239 55317 2248
rect 55371 1784 55413 1793
rect 55371 1744 55372 1784
rect 55412 1744 55413 1784
rect 55371 1735 55413 1744
rect 55275 1532 55317 1541
rect 55275 1492 55276 1532
rect 55316 1492 55317 1532
rect 55275 1483 55317 1492
rect 55276 944 55316 1483
rect 55372 1373 55412 1735
rect 55564 1709 55604 2416
rect 55563 1700 55605 1709
rect 55563 1660 55564 1700
rect 55604 1660 55605 1700
rect 55563 1651 55605 1660
rect 55371 1364 55413 1373
rect 55371 1324 55372 1364
rect 55412 1324 55413 1364
rect 55371 1315 55413 1324
rect 55372 1112 55412 1315
rect 55660 1289 55700 3751
rect 55756 2801 55796 2886
rect 55755 2792 55797 2801
rect 55755 2752 55756 2792
rect 55796 2752 55797 2792
rect 55755 2743 55797 2752
rect 55755 2624 55797 2633
rect 55755 2584 55756 2624
rect 55796 2584 55797 2624
rect 55755 2575 55797 2584
rect 55756 2490 55796 2575
rect 55852 1709 55892 5440
rect 56140 5431 56180 5440
rect 56428 5480 56468 5608
rect 56620 5599 56660 5608
rect 56811 5648 56853 5657
rect 56811 5608 56812 5648
rect 56852 5608 56853 5648
rect 56811 5599 56853 5608
rect 58156 5648 58196 5657
rect 56716 5564 56756 5573
rect 56716 5480 56756 5524
rect 56812 5514 56852 5599
rect 56428 5237 56468 5440
rect 56524 5440 56756 5480
rect 56427 5228 56469 5237
rect 56427 5188 56428 5228
rect 56468 5188 56469 5228
rect 56427 5179 56469 5188
rect 55948 4976 55988 4985
rect 55948 4817 55988 4936
rect 56140 4976 56180 4985
rect 56044 4892 56084 4901
rect 55947 4808 55989 4817
rect 55947 4768 55948 4808
rect 55988 4768 55989 4808
rect 55947 4759 55989 4768
rect 56044 3632 56084 4852
rect 55948 3592 56084 3632
rect 55851 1700 55893 1709
rect 55851 1660 55852 1700
rect 55892 1660 55893 1700
rect 55851 1651 55893 1660
rect 55755 1364 55797 1373
rect 55755 1324 55756 1364
rect 55796 1324 55797 1364
rect 55755 1315 55797 1324
rect 55659 1280 55701 1289
rect 55659 1240 55660 1280
rect 55700 1240 55701 1280
rect 55659 1231 55701 1240
rect 55372 1063 55412 1072
rect 55563 1112 55605 1121
rect 55563 1072 55564 1112
rect 55604 1072 55605 1112
rect 55563 1063 55605 1072
rect 55564 978 55604 1063
rect 55468 944 55508 953
rect 55276 904 55412 944
rect 55372 80 55412 904
rect 55468 365 55508 904
rect 55563 776 55605 785
rect 55563 736 55564 776
rect 55604 736 55605 776
rect 55563 727 55605 736
rect 55467 356 55509 365
rect 55467 316 55468 356
rect 55508 316 55509 356
rect 55467 307 55509 316
rect 55564 80 55604 727
rect 55756 80 55796 1315
rect 55948 1280 55988 3592
rect 56140 3473 56180 4936
rect 56332 4976 56372 4985
rect 56332 4817 56372 4936
rect 56427 4976 56469 4985
rect 56427 4936 56428 4976
rect 56468 4936 56469 4976
rect 56427 4927 56469 4936
rect 56428 4842 56468 4927
rect 56331 4808 56373 4817
rect 56331 4768 56332 4808
rect 56372 4768 56373 4808
rect 56331 4759 56373 4768
rect 56524 4052 56564 5440
rect 58059 5312 58101 5321
rect 58059 5272 58060 5312
rect 58100 5272 58101 5312
rect 58059 5263 58101 5272
rect 56332 4012 56564 4052
rect 56620 5144 56660 5153
rect 56139 3464 56181 3473
rect 56139 3424 56140 3464
rect 56180 3424 56181 3464
rect 56139 3415 56181 3424
rect 56043 2792 56085 2801
rect 56043 2752 56044 2792
rect 56084 2752 56085 2792
rect 56043 2743 56085 2752
rect 56044 2624 56084 2743
rect 56044 2575 56084 2584
rect 56235 2624 56277 2633
rect 56235 2584 56236 2624
rect 56276 2584 56277 2624
rect 56235 2575 56277 2584
rect 56236 2490 56276 2575
rect 56140 2456 56180 2465
rect 55852 1240 55988 1280
rect 56044 2416 56140 2456
rect 55852 533 55892 1240
rect 55947 1112 55989 1121
rect 55947 1072 55948 1112
rect 55988 1072 55989 1112
rect 55947 1063 55989 1072
rect 55851 524 55893 533
rect 55851 484 55852 524
rect 55892 484 55893 524
rect 55851 475 55893 484
rect 55948 80 55988 1063
rect 56044 785 56084 2416
rect 56140 2407 56180 2416
rect 56235 1700 56277 1709
rect 56235 1660 56236 1700
rect 56276 1660 56277 1700
rect 56235 1651 56277 1660
rect 56139 1280 56181 1289
rect 56139 1240 56140 1280
rect 56180 1240 56181 1280
rect 56139 1231 56181 1240
rect 56043 776 56085 785
rect 56043 736 56044 776
rect 56084 736 56085 776
rect 56043 727 56085 736
rect 56140 80 56180 1231
rect 56236 1112 56276 1651
rect 56332 1373 56372 4012
rect 56620 3809 56660 5104
rect 58060 5144 58100 5263
rect 58060 5095 58100 5104
rect 58156 5069 58196 5608
rect 58348 5648 58388 5657
rect 60940 5648 60980 9920
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 71884 5657 71924 9920
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 61228 5648 61268 5657
rect 60940 5608 61076 5648
rect 58252 5480 58292 5489
rect 58155 5060 58197 5069
rect 58155 5020 58156 5060
rect 58196 5020 58197 5060
rect 58155 5011 58197 5020
rect 57964 4976 58004 4985
rect 57772 4724 57812 4733
rect 57676 4684 57772 4724
rect 57099 4136 57141 4145
rect 57099 4096 57100 4136
rect 57140 4096 57141 4136
rect 57099 4087 57141 4096
rect 56619 3800 56661 3809
rect 56619 3760 56620 3800
rect 56660 3760 56661 3800
rect 56619 3751 56661 3760
rect 56620 3473 56660 3558
rect 56619 3464 56661 3473
rect 56619 3424 56620 3464
rect 56660 3424 56661 3464
rect 56619 3415 56661 3424
rect 56908 3464 56948 3475
rect 57100 3473 57140 4087
rect 57676 3641 57716 4684
rect 57772 4675 57812 4684
rect 57964 4565 58004 4936
rect 58060 4976 58100 4985
rect 58060 4817 58100 4936
rect 58059 4808 58101 4817
rect 58059 4768 58060 4808
rect 58100 4768 58101 4808
rect 58059 4759 58101 4768
rect 57963 4556 58005 4565
rect 57963 4516 57964 4556
rect 58004 4516 58005 4556
rect 57963 4507 58005 4516
rect 57675 3632 57717 3641
rect 57675 3592 57676 3632
rect 57716 3592 57717 3632
rect 57675 3583 57717 3592
rect 57867 3632 57909 3641
rect 57867 3592 57868 3632
rect 57908 3592 57909 3632
rect 57867 3583 57909 3592
rect 57099 3464 57141 3473
rect 56908 3389 56948 3424
rect 57004 3424 57100 3464
rect 57140 3424 57141 3464
rect 56907 3380 56949 3389
rect 56907 3340 56908 3380
rect 56948 3340 56949 3380
rect 56907 3331 56949 3340
rect 56619 3296 56661 3305
rect 56619 3256 56620 3296
rect 56660 3256 56661 3296
rect 56619 3247 56661 3256
rect 56428 3212 56468 3221
rect 56428 2540 56468 3172
rect 56620 3162 56660 3247
rect 56908 3212 56948 3221
rect 56428 2500 56564 2540
rect 56331 1364 56373 1373
rect 56331 1324 56332 1364
rect 56372 1324 56373 1364
rect 56331 1315 56373 1324
rect 56427 1196 56469 1205
rect 56427 1156 56428 1196
rect 56468 1156 56469 1196
rect 56427 1147 56469 1156
rect 56236 1063 56276 1072
rect 56428 1112 56468 1147
rect 56428 1061 56468 1072
rect 56332 944 56372 953
rect 56332 785 56372 904
rect 56331 776 56373 785
rect 56331 736 56332 776
rect 56372 736 56373 776
rect 56331 727 56373 736
rect 56331 524 56373 533
rect 56331 484 56332 524
rect 56372 484 56373 524
rect 56331 475 56373 484
rect 56332 80 56372 475
rect 56524 80 56564 2500
rect 56716 1289 56756 1374
rect 56715 1280 56757 1289
rect 56715 1240 56716 1280
rect 56756 1240 56757 1280
rect 56715 1231 56757 1240
rect 56619 1115 56661 1121
rect 56716 1115 56756 1124
rect 56619 1112 56716 1115
rect 56619 1072 56620 1112
rect 56660 1075 56716 1112
rect 56908 1113 56948 3172
rect 57004 2129 57044 3424
rect 57099 3415 57141 3424
rect 57100 3330 57140 3415
rect 57676 2969 57716 3583
rect 57868 3296 57908 3583
rect 57964 3473 58004 4507
rect 57963 3464 58005 3473
rect 57963 3424 57964 3464
rect 58004 3424 58005 3464
rect 58060 3464 58100 4759
rect 58156 4304 58196 5011
rect 58156 4255 58196 4264
rect 58155 4136 58197 4145
rect 58155 4096 58156 4136
rect 58196 4096 58197 4136
rect 58155 4087 58197 4096
rect 58156 4002 58196 4087
rect 58156 3464 58196 3473
rect 58060 3424 58156 3464
rect 57963 3415 58005 3424
rect 58156 3415 58196 3424
rect 58252 3389 58292 5440
rect 58348 4145 58388 5608
rect 58827 5564 58869 5573
rect 58827 5524 58828 5564
rect 58868 5524 58869 5564
rect 58827 5515 58869 5524
rect 58731 5312 58773 5321
rect 58731 5272 58732 5312
rect 58772 5272 58773 5312
rect 58731 5263 58773 5272
rect 58732 5144 58772 5263
rect 58732 5095 58772 5104
rect 58636 4976 58676 4985
rect 58539 4808 58581 4817
rect 58539 4768 58540 4808
rect 58580 4768 58581 4808
rect 58539 4759 58581 4768
rect 58443 4724 58485 4733
rect 58443 4684 58444 4724
rect 58484 4684 58485 4724
rect 58443 4675 58485 4684
rect 58444 4590 58484 4675
rect 58347 4136 58389 4145
rect 58347 4096 58348 4136
rect 58388 4096 58389 4136
rect 58347 4087 58389 4096
rect 58540 4136 58580 4759
rect 58636 4220 58676 4936
rect 58732 4976 58772 4985
rect 58828 4976 58868 5515
rect 61036 5489 61076 5608
rect 61131 5564 61173 5573
rect 61131 5524 61132 5564
rect 61172 5524 61173 5564
rect 61131 5515 61173 5524
rect 60940 5480 60980 5489
rect 58923 5312 58965 5321
rect 58923 5272 58924 5312
rect 58964 5272 58965 5312
rect 58923 5263 58965 5272
rect 58772 4936 58868 4976
rect 58732 4817 58772 4936
rect 58731 4808 58773 4817
rect 58731 4768 58732 4808
rect 58772 4768 58773 4808
rect 58731 4759 58773 4768
rect 58636 4180 58772 4220
rect 58348 3968 58388 3977
rect 58348 3809 58388 3928
rect 58347 3800 58389 3809
rect 58540 3800 58580 4096
rect 58732 4136 58772 4180
rect 58347 3760 58348 3800
rect 58388 3760 58389 3800
rect 58347 3751 58389 3760
rect 58537 3760 58580 3800
rect 58636 4052 58676 4061
rect 58348 3473 58388 3558
rect 58537 3548 58577 3760
rect 58636 3725 58676 4012
rect 58732 3893 58772 4096
rect 58731 3884 58773 3893
rect 58731 3844 58732 3884
rect 58772 3844 58773 3884
rect 58731 3835 58773 3844
rect 58635 3716 58677 3725
rect 58635 3676 58636 3716
rect 58676 3676 58677 3716
rect 58635 3667 58677 3676
rect 58537 3508 58676 3548
rect 58347 3464 58389 3473
rect 58636 3464 58676 3508
rect 58924 3473 58964 5263
rect 60459 5144 60501 5153
rect 60459 5104 60460 5144
rect 60500 5104 60501 5144
rect 60459 5095 60501 5104
rect 60460 4976 60500 5095
rect 60364 4936 60460 4976
rect 59115 4724 59157 4733
rect 59115 4684 59116 4724
rect 59156 4684 59157 4724
rect 59115 4675 59157 4684
rect 59020 4313 59060 4398
rect 59019 4304 59061 4313
rect 59019 4264 59020 4304
rect 59060 4264 59061 4304
rect 59019 4255 59061 4264
rect 59019 4136 59061 4145
rect 59019 4096 59020 4136
rect 59060 4096 59061 4136
rect 59019 4087 59061 4096
rect 59020 4002 59060 4087
rect 59019 3884 59061 3893
rect 59019 3844 59020 3884
rect 59060 3844 59061 3884
rect 59019 3835 59061 3844
rect 58347 3424 58348 3464
rect 58388 3451 58580 3464
rect 58388 3424 58540 3451
rect 58347 3415 58389 3424
rect 58540 3402 58580 3411
rect 58636 3389 58676 3424
rect 58828 3464 58868 3473
rect 58923 3464 58965 3473
rect 58868 3424 58924 3464
rect 58964 3424 58965 3464
rect 58828 3415 58868 3424
rect 58923 3415 58965 3424
rect 59020 3464 59060 3835
rect 59116 3641 59156 4675
rect 59403 4304 59445 4313
rect 59403 4264 59404 4304
rect 59444 4264 59445 4304
rect 59403 4255 59445 4264
rect 59404 4136 59444 4255
rect 60364 4145 60404 4936
rect 60460 4927 60500 4936
rect 60843 4976 60885 4985
rect 60843 4936 60844 4976
rect 60884 4936 60885 4976
rect 60843 4927 60885 4936
rect 60844 4842 60884 4927
rect 60459 4808 60501 4817
rect 60459 4768 60460 4808
rect 60500 4768 60501 4808
rect 60459 4759 60501 4768
rect 60460 4674 60500 4759
rect 60652 4724 60692 4733
rect 60844 4724 60884 4733
rect 60692 4684 60788 4724
rect 60652 4675 60692 4684
rect 59404 4087 59444 4096
rect 59595 4136 59637 4145
rect 59595 4096 59596 4136
rect 59636 4096 59637 4136
rect 59595 4087 59637 4096
rect 60363 4136 60405 4145
rect 60363 4096 60364 4136
rect 60404 4096 60405 4136
rect 60363 4087 60405 4096
rect 59596 4002 59636 4087
rect 59212 3968 59252 3977
rect 59500 3968 59540 3977
rect 59115 3632 59157 3641
rect 59115 3592 59116 3632
rect 59156 3592 59157 3632
rect 59115 3583 59157 3592
rect 59020 3415 59060 3424
rect 59116 3464 59156 3475
rect 58251 3380 58293 3389
rect 58251 3340 58252 3380
rect 58292 3340 58293 3380
rect 58251 3331 58293 3340
rect 58635 3380 58677 3389
rect 58635 3340 58636 3380
rect 58676 3340 58677 3380
rect 58635 3331 58677 3340
rect 58539 3296 58581 3305
rect 58636 3300 58676 3331
rect 58924 3330 58964 3415
rect 59116 3389 59156 3424
rect 59115 3380 59157 3389
rect 59115 3340 59116 3380
rect 59156 3340 59157 3380
rect 59115 3331 59157 3340
rect 57868 3256 58004 3296
rect 57675 2960 57717 2969
rect 57675 2920 57676 2960
rect 57716 2920 57717 2960
rect 57675 2911 57717 2920
rect 57964 2885 58004 3256
rect 58539 3256 58540 3296
rect 58580 3256 58581 3296
rect 58539 3247 58581 3256
rect 58252 3212 58292 3221
rect 57963 2876 58005 2885
rect 57963 2836 57964 2876
rect 58004 2836 58005 2876
rect 57963 2827 58005 2836
rect 58252 2801 58292 3172
rect 58251 2792 58293 2801
rect 58251 2752 58252 2792
rect 58292 2752 58293 2792
rect 58251 2743 58293 2752
rect 58540 2372 58580 3247
rect 58828 3212 58868 3221
rect 58868 3172 59156 3212
rect 58828 3163 58868 3172
rect 58636 2792 58676 2801
rect 58676 2752 59060 2792
rect 58636 2743 58676 2752
rect 58635 2624 58677 2633
rect 58635 2584 58636 2624
rect 58676 2584 58677 2624
rect 58635 2575 58677 2584
rect 58923 2624 58965 2633
rect 58923 2584 58924 2624
rect 58964 2584 58965 2624
rect 58923 2575 58965 2584
rect 58636 2490 58676 2575
rect 58828 2456 58868 2465
rect 58540 2332 58676 2372
rect 57003 2120 57045 2129
rect 57003 2080 57004 2120
rect 57044 2080 57045 2120
rect 57003 2071 57045 2080
rect 57483 2120 57525 2129
rect 57483 2080 57484 2120
rect 57524 2080 57525 2120
rect 57483 2071 57525 2080
rect 58059 2120 58101 2129
rect 58059 2080 58060 2120
rect 58100 2080 58101 2120
rect 58059 2071 58101 2080
rect 57004 1952 57044 2071
rect 57387 2036 57429 2045
rect 57387 1996 57388 2036
rect 57428 1996 57429 2036
rect 57387 1987 57429 1996
rect 57004 1709 57044 1912
rect 57196 1952 57236 1963
rect 57196 1877 57236 1912
rect 57195 1868 57237 1877
rect 57100 1828 57196 1868
rect 57236 1828 57237 1868
rect 57003 1700 57045 1709
rect 57003 1660 57004 1700
rect 57044 1660 57045 1700
rect 57003 1651 57045 1660
rect 56660 1072 56661 1075
rect 56619 1063 56661 1072
rect 56716 1066 56756 1075
rect 56813 1073 56948 1113
rect 57004 1115 57044 1651
rect 57100 1532 57140 1828
rect 57195 1819 57237 1828
rect 57388 1784 57428 1987
rect 57484 1952 57524 2071
rect 57867 2036 57909 2045
rect 57867 1996 57868 2036
rect 57908 1996 57909 2036
rect 57867 1987 57909 1996
rect 57484 1903 57524 1912
rect 57868 1952 57908 1987
rect 57868 1901 57908 1912
rect 58060 1952 58100 2071
rect 58443 2036 58485 2045
rect 58443 1996 58444 2036
rect 58484 1996 58485 2036
rect 58443 1987 58485 1996
rect 58060 1903 58100 1912
rect 57484 1784 57524 1793
rect 57388 1744 57484 1784
rect 57484 1735 57524 1744
rect 57196 1700 57236 1709
rect 57676 1700 57716 1709
rect 57236 1660 57428 1700
rect 57196 1651 57236 1660
rect 57100 1492 57236 1532
rect 57196 1280 57236 1492
rect 57196 1231 57236 1240
rect 57099 1115 57141 1121
rect 57196 1115 57236 1121
rect 57004 1112 57236 1115
rect 57004 1075 57100 1112
rect 56813 1028 56853 1073
rect 57099 1072 57100 1075
rect 57140 1075 57196 1112
rect 57140 1072 57141 1075
rect 57099 1063 57141 1072
rect 57388 1112 57428 1660
rect 57388 1072 57524 1112
rect 57196 1063 57236 1072
rect 56812 988 56853 1028
rect 56812 776 56852 988
rect 56716 736 56852 776
rect 56908 944 56948 953
rect 57100 951 57140 1063
rect 57388 944 57428 953
rect 56716 80 56756 736
rect 56908 80 56948 904
rect 57292 904 57388 944
rect 57099 776 57141 785
rect 57099 736 57100 776
rect 57140 736 57141 776
rect 57099 727 57141 736
rect 57100 80 57140 727
rect 57292 80 57332 904
rect 57388 895 57428 904
rect 57484 80 57524 1072
rect 57676 80 57716 1660
rect 57868 1700 57908 1709
rect 57771 1448 57813 1457
rect 57771 1408 57772 1448
rect 57812 1408 57813 1448
rect 57771 1399 57813 1408
rect 57772 1280 57812 1399
rect 57772 1231 57812 1240
rect 57771 1112 57813 1121
rect 57771 1072 57772 1112
rect 57812 1072 57813 1112
rect 57771 1063 57813 1072
rect 57772 978 57812 1063
rect 57868 80 57908 1660
rect 58155 1448 58197 1457
rect 58155 1408 58156 1448
rect 58196 1408 58197 1448
rect 58155 1399 58197 1408
rect 58156 1112 58196 1399
rect 58156 1063 58196 1072
rect 58347 1112 58389 1121
rect 58347 1072 58348 1112
rect 58388 1072 58389 1112
rect 58347 1063 58389 1072
rect 58348 978 58388 1063
rect 57964 944 58004 953
rect 58252 944 58292 953
rect 58004 904 58100 944
rect 57964 895 58004 904
rect 58060 80 58100 904
rect 58252 80 58292 904
rect 58444 80 58484 1987
rect 58636 80 58676 2332
rect 58731 1952 58773 1961
rect 58731 1912 58732 1952
rect 58772 1912 58773 1952
rect 58731 1903 58773 1912
rect 58732 1818 58772 1903
rect 58731 1700 58773 1709
rect 58731 1660 58732 1700
rect 58772 1660 58773 1700
rect 58731 1651 58773 1660
rect 58732 1566 58772 1651
rect 58828 80 58868 2416
rect 58924 1961 58964 2575
rect 59020 2129 59060 2752
rect 59116 2465 59156 3172
rect 59115 2456 59157 2465
rect 59115 2416 59116 2456
rect 59156 2416 59157 2456
rect 59115 2407 59157 2416
rect 59019 2120 59061 2129
rect 59019 2080 59020 2120
rect 59060 2080 59061 2120
rect 59019 2071 59061 2080
rect 58923 1952 58965 1961
rect 58923 1912 58924 1952
rect 58964 1912 58965 1952
rect 58923 1903 58965 1912
rect 58924 1818 58964 1903
rect 59019 1700 59061 1709
rect 59019 1660 59020 1700
rect 59060 1660 59061 1700
rect 59019 1651 59061 1660
rect 59020 80 59060 1651
rect 59115 1112 59157 1121
rect 59115 1072 59116 1112
rect 59156 1072 59157 1112
rect 59115 1063 59157 1072
rect 59116 978 59156 1063
rect 59212 80 59252 3928
rect 59404 3928 59500 3968
rect 59307 3464 59349 3473
rect 59307 3424 59308 3464
rect 59348 3424 59349 3464
rect 59307 3415 59349 3424
rect 59308 3330 59348 3415
rect 59308 3212 59348 3221
rect 59308 1709 59348 3172
rect 59307 1700 59349 1709
rect 59307 1660 59308 1700
rect 59348 1660 59349 1700
rect 59307 1651 59349 1660
rect 59308 1289 59348 1374
rect 59307 1280 59349 1289
rect 59307 1240 59308 1280
rect 59348 1240 59349 1280
rect 59307 1231 59349 1240
rect 59308 1112 59348 1121
rect 59308 953 59348 1072
rect 59307 944 59349 953
rect 59307 904 59308 944
rect 59348 904 59349 944
rect 59307 895 59349 904
rect 59404 80 59444 3928
rect 59500 3919 59540 3928
rect 60651 3716 60693 3725
rect 60651 3676 60652 3716
rect 60692 3676 60693 3716
rect 60651 3667 60693 3676
rect 60652 2885 60692 3667
rect 60651 2876 60693 2885
rect 60651 2836 60652 2876
rect 60692 2836 60693 2876
rect 60651 2827 60693 2836
rect 60459 2624 60501 2633
rect 60459 2584 60460 2624
rect 60500 2584 60501 2624
rect 60459 2575 60501 2584
rect 60652 2624 60692 2827
rect 60652 2575 60692 2584
rect 60460 1961 60500 2575
rect 60555 2456 60597 2465
rect 60555 2416 60556 2456
rect 60596 2416 60597 2456
rect 60555 2407 60597 2416
rect 60556 2322 60596 2407
rect 59979 1952 60021 1961
rect 59979 1912 59980 1952
rect 60020 1912 60021 1952
rect 59979 1903 60021 1912
rect 60172 1952 60212 1961
rect 59980 1818 60020 1903
rect 60076 1868 60116 1877
rect 59499 1616 59541 1625
rect 59499 1576 59500 1616
rect 59540 1576 59541 1616
rect 59499 1567 59541 1576
rect 59500 1280 59540 1567
rect 59596 1280 59636 1289
rect 59500 1240 59596 1280
rect 59500 953 59540 1240
rect 59596 1231 59636 1240
rect 59883 1280 59925 1289
rect 59883 1240 59884 1280
rect 59924 1240 59925 1280
rect 59883 1231 59925 1240
rect 59595 1112 59637 1121
rect 59595 1072 59596 1112
rect 59636 1072 59637 1112
rect 59595 1063 59637 1072
rect 59596 978 59636 1063
rect 59499 944 59541 953
rect 59788 944 59828 953
rect 59499 904 59500 944
rect 59540 904 59541 944
rect 59499 895 59541 904
rect 59692 904 59788 944
rect 59692 524 59732 904
rect 59788 895 59828 904
rect 59884 524 59924 1231
rect 59596 484 59732 524
rect 59788 484 59924 524
rect 59980 944 60020 953
rect 59596 80 59636 484
rect 59788 80 59828 484
rect 59980 80 60020 904
rect 60076 860 60116 1828
rect 60172 1541 60212 1912
rect 60459 1952 60501 1961
rect 60459 1912 60460 1952
rect 60500 1912 60501 1952
rect 60459 1903 60501 1912
rect 60651 1784 60693 1793
rect 60651 1744 60652 1784
rect 60692 1744 60693 1784
rect 60651 1735 60693 1744
rect 60267 1700 60309 1709
rect 60267 1660 60268 1700
rect 60308 1660 60309 1700
rect 60267 1651 60309 1660
rect 60171 1532 60213 1541
rect 60171 1492 60172 1532
rect 60212 1492 60213 1532
rect 60171 1483 60213 1492
rect 60172 1280 60212 1483
rect 60172 1231 60212 1240
rect 60171 1112 60213 1121
rect 60171 1072 60172 1112
rect 60212 1072 60213 1112
rect 60171 1063 60213 1072
rect 60172 978 60212 1063
rect 60076 820 60212 860
rect 60172 80 60212 820
rect 60268 197 60308 1651
rect 60652 1289 60692 1735
rect 60651 1280 60693 1289
rect 60651 1240 60652 1280
rect 60692 1240 60693 1280
rect 60651 1231 60693 1240
rect 60651 1112 60693 1121
rect 60651 1072 60652 1112
rect 60692 1072 60693 1112
rect 60651 1063 60693 1072
rect 60652 978 60692 1063
rect 60460 944 60500 953
rect 60364 904 60460 944
rect 60267 188 60309 197
rect 60267 148 60268 188
rect 60308 148 60309 188
rect 60267 139 60309 148
rect 60364 80 60404 904
rect 60460 895 60500 904
rect 60555 944 60597 953
rect 60555 904 60556 944
rect 60596 904 60597 944
rect 60555 895 60597 904
rect 60556 80 60596 895
rect 60748 80 60788 4684
rect 60844 944 60884 4684
rect 60940 4649 60980 5440
rect 61035 5480 61077 5489
rect 61035 5440 61036 5480
rect 61076 5440 61077 5480
rect 61035 5431 61077 5440
rect 61036 5346 61076 5431
rect 61132 5430 61172 5515
rect 61228 5321 61268 5608
rect 61324 5648 61364 5657
rect 61227 5312 61269 5321
rect 61227 5272 61228 5312
rect 61268 5272 61269 5312
rect 61227 5263 61269 5272
rect 61035 5144 61077 5153
rect 61035 5104 61036 5144
rect 61076 5104 61077 5144
rect 61035 5095 61077 5104
rect 61036 4976 61076 5095
rect 61324 4985 61364 5608
rect 61515 5648 61557 5657
rect 61515 5608 61516 5648
rect 61556 5608 61557 5648
rect 61515 5599 61557 5608
rect 61708 5648 61748 5657
rect 61516 5480 61556 5599
rect 61516 5431 61556 5440
rect 61515 5312 61557 5321
rect 61515 5272 61516 5312
rect 61556 5272 61557 5312
rect 61515 5263 61557 5272
rect 61419 5228 61461 5237
rect 61419 5188 61420 5228
rect 61460 5188 61461 5228
rect 61419 5179 61461 5188
rect 61036 4733 61076 4936
rect 61228 4976 61268 4985
rect 61228 4901 61268 4936
rect 61323 4976 61365 4985
rect 61323 4936 61324 4976
rect 61364 4936 61365 4976
rect 61323 4927 61365 4936
rect 61227 4892 61269 4901
rect 61227 4852 61228 4892
rect 61268 4852 61269 4892
rect 61227 4843 61269 4852
rect 61035 4724 61077 4733
rect 61035 4684 61036 4724
rect 61076 4684 61077 4724
rect 61035 4675 61077 4684
rect 60939 4640 60981 4649
rect 60939 4600 60940 4640
rect 60980 4600 60981 4640
rect 60939 4591 60981 4600
rect 61228 4061 61268 4843
rect 61324 4842 61364 4927
rect 61323 4724 61365 4733
rect 61323 4684 61324 4724
rect 61364 4684 61365 4724
rect 61323 4675 61365 4684
rect 61324 4590 61364 4675
rect 61420 4136 61460 5179
rect 61516 4976 61556 5263
rect 61708 4985 61748 5608
rect 61804 5648 61844 5657
rect 61804 5312 61844 5608
rect 61899 5648 61941 5657
rect 61899 5608 61900 5648
rect 61940 5608 61941 5648
rect 61899 5599 61941 5608
rect 61996 5648 62036 5657
rect 61900 5514 61940 5599
rect 61996 5489 62036 5608
rect 62571 5648 62613 5657
rect 62571 5608 62572 5648
rect 62612 5608 62613 5648
rect 62571 5599 62613 5608
rect 71883 5648 71925 5657
rect 71883 5608 71884 5648
rect 71924 5608 71925 5648
rect 71883 5599 71925 5608
rect 73323 5648 73365 5657
rect 73323 5608 73324 5648
rect 73364 5608 73365 5648
rect 73323 5599 73365 5608
rect 61995 5480 62037 5489
rect 61995 5440 61996 5480
rect 62036 5440 62037 5480
rect 61995 5431 62037 5440
rect 62379 5480 62421 5489
rect 62379 5440 62380 5480
rect 62420 5440 62421 5480
rect 62379 5431 62421 5440
rect 61899 5312 61941 5321
rect 61804 5272 61900 5312
rect 61940 5272 61941 5312
rect 61899 5263 61941 5272
rect 61900 5144 61940 5263
rect 61900 5095 61940 5104
rect 61803 5060 61845 5069
rect 61803 5020 61804 5060
rect 61844 5020 61845 5060
rect 61803 5011 61845 5020
rect 62187 5060 62229 5069
rect 62187 5020 62188 5060
rect 62228 5020 62229 5060
rect 62187 5011 62229 5020
rect 61707 4976 61749 4985
rect 61556 4936 61652 4976
rect 61516 4927 61556 4936
rect 61516 4136 61556 4145
rect 61420 4096 61516 4136
rect 61227 4052 61269 4061
rect 61227 4012 61228 4052
rect 61268 4012 61269 4052
rect 61227 4003 61269 4012
rect 61516 3977 61556 4096
rect 61324 3968 61364 3977
rect 60939 2876 60981 2885
rect 60939 2836 60940 2876
rect 60980 2836 60981 2876
rect 60939 2827 60981 2836
rect 60940 2792 60980 2827
rect 60940 2741 60980 2752
rect 61324 2717 61364 3928
rect 61515 3968 61557 3977
rect 61515 3928 61516 3968
rect 61556 3928 61557 3968
rect 61515 3919 61557 3928
rect 61612 3968 61652 4936
rect 61707 4936 61708 4976
rect 61748 4936 61749 4976
rect 61707 4927 61749 4936
rect 61804 4136 61844 5011
rect 61899 4976 61941 4985
rect 61899 4936 61900 4976
rect 61940 4936 61941 4976
rect 61899 4927 61941 4936
rect 61996 4976 62036 4985
rect 61900 4808 61940 4927
rect 61996 4892 62036 4936
rect 62188 4926 62228 5011
rect 62380 4976 62420 5431
rect 62572 4976 62612 5599
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 73324 4985 73364 5599
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 82156 4985 82196 5070
rect 62420 4936 62516 4976
rect 62380 4927 62420 4936
rect 62091 4892 62133 4901
rect 61996 4852 62092 4892
rect 62132 4852 62133 4892
rect 62091 4843 62133 4852
rect 61900 4768 62036 4808
rect 61899 4136 61941 4145
rect 61804 4096 61900 4136
rect 61940 4096 61941 4136
rect 61899 4087 61941 4096
rect 61900 4002 61940 4087
rect 61996 3977 62036 4768
rect 62092 4565 62132 4843
rect 62379 4724 62421 4733
rect 62379 4684 62380 4724
rect 62420 4684 62421 4724
rect 62379 4675 62421 4684
rect 62380 4590 62420 4675
rect 62091 4556 62133 4565
rect 62091 4516 62092 4556
rect 62132 4516 62133 4556
rect 62091 4507 62133 4516
rect 62476 4313 62516 4936
rect 62572 4927 62612 4936
rect 62667 4976 62709 4985
rect 62667 4936 62668 4976
rect 62708 4936 62709 4976
rect 62667 4927 62709 4936
rect 66892 4976 66932 4985
rect 62668 4481 62708 4927
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 62667 4472 62709 4481
rect 62667 4432 62668 4472
rect 62708 4432 62709 4472
rect 62667 4423 62709 4432
rect 66892 4397 66932 4936
rect 67179 4976 67221 4985
rect 67179 4936 67180 4976
rect 67220 4936 67221 4976
rect 67179 4927 67221 4936
rect 73323 4976 73365 4985
rect 73323 4936 73324 4976
rect 73364 4936 73365 4976
rect 73323 4927 73365 4936
rect 73612 4976 73652 4985
rect 67180 4842 67220 4927
rect 69099 4808 69141 4817
rect 69099 4768 69100 4808
rect 69140 4768 69141 4808
rect 69099 4759 69141 4768
rect 67180 4724 67220 4733
rect 66891 4388 66933 4397
rect 66891 4348 66892 4388
rect 66932 4348 66933 4388
rect 66891 4339 66933 4348
rect 62475 4304 62517 4313
rect 62475 4264 62476 4304
rect 62516 4264 62517 4304
rect 62475 4255 62517 4264
rect 62284 4136 62324 4147
rect 62284 4061 62324 4096
rect 62475 4136 62517 4145
rect 62475 4096 62476 4136
rect 62516 4096 62517 4136
rect 62475 4087 62517 4096
rect 66507 4136 66549 4145
rect 66507 4096 66508 4136
rect 66548 4096 66549 4136
rect 66507 4087 66549 4096
rect 66796 4136 66836 4145
rect 62283 4052 62325 4061
rect 62283 4012 62284 4052
rect 62324 4012 62325 4052
rect 62283 4003 62325 4012
rect 62380 4052 62420 4061
rect 61612 3464 61652 3928
rect 61803 3968 61845 3977
rect 61803 3928 61804 3968
rect 61844 3928 61845 3968
rect 61803 3919 61845 3928
rect 61995 3968 62037 3977
rect 61995 3928 61996 3968
rect 62036 3928 62037 3968
rect 61995 3919 62037 3928
rect 62092 3968 62132 3977
rect 61612 3415 61652 3424
rect 61804 3464 61844 3919
rect 61804 3415 61844 3424
rect 61708 3212 61748 3221
rect 61420 2801 61460 2886
rect 61419 2792 61461 2801
rect 61419 2752 61420 2792
rect 61460 2752 61461 2792
rect 61419 2743 61461 2752
rect 61323 2708 61365 2717
rect 61323 2668 61324 2708
rect 61364 2668 61365 2708
rect 61323 2659 61365 2668
rect 61708 2633 61748 3172
rect 61803 2792 61845 2801
rect 61803 2752 61804 2792
rect 61844 2752 61845 2792
rect 61803 2743 61845 2752
rect 60939 2624 60981 2633
rect 60939 2584 60940 2624
rect 60980 2584 60981 2624
rect 60939 2575 60981 2584
rect 61419 2624 61461 2633
rect 61419 2584 61420 2624
rect 61460 2584 61461 2624
rect 61419 2575 61461 2584
rect 61707 2624 61749 2633
rect 61707 2584 61708 2624
rect 61748 2584 61749 2624
rect 61707 2575 61749 2584
rect 61804 2624 61844 2743
rect 61995 2708 62037 2717
rect 61995 2668 61996 2708
rect 62036 2668 62037 2708
rect 61995 2659 62037 2668
rect 61804 2575 61844 2584
rect 61996 2624 62036 2659
rect 60940 2490 60980 2575
rect 61420 2490 61460 2575
rect 61996 2573 62036 2584
rect 61132 2456 61172 2465
rect 61323 2456 61365 2465
rect 61612 2456 61652 2465
rect 61900 2456 61940 2465
rect 61172 2416 61268 2456
rect 61132 2407 61172 2416
rect 60939 1280 60981 1289
rect 60939 1240 60940 1280
rect 60980 1240 60981 1280
rect 60939 1231 60981 1240
rect 60940 1112 60980 1231
rect 61132 1121 61172 1206
rect 60940 1063 60980 1072
rect 61131 1112 61173 1121
rect 61131 1072 61132 1112
rect 61172 1072 61173 1112
rect 61131 1063 61173 1072
rect 61035 944 61077 953
rect 61228 944 61268 2416
rect 61323 2416 61324 2456
rect 61364 2416 61365 2456
rect 61323 2407 61365 2416
rect 61516 2416 61612 2456
rect 60844 904 60980 944
rect 60940 80 60980 904
rect 61035 904 61036 944
rect 61076 904 61077 944
rect 61035 895 61077 904
rect 61132 904 61268 944
rect 61036 810 61076 895
rect 61132 80 61172 904
rect 61324 80 61364 2407
rect 61516 80 61556 2416
rect 61612 2407 61652 2416
rect 61708 2416 61900 2456
rect 61708 80 61748 2416
rect 61900 2407 61940 2416
rect 61899 1868 61941 1877
rect 61899 1828 61900 1868
rect 61940 1828 61941 1868
rect 61899 1819 61941 1828
rect 61900 80 61940 1819
rect 62092 80 62132 3928
rect 62380 1877 62420 4012
rect 62476 4002 62516 4087
rect 66508 4002 66548 4087
rect 66796 3977 66836 4096
rect 66987 4136 67029 4145
rect 66987 4096 66988 4136
rect 67028 4096 67029 4136
rect 66987 4087 67029 4096
rect 66892 4052 66932 4061
rect 66316 3968 66356 3977
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 64011 3716 64053 3725
rect 64011 3676 64012 3716
rect 64052 3676 64053 3716
rect 64011 3667 64053 3676
rect 63147 3464 63189 3473
rect 63147 3424 63148 3464
rect 63188 3424 63189 3464
rect 63147 3415 63189 3424
rect 63340 3464 63380 3473
rect 63148 3330 63188 3415
rect 63340 3305 63380 3424
rect 63435 3464 63477 3473
rect 63435 3424 63436 3464
rect 63476 3424 63477 3464
rect 63435 3415 63477 3424
rect 63819 3464 63861 3473
rect 63819 3424 63820 3464
rect 63860 3424 63861 3464
rect 63819 3415 63861 3424
rect 64012 3464 64052 3667
rect 66316 3557 66356 3928
rect 66603 3968 66645 3977
rect 66603 3928 66604 3968
rect 66644 3928 66645 3968
rect 66603 3919 66645 3928
rect 66795 3968 66837 3977
rect 66795 3928 66796 3968
rect 66836 3928 66837 3968
rect 66795 3919 66837 3928
rect 66411 3884 66453 3893
rect 66411 3844 66412 3884
rect 66452 3844 66453 3884
rect 66411 3835 66453 3844
rect 65451 3548 65493 3557
rect 65451 3508 65452 3548
rect 65492 3508 65493 3548
rect 65451 3499 65493 3508
rect 65643 3548 65685 3557
rect 65643 3508 65644 3548
rect 65684 3508 65685 3548
rect 65643 3499 65685 3508
rect 66027 3548 66069 3557
rect 66027 3508 66028 3548
rect 66068 3508 66069 3548
rect 66027 3499 66069 3508
rect 66315 3548 66357 3557
rect 66315 3508 66316 3548
rect 66356 3508 66357 3548
rect 66315 3499 66357 3508
rect 64203 3464 64245 3473
rect 64052 3424 64148 3464
rect 64012 3415 64052 3424
rect 63339 3296 63381 3305
rect 63339 3256 63340 3296
rect 63380 3256 63381 3296
rect 63339 3247 63381 3256
rect 63244 3212 63284 3221
rect 63148 3172 63244 3212
rect 62859 2792 62901 2801
rect 62859 2752 62860 2792
rect 62900 2752 62901 2792
rect 62859 2743 62901 2752
rect 62860 2624 62900 2743
rect 63052 2633 63092 2718
rect 62860 2540 62900 2584
rect 63051 2624 63093 2633
rect 63051 2584 63052 2624
rect 63092 2584 63093 2624
rect 63051 2575 63093 2584
rect 62764 2500 62900 2540
rect 62956 2540 62996 2549
rect 62571 1952 62613 1961
rect 62571 1912 62572 1952
rect 62612 1912 62613 1952
rect 62571 1903 62613 1912
rect 62764 1952 62804 2500
rect 62764 1903 62804 1912
rect 62379 1868 62421 1877
rect 62379 1828 62380 1868
rect 62420 1828 62421 1868
rect 62379 1819 62421 1828
rect 62572 1818 62612 1903
rect 62668 1700 62708 1709
rect 62284 1660 62668 1700
rect 62284 80 62324 1660
rect 62668 1651 62708 1660
rect 62956 1364 62996 2500
rect 63052 1373 63092 1458
rect 62572 1324 62996 1364
rect 63051 1364 63093 1373
rect 63051 1324 63052 1364
rect 63092 1324 63093 1364
rect 62475 944 62517 953
rect 62475 904 62476 944
rect 62516 904 62517 944
rect 62475 895 62517 904
rect 62476 80 62516 895
rect 62572 860 62612 1324
rect 63051 1315 63093 1324
rect 62668 1121 62708 1206
rect 63051 1196 63093 1205
rect 63051 1156 63052 1196
rect 63092 1156 63093 1196
rect 63051 1147 63093 1156
rect 62667 1112 62709 1121
rect 62667 1072 62668 1112
rect 62708 1072 62709 1112
rect 63052 1112 63092 1147
rect 62667 1063 62709 1072
rect 62860 1101 62900 1110
rect 63052 1061 63092 1072
rect 63148 1109 63188 3172
rect 63244 3163 63284 3172
rect 63436 3128 63476 3415
rect 63820 3330 63860 3415
rect 63916 3212 63956 3221
rect 63956 3172 64052 3212
rect 63916 3163 63956 3172
rect 63340 3088 63476 3128
rect 63340 2801 63380 3088
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 63339 2792 63381 2801
rect 63339 2752 63340 2792
rect 63380 2752 63381 2792
rect 63339 2743 63381 2752
rect 63340 2624 63380 2743
rect 63532 2633 63572 2718
rect 63340 2575 63380 2584
rect 63531 2624 63573 2633
rect 63531 2584 63532 2624
rect 63572 2584 63573 2624
rect 63531 2575 63573 2584
rect 63436 2540 63476 2549
rect 63436 1280 63476 2500
rect 64012 1709 64052 3172
rect 64108 2297 64148 3424
rect 64203 3424 64204 3464
rect 64244 3424 64245 3464
rect 64203 3415 64245 3424
rect 64396 3464 64436 3473
rect 64204 3330 64244 3415
rect 64300 3212 64340 3221
rect 64203 2960 64245 2969
rect 64203 2920 64204 2960
rect 64244 2920 64245 2960
rect 64203 2911 64245 2920
rect 64204 2633 64244 2911
rect 64203 2624 64245 2633
rect 64203 2584 64204 2624
rect 64244 2584 64245 2624
rect 64203 2575 64245 2584
rect 64107 2288 64149 2297
rect 64107 2248 64108 2288
rect 64148 2248 64149 2288
rect 64107 2239 64149 2248
rect 64011 1700 64053 1709
rect 64011 1660 64012 1700
rect 64052 1660 64053 1700
rect 64011 1651 64053 1660
rect 64300 1616 64340 3172
rect 64396 3053 64436 3424
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 64780 3464 64820 3475
rect 64588 3330 64628 3415
rect 64780 3389 64820 3424
rect 65259 3464 65301 3473
rect 65259 3424 65260 3464
rect 65300 3424 65301 3464
rect 65259 3415 65301 3424
rect 65452 3464 65492 3499
rect 64779 3380 64821 3389
rect 64779 3340 64780 3380
rect 64820 3340 64821 3380
rect 64779 3331 64821 3340
rect 64684 3212 64724 3221
rect 64395 3044 64437 3053
rect 64395 3004 64396 3044
rect 64436 3004 64437 3044
rect 64395 2995 64437 3004
rect 64396 2213 64436 2995
rect 64395 2204 64437 2213
rect 64395 2164 64396 2204
rect 64436 2164 64437 2204
rect 64395 2155 64437 2164
rect 64204 1576 64340 1616
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 64204 1373 64244 1576
rect 64684 1373 64724 3172
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 65260 2120 65300 3415
rect 65452 3389 65492 3424
rect 65644 3464 65684 3499
rect 65644 3413 65684 3424
rect 65835 3464 65877 3473
rect 65835 3424 65836 3464
rect 65876 3424 65877 3464
rect 65835 3415 65877 3424
rect 66028 3464 66068 3499
rect 65451 3380 65493 3389
rect 65451 3340 65452 3380
rect 65492 3340 65493 3380
rect 65451 3331 65493 3340
rect 65452 3300 65492 3331
rect 65836 3330 65876 3415
rect 66028 3413 66068 3424
rect 66219 3464 66261 3473
rect 66219 3424 66220 3464
rect 66260 3424 66261 3464
rect 66219 3415 66261 3424
rect 66220 3330 66260 3415
rect 65355 3212 65397 3221
rect 65740 3212 65780 3221
rect 66124 3212 66164 3221
rect 65355 3172 65356 3212
rect 65396 3172 65397 3212
rect 65355 3163 65397 3172
rect 65644 3172 65740 3212
rect 65356 3078 65396 3163
rect 64876 2080 65300 2120
rect 64876 1952 64916 2080
rect 64876 1903 64916 1912
rect 65067 1952 65109 1961
rect 65067 1912 65068 1952
rect 65108 1912 65109 1952
rect 65067 1903 65109 1912
rect 65068 1818 65108 1903
rect 64972 1700 65012 1709
rect 65012 1660 65300 1700
rect 64972 1651 65012 1660
rect 64203 1364 64245 1373
rect 64203 1324 64204 1364
rect 64244 1324 64245 1364
rect 64203 1315 64245 1324
rect 64683 1364 64725 1373
rect 64683 1324 64684 1364
rect 64724 1324 64725 1364
rect 64683 1315 64725 1324
rect 63340 1240 63476 1280
rect 63723 1280 63765 1289
rect 63723 1240 63724 1280
rect 63764 1240 63765 1280
rect 63244 1121 63284 1206
rect 63243 1112 63285 1121
rect 63148 1069 63189 1109
rect 62860 953 62900 1061
rect 62763 944 62805 953
rect 62763 904 62764 944
rect 62804 904 62805 944
rect 62860 944 62906 953
rect 62860 904 62865 944
rect 62905 904 62906 944
rect 62763 895 62805 904
rect 62864 895 62906 904
rect 62572 820 62708 860
rect 62668 80 62708 820
rect 62764 810 62804 895
rect 63149 860 63189 1069
rect 63243 1072 63244 1112
rect 63284 1072 63285 1112
rect 63243 1063 63285 1072
rect 63243 944 63285 953
rect 63243 904 63244 944
rect 63284 904 63285 944
rect 63340 944 63380 1240
rect 63723 1231 63765 1240
rect 64875 1280 64917 1289
rect 64875 1240 64876 1280
rect 64916 1240 64917 1280
rect 64875 1231 64917 1240
rect 63531 1196 63573 1205
rect 63436 1156 63532 1196
rect 63572 1156 63573 1196
rect 63436 1112 63476 1156
rect 63531 1147 63573 1156
rect 63436 1063 63476 1072
rect 63627 1112 63669 1121
rect 63627 1072 63628 1112
rect 63668 1072 63669 1112
rect 63627 1063 63669 1072
rect 63724 1112 63764 1231
rect 64011 1196 64053 1205
rect 64011 1156 64012 1196
rect 64052 1156 64053 1196
rect 64011 1147 64053 1156
rect 64395 1196 64437 1205
rect 64395 1156 64396 1196
rect 64436 1156 64437 1196
rect 64395 1147 64437 1156
rect 63820 1125 63860 1140
rect 63724 1085 63820 1112
rect 63724 1072 63860 1085
rect 64012 1112 64052 1147
rect 63628 978 63668 1063
rect 63531 944 63573 953
rect 63340 904 63476 944
rect 63243 895 63285 904
rect 63148 820 63189 860
rect 63148 776 63188 820
rect 63052 736 63188 776
rect 62859 524 62901 533
rect 62859 484 62860 524
rect 62900 484 62901 524
rect 62859 475 62901 484
rect 62860 80 62900 475
rect 63052 80 63092 736
rect 63244 80 63284 895
rect 63436 80 63476 904
rect 63531 904 63532 944
rect 63572 904 63573 944
rect 63531 895 63573 904
rect 63532 810 63572 895
rect 63724 785 63764 1072
rect 64012 1061 64052 1072
rect 64204 1112 64244 1121
rect 64299 1112 64341 1121
rect 64244 1072 64300 1112
rect 64340 1072 64341 1112
rect 64204 1063 64244 1072
rect 64299 1063 64341 1072
rect 64396 1112 64436 1147
rect 64588 1121 64628 1206
rect 64779 1196 64821 1205
rect 64779 1156 64780 1196
rect 64820 1156 64821 1196
rect 64779 1147 64821 1156
rect 64396 1061 64436 1072
rect 64587 1112 64629 1121
rect 64587 1072 64588 1112
rect 64628 1072 64629 1112
rect 64587 1063 64629 1072
rect 64780 1112 64820 1147
rect 64780 1061 64820 1072
rect 64876 953 64916 1231
rect 65163 1196 65205 1205
rect 65163 1156 65164 1196
rect 65204 1156 65205 1196
rect 65163 1147 65205 1156
rect 64972 1112 65012 1123
rect 64972 1037 65012 1072
rect 65164 1112 65204 1147
rect 65164 1061 65204 1072
rect 64971 1028 65013 1037
rect 64971 988 64972 1028
rect 65012 988 65013 1028
rect 64971 979 65013 988
rect 65068 953 65108 1038
rect 63819 944 63861 953
rect 63819 904 63820 944
rect 63860 904 63861 944
rect 63819 895 63861 904
rect 63916 944 63956 953
rect 63723 776 63765 785
rect 63723 736 63724 776
rect 63764 736 63765 776
rect 63723 727 63765 736
rect 63627 524 63669 533
rect 63627 484 63628 524
rect 63668 484 63669 524
rect 63627 475 63669 484
rect 63628 80 63668 475
rect 63820 80 63860 895
rect 63916 533 63956 904
rect 64203 944 64245 953
rect 64203 904 64204 944
rect 64244 904 64245 944
rect 64203 895 64245 904
rect 64299 944 64341 953
rect 64684 944 64724 953
rect 64299 904 64300 944
rect 64340 904 64341 944
rect 64299 895 64341 904
rect 64396 904 64684 944
rect 63915 524 63957 533
rect 64204 524 64244 895
rect 64300 810 64340 895
rect 64396 860 64436 904
rect 64684 895 64724 904
rect 64875 944 64917 953
rect 64875 904 64876 944
rect 64916 904 64917 944
rect 64875 895 64917 904
rect 65067 944 65109 953
rect 65067 904 65068 944
rect 65108 904 65109 944
rect 65067 895 65109 904
rect 64393 820 64436 860
rect 64393 776 64433 820
rect 64683 776 64725 785
rect 64393 736 64436 776
rect 63915 484 63916 524
rect 63956 484 63957 524
rect 63915 475 63957 484
rect 64012 484 64244 524
rect 64012 80 64052 484
rect 64203 104 64245 113
rect 64203 80 64204 104
rect 20084 64 20104 80
rect 20024 0 20104 64
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 0 33544 80
rect 33656 0 33736 80
rect 33848 0 33928 80
rect 34040 0 34120 80
rect 34232 0 34312 80
rect 34424 0 34504 80
rect 34616 0 34696 80
rect 34808 0 34888 80
rect 35000 0 35080 80
rect 35192 0 35272 80
rect 35384 0 35464 80
rect 35576 0 35656 80
rect 35768 0 35848 80
rect 35960 0 36040 80
rect 36152 0 36232 80
rect 36344 0 36424 80
rect 36536 0 36616 80
rect 36728 0 36808 80
rect 36920 0 37000 80
rect 37112 0 37192 80
rect 37304 0 37384 80
rect 37496 0 37576 80
rect 37688 0 37768 80
rect 37880 0 37960 80
rect 38072 0 38152 80
rect 38264 0 38344 80
rect 38456 0 38536 80
rect 38648 0 38728 80
rect 38840 0 38920 80
rect 39032 0 39112 80
rect 39224 0 39304 80
rect 39416 0 39496 80
rect 39608 0 39688 80
rect 39800 0 39880 80
rect 39992 0 40072 80
rect 40184 0 40264 80
rect 40376 0 40456 80
rect 40568 0 40648 80
rect 40760 0 40840 80
rect 40952 0 41032 80
rect 41144 0 41224 80
rect 41336 0 41416 80
rect 41528 0 41608 80
rect 41720 0 41800 80
rect 41912 0 41992 80
rect 42104 0 42184 80
rect 42296 0 42376 80
rect 42488 0 42568 80
rect 42680 0 42760 80
rect 42872 0 42952 80
rect 43064 0 43144 80
rect 43256 0 43336 80
rect 43448 0 43528 80
rect 43640 0 43720 80
rect 43832 0 43912 80
rect 44024 0 44104 80
rect 44216 0 44296 80
rect 44408 0 44488 80
rect 44600 0 44680 80
rect 44792 0 44872 80
rect 44984 0 45064 80
rect 45176 0 45256 80
rect 45368 0 45448 80
rect 45560 0 45640 80
rect 45752 0 45832 80
rect 45944 0 46024 80
rect 46136 0 46216 80
rect 46328 0 46408 80
rect 46520 0 46600 80
rect 46712 0 46792 80
rect 46904 0 46984 80
rect 47096 0 47176 80
rect 47288 0 47368 80
rect 47480 0 47560 80
rect 47672 0 47752 80
rect 47864 0 47944 80
rect 48056 0 48136 80
rect 48248 0 48328 80
rect 48440 0 48520 80
rect 48632 0 48712 80
rect 48824 0 48904 80
rect 49016 0 49096 80
rect 49208 0 49288 80
rect 49400 0 49480 80
rect 49592 0 49672 80
rect 49784 0 49864 80
rect 49976 0 50056 80
rect 50168 0 50248 80
rect 50360 0 50440 80
rect 50552 0 50632 80
rect 50744 0 50824 80
rect 50936 0 51016 80
rect 51128 0 51208 80
rect 51320 0 51400 80
rect 51512 0 51592 80
rect 51704 0 51784 80
rect 51896 0 51976 80
rect 52088 0 52168 80
rect 52280 0 52360 80
rect 52472 0 52552 80
rect 52664 0 52744 80
rect 52856 0 52936 80
rect 53048 0 53128 80
rect 53240 0 53320 80
rect 53432 0 53512 80
rect 53624 0 53704 80
rect 53816 0 53896 80
rect 54008 0 54088 80
rect 54200 0 54280 80
rect 54392 0 54472 80
rect 54584 0 54664 80
rect 54776 0 54856 80
rect 54968 0 55048 80
rect 55160 0 55240 80
rect 55352 0 55432 80
rect 55544 0 55624 80
rect 55736 0 55816 80
rect 55928 0 56008 80
rect 56120 0 56200 80
rect 56312 0 56392 80
rect 56504 0 56584 80
rect 56696 0 56776 80
rect 56888 0 56968 80
rect 57080 0 57160 80
rect 57272 0 57352 80
rect 57464 0 57544 80
rect 57656 0 57736 80
rect 57848 0 57928 80
rect 58040 0 58120 80
rect 58232 0 58312 80
rect 58424 0 58504 80
rect 58616 0 58696 80
rect 58808 0 58888 80
rect 59000 0 59080 80
rect 59192 0 59272 80
rect 59384 0 59464 80
rect 59576 0 59656 80
rect 59768 0 59848 80
rect 59960 0 60040 80
rect 60152 0 60232 80
rect 60344 0 60424 80
rect 60536 0 60616 80
rect 60728 0 60808 80
rect 60920 0 61000 80
rect 61112 0 61192 80
rect 61304 0 61384 80
rect 61496 0 61576 80
rect 61688 0 61768 80
rect 61880 0 61960 80
rect 62072 0 62152 80
rect 62264 0 62344 80
rect 62456 0 62536 80
rect 62648 0 62728 80
rect 62840 0 62920 80
rect 63032 0 63112 80
rect 63224 0 63304 80
rect 63416 0 63496 80
rect 63608 0 63688 80
rect 63800 0 63880 80
rect 63992 0 64072 80
rect 64184 64 64204 80
rect 64244 80 64245 104
rect 64396 80 64436 736
rect 64683 736 64684 776
rect 64724 736 64725 776
rect 64683 727 64725 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 64587 524 64629 533
rect 64587 484 64588 524
rect 64628 484 64629 524
rect 64684 524 64724 727
rect 65260 608 65300 1660
rect 65548 1205 65588 1207
rect 65547 1196 65589 1205
rect 65547 1156 65548 1196
rect 65588 1156 65589 1196
rect 65547 1147 65589 1156
rect 65356 1112 65396 1121
rect 65451 1112 65493 1121
rect 65451 1109 65452 1112
rect 65396 1072 65452 1109
rect 65492 1072 65493 1112
rect 65356 1069 65493 1072
rect 65356 1063 65396 1069
rect 65451 1063 65493 1069
rect 65548 1112 65588 1147
rect 65548 1063 65588 1072
rect 65355 944 65397 953
rect 65355 904 65356 944
rect 65396 904 65397 944
rect 65355 895 65397 904
rect 65452 944 65492 953
rect 64972 568 65300 608
rect 64684 484 64820 524
rect 64587 475 64629 484
rect 64588 80 64628 475
rect 64780 80 64820 484
rect 64972 80 65012 568
rect 65163 440 65205 449
rect 65163 400 65164 440
rect 65204 400 65205 440
rect 65163 391 65205 400
rect 65164 80 65204 391
rect 65356 80 65396 895
rect 65452 449 65492 904
rect 65547 944 65589 953
rect 65547 904 65548 944
rect 65588 904 65589 944
rect 65644 944 65684 3172
rect 65740 3163 65780 3172
rect 66028 3172 66124 3212
rect 65740 1121 65780 1206
rect 65931 1196 65973 1205
rect 65931 1156 65932 1196
rect 65972 1156 65973 1196
rect 65931 1147 65973 1156
rect 65739 1112 65781 1121
rect 65739 1072 65740 1112
rect 65780 1072 65781 1112
rect 65739 1063 65781 1072
rect 65932 1112 65972 1147
rect 65932 1061 65972 1072
rect 65835 944 65877 953
rect 65644 904 65780 944
rect 65547 895 65589 904
rect 65451 440 65493 449
rect 65451 400 65452 440
rect 65492 400 65493 440
rect 65451 391 65493 400
rect 65548 80 65588 895
rect 65740 80 65780 904
rect 65835 904 65836 944
rect 65876 904 65877 944
rect 65835 895 65877 904
rect 65836 810 65876 895
rect 66028 860 66068 3172
rect 66124 3163 66164 3172
rect 66412 2708 66452 3835
rect 66604 3834 66644 3919
rect 66892 3632 66932 4012
rect 66988 4002 67028 4087
rect 67180 3977 67220 4684
rect 69100 4229 69140 4759
rect 73324 4724 73364 4733
rect 68523 4220 68565 4229
rect 68523 4180 68524 4220
rect 68564 4180 68565 4220
rect 68523 4171 68565 4180
rect 69099 4220 69141 4229
rect 69099 4180 69100 4220
rect 69140 4180 69141 4220
rect 69099 4171 69141 4180
rect 68524 4136 68564 4171
rect 68524 4085 68564 4096
rect 68908 4136 68948 4145
rect 68908 3977 68948 4096
rect 69100 4136 69140 4171
rect 73324 4145 73364 4684
rect 73612 4313 73652 4936
rect 73803 4976 73845 4985
rect 73803 4936 73804 4976
rect 73844 4936 73845 4976
rect 73803 4927 73845 4936
rect 74092 4976 74132 4985
rect 73804 4842 73844 4927
rect 74092 4892 74132 4936
rect 74283 4976 74325 4985
rect 74283 4936 74284 4976
rect 74324 4936 74325 4976
rect 74283 4927 74325 4936
rect 74476 4976 74516 4985
rect 82155 4976 82197 4985
rect 73996 4852 74132 4892
rect 73611 4304 73653 4313
rect 73611 4264 73612 4304
rect 73652 4264 73653 4304
rect 73996 4304 74036 4852
rect 74092 4724 74132 4733
rect 74092 4481 74132 4684
rect 74187 4640 74229 4649
rect 74187 4600 74188 4640
rect 74228 4600 74229 4640
rect 74187 4591 74229 4600
rect 74091 4472 74133 4481
rect 74091 4432 74092 4472
rect 74132 4432 74133 4472
rect 74091 4423 74133 4432
rect 74091 4304 74133 4313
rect 73996 4264 74092 4304
rect 74132 4264 74133 4304
rect 73611 4255 73653 4264
rect 74091 4255 74133 4264
rect 69100 4086 69140 4096
rect 73323 4136 73365 4145
rect 73323 4096 73324 4136
rect 73364 4096 73365 4136
rect 73323 4087 73365 4096
rect 74092 4136 74132 4255
rect 74188 4145 74228 4591
rect 74284 4229 74324 4927
rect 74380 4892 74420 4903
rect 74380 4817 74420 4852
rect 74379 4808 74421 4817
rect 74379 4768 74380 4808
rect 74420 4768 74421 4808
rect 74379 4759 74421 4768
rect 74476 4313 74516 4936
rect 82060 4936 82156 4976
rect 82196 4936 82197 4976
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 80523 4472 80565 4481
rect 80523 4432 80524 4472
rect 80564 4432 80565 4472
rect 80523 4423 80565 4432
rect 74475 4304 74517 4313
rect 74475 4264 74476 4304
rect 74516 4264 74517 4304
rect 74475 4255 74517 4264
rect 74667 4304 74709 4313
rect 74667 4264 74668 4304
rect 74708 4264 74709 4304
rect 74667 4255 74709 4264
rect 74283 4220 74325 4229
rect 74283 4180 74284 4220
rect 74324 4180 74325 4220
rect 74283 4171 74325 4180
rect 74092 4087 74132 4096
rect 74187 4136 74229 4145
rect 74187 4096 74188 4136
rect 74228 4096 74229 4136
rect 74187 4087 74229 4096
rect 74284 4136 74324 4171
rect 74284 4086 74324 4096
rect 74379 4136 74421 4145
rect 74379 4096 74380 4136
rect 74420 4096 74421 4136
rect 74379 4087 74421 4096
rect 69004 4052 69044 4061
rect 67179 3968 67221 3977
rect 67179 3928 67180 3968
rect 67220 3928 67221 3968
rect 67179 3919 67221 3928
rect 68427 3968 68469 3977
rect 68427 3928 68428 3968
rect 68468 3928 68469 3968
rect 68427 3919 68469 3928
rect 68716 3968 68756 3977
rect 68428 3834 68468 3919
rect 67371 3632 67413 3641
rect 66892 3592 67124 3632
rect 66795 3464 66837 3473
rect 66795 3424 66796 3464
rect 66836 3424 66837 3464
rect 66795 3415 66837 3424
rect 66988 3464 67028 3473
rect 66124 2668 66452 2708
rect 66124 1121 66164 2668
rect 66796 2549 66836 3415
rect 66988 3305 67028 3424
rect 66987 3296 67029 3305
rect 66987 3256 66988 3296
rect 67028 3256 67029 3296
rect 66987 3247 67029 3256
rect 66892 3212 66932 3221
rect 66795 2540 66837 2549
rect 66412 2500 66796 2540
rect 66836 2500 66837 2540
rect 66892 2540 66932 3172
rect 66892 2500 67028 2540
rect 66412 1952 66452 2500
rect 66795 2491 66837 2500
rect 66603 2372 66645 2381
rect 66603 2332 66604 2372
rect 66644 2332 66645 2372
rect 66603 2323 66645 2332
rect 66412 1903 66452 1912
rect 66604 1952 66644 2323
rect 66604 1903 66644 1912
rect 66508 1700 66548 1709
rect 66412 1660 66508 1700
rect 66315 1196 66357 1205
rect 66315 1156 66316 1196
rect 66356 1156 66357 1196
rect 66315 1147 66357 1156
rect 66123 1112 66165 1121
rect 66123 1072 66124 1112
rect 66164 1072 66165 1112
rect 66123 1063 66165 1072
rect 66316 1112 66356 1147
rect 66316 1061 66356 1072
rect 66220 944 66260 953
rect 66028 820 66164 860
rect 65931 524 65973 533
rect 65931 484 65932 524
rect 65972 484 65973 524
rect 65931 475 65973 484
rect 65932 80 65972 475
rect 66124 80 66164 820
rect 66220 533 66260 904
rect 66412 860 66452 1660
rect 66508 1651 66548 1660
rect 66892 1373 66932 1458
rect 66891 1364 66933 1373
rect 66891 1324 66892 1364
rect 66932 1324 66933 1364
rect 66891 1315 66933 1324
rect 66507 1280 66549 1289
rect 66507 1240 66508 1280
rect 66548 1240 66549 1280
rect 66507 1231 66549 1240
rect 66508 1112 66548 1231
rect 66700 1205 66740 1207
rect 66604 1196 66644 1205
rect 66508 1063 66548 1072
rect 66597 1156 66604 1196
rect 66597 1147 66644 1156
rect 66699 1196 66741 1205
rect 66699 1156 66700 1196
rect 66740 1156 66741 1196
rect 66699 1147 66741 1156
rect 66796 1156 66925 1196
rect 66597 944 66637 1147
rect 66700 1112 66740 1147
rect 66700 1063 66740 1072
rect 66699 944 66741 953
rect 66597 904 66644 944
rect 66412 820 66548 860
rect 66219 524 66261 533
rect 66219 484 66220 524
rect 66260 484 66261 524
rect 66219 475 66261 484
rect 66315 440 66357 449
rect 66315 400 66316 440
rect 66356 400 66357 440
rect 66315 391 66357 400
rect 66316 80 66356 391
rect 66508 80 66548 820
rect 66604 449 66644 904
rect 66699 904 66700 944
rect 66740 904 66741 944
rect 66699 895 66741 904
rect 66603 440 66645 449
rect 66603 400 66604 440
rect 66644 400 66645 440
rect 66603 391 66645 400
rect 66700 80 66740 895
rect 66796 617 66836 1156
rect 66885 1125 66925 1156
rect 66885 1076 66925 1085
rect 66988 1028 67028 2500
rect 67084 1205 67124 3592
rect 67371 3592 67372 3632
rect 67412 3592 67413 3632
rect 67371 3583 67413 3592
rect 67179 3464 67221 3473
rect 67179 3424 67180 3464
rect 67220 3424 67221 3464
rect 67179 3415 67221 3424
rect 67372 3464 67412 3583
rect 68619 3548 68661 3557
rect 68619 3508 68620 3548
rect 68660 3508 68661 3548
rect 68619 3499 68661 3508
rect 67372 3415 67412 3424
rect 68620 3464 68660 3499
rect 68716 3464 68756 3928
rect 68907 3968 68949 3977
rect 68907 3928 68908 3968
rect 68948 3928 68949 3968
rect 68907 3919 68949 3928
rect 69004 3632 69044 4012
rect 74380 4002 74420 4087
rect 74092 3968 74132 3977
rect 73996 3928 74092 3968
rect 74668 3968 74708 4255
rect 74763 4220 74805 4229
rect 74763 4180 74764 4220
rect 74804 4180 74805 4220
rect 74763 4171 74805 4180
rect 74764 4136 74804 4171
rect 74764 4085 74804 4096
rect 74859 4136 74901 4145
rect 74859 4096 74860 4136
rect 74900 4096 74901 4136
rect 74859 4087 74901 4096
rect 80331 4136 80373 4145
rect 80331 4096 80332 4136
rect 80372 4096 80373 4136
rect 80331 4087 80373 4096
rect 80524 4136 80564 4423
rect 82060 4397 82100 4936
rect 82155 4927 82197 4936
rect 82348 4976 82388 4987
rect 82828 4985 82868 9920
rect 93772 9260 93812 9920
rect 93676 9220 93812 9260
rect 93676 4985 93716 9220
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 82348 4901 82388 4936
rect 82827 4976 82869 4985
rect 82827 4936 82828 4976
rect 82868 4936 82869 4976
rect 82827 4927 82869 4936
rect 93675 4976 93717 4985
rect 93675 4936 93676 4976
rect 93716 4936 93717 4976
rect 93675 4927 93717 4936
rect 82347 4892 82389 4901
rect 82347 4852 82348 4892
rect 82388 4852 82389 4892
rect 82347 4843 82389 4852
rect 91755 4808 91797 4817
rect 91755 4768 91756 4808
rect 91796 4768 91797 4808
rect 91755 4759 91797 4768
rect 82156 4724 82196 4733
rect 82059 4388 82101 4397
rect 82059 4348 82060 4388
rect 82100 4348 82101 4388
rect 82059 4339 82101 4348
rect 82156 4229 82196 4684
rect 86571 4640 86613 4649
rect 86571 4600 86572 4640
rect 86612 4600 86613 4640
rect 86571 4591 86613 4600
rect 82155 4220 82197 4229
rect 82155 4180 82156 4220
rect 82196 4180 82197 4220
rect 82155 4171 82197 4180
rect 86572 4145 86612 4591
rect 86667 4220 86709 4229
rect 86667 4180 86668 4220
rect 86708 4180 86709 4220
rect 86667 4171 86709 4180
rect 80811 4136 80853 4145
rect 80564 4096 80756 4136
rect 80524 4087 80564 4096
rect 74860 4002 74900 4087
rect 75052 4052 75092 4061
rect 74764 3968 74804 3977
rect 74668 3928 74764 3968
rect 72075 3800 72117 3809
rect 72075 3760 72076 3800
rect 72116 3760 72117 3800
rect 72075 3751 72117 3760
rect 70155 3716 70197 3725
rect 70155 3676 70156 3716
rect 70196 3676 70197 3716
rect 70155 3667 70197 3676
rect 68908 3592 69044 3632
rect 68811 3464 68853 3473
rect 68716 3424 68812 3464
rect 68852 3424 68853 3464
rect 67180 3330 67220 3415
rect 68620 3413 68660 3424
rect 68811 3415 68853 3424
rect 68812 3330 68852 3415
rect 67371 3296 67413 3305
rect 67371 3256 67372 3296
rect 67412 3256 67413 3296
rect 67371 3247 67413 3256
rect 67276 3212 67316 3221
rect 67180 3172 67276 3212
rect 67083 1196 67125 1205
rect 67083 1156 67084 1196
rect 67124 1156 67125 1196
rect 67083 1147 67125 1156
rect 67084 1112 67124 1147
rect 67084 1063 67124 1072
rect 66902 988 67028 1028
rect 66902 944 66942 988
rect 66892 904 66942 944
rect 67083 944 67125 953
rect 67083 904 67084 944
rect 67124 904 67125 944
rect 67180 944 67220 3172
rect 67276 3163 67316 3172
rect 67372 3053 67412 3247
rect 68716 3212 68756 3221
rect 68332 3172 68716 3212
rect 67371 3044 67413 3053
rect 67371 3004 67372 3044
rect 67412 3004 67413 3044
rect 67371 2995 67413 3004
rect 67371 2624 67413 2633
rect 67371 2584 67372 2624
rect 67412 2584 67413 2624
rect 67371 2575 67413 2584
rect 67564 2624 67604 2633
rect 67372 2490 67412 2575
rect 67468 2540 67508 2549
rect 67468 1448 67508 2500
rect 67564 2465 67604 2584
rect 67563 2456 67605 2465
rect 67563 2416 67564 2456
rect 67604 2416 67605 2456
rect 67563 2407 67605 2416
rect 67564 1952 67604 2407
rect 67660 1952 67700 1961
rect 67564 1912 67660 1952
rect 67660 1903 67700 1912
rect 67851 1952 67893 1961
rect 67851 1912 67852 1952
rect 67892 1912 67893 1952
rect 67851 1903 67893 1912
rect 67852 1818 67892 1903
rect 67756 1700 67796 1709
rect 67796 1660 67988 1700
rect 67756 1651 67796 1660
rect 67468 1408 67604 1448
rect 67275 1196 67317 1205
rect 67275 1156 67276 1196
rect 67316 1156 67317 1196
rect 67275 1147 67317 1156
rect 67276 1112 67316 1147
rect 67276 1061 67316 1072
rect 67467 1112 67509 1121
rect 67467 1072 67468 1112
rect 67508 1072 67509 1112
rect 67467 1063 67509 1072
rect 67468 978 67508 1063
rect 67371 944 67413 953
rect 67180 904 67316 944
rect 66795 608 66837 617
rect 66795 568 66796 608
rect 66836 568 66837 608
rect 66795 559 66837 568
rect 66796 449 66836 559
rect 66795 440 66837 449
rect 66795 400 66796 440
rect 66836 400 66837 440
rect 66795 391 66837 400
rect 66892 80 66932 904
rect 67083 895 67125 904
rect 67084 80 67124 895
rect 67276 80 67316 904
rect 67371 904 67372 944
rect 67412 904 67413 944
rect 67371 895 67413 904
rect 67372 810 67412 895
rect 67564 776 67604 1408
rect 67852 1121 67892 1206
rect 67660 1112 67700 1121
rect 67660 860 67700 1072
rect 67851 1112 67893 1121
rect 67851 1072 67852 1112
rect 67892 1072 67893 1112
rect 67851 1063 67893 1072
rect 67756 1028 67796 1037
rect 67756 944 67796 988
rect 67756 904 67892 944
rect 67660 820 67796 860
rect 67564 736 67700 776
rect 67467 692 67509 701
rect 67467 652 67468 692
rect 67508 652 67509 692
rect 67467 643 67509 652
rect 67468 80 67508 643
rect 67660 80 67700 736
rect 67756 617 67796 820
rect 67852 701 67892 904
rect 67948 860 67988 1660
rect 68043 1196 68085 1205
rect 68043 1156 68044 1196
rect 68084 1156 68085 1196
rect 68043 1147 68085 1156
rect 68044 1112 68084 1147
rect 68236 1121 68276 1206
rect 68044 1061 68084 1072
rect 68235 1112 68277 1121
rect 68235 1072 68236 1112
rect 68276 1072 68277 1112
rect 68235 1063 68277 1072
rect 68140 944 68180 953
rect 67948 820 68084 860
rect 67851 692 67893 701
rect 67851 652 67852 692
rect 67892 652 67893 692
rect 67851 643 67893 652
rect 67755 608 67797 617
rect 67755 568 67756 608
rect 67796 568 67797 608
rect 67755 559 67797 568
rect 67756 197 67796 559
rect 67851 524 67893 533
rect 67851 484 67852 524
rect 67892 484 67893 524
rect 67851 475 67893 484
rect 67755 188 67797 197
rect 67755 148 67756 188
rect 67796 148 67797 188
rect 67755 139 67797 148
rect 67852 80 67892 475
rect 68044 80 68084 820
rect 68140 533 68180 904
rect 68235 944 68277 953
rect 68235 904 68236 944
rect 68276 904 68277 944
rect 68332 944 68372 3172
rect 68716 3163 68756 3172
rect 68715 1616 68757 1625
rect 68715 1576 68716 1616
rect 68756 1576 68757 1616
rect 68715 1567 68757 1576
rect 68428 1121 68468 1206
rect 68620 1121 68660 1206
rect 68427 1112 68469 1121
rect 68427 1072 68428 1112
rect 68468 1072 68469 1112
rect 68427 1063 68469 1072
rect 68619 1112 68661 1121
rect 68619 1072 68620 1112
rect 68660 1072 68661 1112
rect 68619 1063 68661 1072
rect 68523 944 68565 953
rect 68332 904 68468 944
rect 68235 895 68277 904
rect 68139 524 68181 533
rect 68139 484 68140 524
rect 68180 484 68181 524
rect 68139 475 68181 484
rect 68236 80 68276 895
rect 68428 80 68468 904
rect 68523 904 68524 944
rect 68564 904 68565 944
rect 68716 944 68756 1567
rect 68812 1121 68852 1206
rect 68811 1112 68853 1121
rect 68811 1072 68812 1112
rect 68852 1072 68853 1112
rect 68908 1112 68948 3592
rect 69771 3548 69813 3557
rect 69771 3508 69772 3548
rect 69812 3508 69813 3548
rect 69771 3499 69813 3508
rect 69004 3464 69044 3473
rect 69004 2717 69044 3424
rect 69195 3464 69237 3473
rect 69195 3424 69196 3464
rect 69236 3424 69237 3464
rect 69195 3415 69237 3424
rect 69388 3464 69428 3473
rect 69196 3330 69236 3415
rect 69100 3212 69140 3221
rect 69003 2708 69045 2717
rect 69003 2668 69004 2708
rect 69044 2668 69045 2708
rect 69003 2659 69045 2668
rect 69004 2213 69044 2659
rect 69003 2204 69045 2213
rect 69003 2164 69004 2204
rect 69044 2164 69045 2204
rect 69003 2155 69045 2164
rect 69100 1625 69140 3172
rect 69388 3137 69428 3424
rect 69579 3464 69621 3473
rect 69579 3424 69580 3464
rect 69620 3424 69621 3464
rect 69579 3415 69621 3424
rect 69772 3464 69812 3499
rect 69580 3330 69620 3415
rect 69772 3413 69812 3424
rect 69963 3464 70005 3473
rect 69963 3424 69964 3464
rect 70004 3424 70005 3464
rect 69963 3415 70005 3424
rect 70156 3464 70196 3667
rect 71307 3548 71349 3557
rect 71307 3508 71308 3548
rect 71348 3508 71349 3548
rect 71307 3499 71349 3508
rect 71691 3548 71733 3557
rect 71691 3508 71692 3548
rect 71732 3508 71733 3548
rect 71691 3499 71733 3508
rect 70156 3415 70196 3424
rect 70347 3464 70389 3473
rect 70347 3424 70348 3464
rect 70388 3424 70389 3464
rect 70347 3415 70389 3424
rect 70540 3464 70580 3473
rect 69964 3330 70004 3415
rect 70348 3330 70388 3415
rect 70540 3305 70580 3424
rect 70731 3464 70773 3473
rect 70731 3424 70732 3464
rect 70772 3424 70773 3464
rect 70731 3415 70773 3424
rect 70924 3464 70964 3473
rect 70732 3330 70772 3415
rect 70539 3296 70581 3305
rect 70539 3256 70540 3296
rect 70580 3256 70581 3296
rect 70539 3247 70581 3256
rect 69484 3212 69524 3221
rect 69868 3212 69908 3221
rect 70252 3212 70292 3221
rect 69387 3128 69429 3137
rect 69387 3088 69388 3128
rect 69428 3088 69429 3128
rect 69387 3079 69429 3088
rect 69388 2885 69428 3079
rect 69387 2876 69429 2885
rect 69387 2836 69388 2876
rect 69428 2836 69429 2876
rect 69387 2827 69429 2836
rect 69484 2540 69524 3172
rect 69196 2500 69524 2540
rect 69580 3172 69868 3212
rect 69099 1616 69141 1625
rect 69099 1576 69100 1616
rect 69140 1576 69141 1616
rect 69099 1567 69141 1576
rect 69196 1280 69236 2500
rect 69387 1448 69429 1457
rect 69387 1408 69388 1448
rect 69428 1408 69429 1448
rect 69387 1399 69429 1408
rect 69100 1240 69236 1280
rect 69003 1112 69045 1121
rect 68908 1072 69004 1112
rect 69044 1072 69045 1112
rect 68811 1063 68853 1072
rect 69003 1063 69045 1072
rect 69004 978 69044 1063
rect 68908 944 68948 953
rect 68716 904 68852 944
rect 68523 895 68565 904
rect 68524 810 68564 895
rect 68619 692 68661 701
rect 68619 652 68620 692
rect 68660 652 68661 692
rect 68619 643 68661 652
rect 68620 80 68660 643
rect 68812 80 68852 904
rect 68908 701 68948 904
rect 69100 860 69140 1240
rect 69195 1112 69237 1121
rect 69195 1072 69196 1112
rect 69236 1072 69237 1112
rect 69195 1063 69237 1072
rect 69388 1112 69428 1399
rect 69580 1364 69620 3172
rect 69868 3163 69908 3172
rect 70060 3172 70252 3212
rect 70060 2540 70100 3172
rect 70252 3163 70292 3172
rect 70636 3212 70676 3221
rect 69388 1063 69428 1072
rect 69484 1324 69620 1364
rect 69868 2500 70100 2540
rect 69196 978 69236 1063
rect 69292 944 69332 953
rect 69100 820 69236 860
rect 68907 692 68949 701
rect 68907 652 68908 692
rect 68948 652 68949 692
rect 68907 643 68949 652
rect 69003 524 69045 533
rect 69003 484 69004 524
rect 69044 484 69045 524
rect 69003 475 69045 484
rect 69004 80 69044 475
rect 69196 80 69236 820
rect 69292 533 69332 904
rect 69387 944 69429 953
rect 69387 904 69388 944
rect 69428 904 69429 944
rect 69484 944 69524 1324
rect 69771 1196 69813 1205
rect 69771 1156 69772 1196
rect 69812 1156 69813 1196
rect 69771 1147 69813 1156
rect 69590 1112 69630 1118
rect 69675 1112 69717 1121
rect 69590 1109 69676 1112
rect 69630 1072 69676 1109
rect 69716 1072 69717 1112
rect 69590 1060 69630 1069
rect 69675 1063 69717 1072
rect 69772 1112 69812 1147
rect 69772 1061 69812 1072
rect 69675 944 69717 953
rect 69484 904 69620 944
rect 69387 895 69429 904
rect 69291 524 69333 533
rect 69291 484 69292 524
rect 69332 484 69333 524
rect 69291 475 69333 484
rect 69388 80 69428 895
rect 69580 80 69620 904
rect 69675 904 69676 944
rect 69716 904 69717 944
rect 69675 895 69717 904
rect 69676 810 69716 895
rect 69868 860 69908 2500
rect 70636 1289 70676 3172
rect 70924 3053 70964 3424
rect 71115 3464 71157 3473
rect 71115 3424 71116 3464
rect 71156 3424 71157 3464
rect 71115 3415 71157 3424
rect 71308 3464 71348 3499
rect 71116 3330 71156 3415
rect 71308 3413 71348 3424
rect 71499 3464 71541 3473
rect 71499 3424 71500 3464
rect 71540 3424 71541 3464
rect 71499 3415 71541 3424
rect 71692 3464 71732 3499
rect 71500 3330 71540 3415
rect 71692 3389 71732 3424
rect 71883 3464 71925 3473
rect 71883 3424 71884 3464
rect 71924 3424 71925 3464
rect 71883 3415 71925 3424
rect 72076 3464 72116 3751
rect 73323 3632 73365 3641
rect 73323 3592 73324 3632
rect 73364 3592 73365 3632
rect 73323 3583 73365 3592
rect 71691 3380 71733 3389
rect 71691 3340 71692 3380
rect 71732 3340 71733 3380
rect 71691 3331 71733 3340
rect 71692 3300 71732 3331
rect 71884 3330 71924 3415
rect 71020 3212 71060 3221
rect 71404 3212 71444 3221
rect 70923 3044 70965 3053
rect 70923 3004 70924 3044
rect 70964 3004 70965 3044
rect 70923 2995 70965 3004
rect 70924 2801 70964 2995
rect 70923 2792 70965 2801
rect 70923 2752 70924 2792
rect 70964 2752 70965 2792
rect 70923 2743 70965 2752
rect 71020 2540 71060 3172
rect 70828 2500 71060 2540
rect 71212 3172 71404 3212
rect 70731 1532 70773 1541
rect 70731 1492 70732 1532
rect 70772 1492 70773 1532
rect 70731 1483 70773 1492
rect 70732 1364 70772 1483
rect 70732 1315 70772 1324
rect 70251 1280 70293 1289
rect 70251 1240 70252 1280
rect 70292 1240 70293 1280
rect 70251 1231 70293 1240
rect 70635 1280 70677 1289
rect 70635 1240 70636 1280
rect 70676 1240 70677 1280
rect 70635 1231 70677 1240
rect 70155 1196 70197 1205
rect 70155 1156 70156 1196
rect 70196 1156 70197 1196
rect 70155 1147 70197 1156
rect 69963 1112 70005 1121
rect 69963 1072 69964 1112
rect 70004 1072 70005 1112
rect 69963 1063 70005 1072
rect 70156 1112 70196 1147
rect 69964 978 70004 1063
rect 70156 1061 70196 1072
rect 70060 944 70100 953
rect 69868 820 70004 860
rect 69771 524 69813 533
rect 69771 484 69772 524
rect 69812 484 69813 524
rect 69771 475 69813 484
rect 69772 80 69812 475
rect 69964 80 70004 820
rect 70060 533 70100 904
rect 70155 944 70197 953
rect 70155 904 70156 944
rect 70196 904 70197 944
rect 70155 895 70197 904
rect 70059 524 70101 533
rect 70059 484 70060 524
rect 70100 484 70101 524
rect 70059 475 70101 484
rect 70156 80 70196 895
rect 70252 860 70292 1231
rect 70520 1196 70562 1205
rect 70520 1156 70521 1196
rect 70561 1156 70562 1196
rect 70520 1147 70562 1156
rect 70347 1112 70389 1121
rect 70347 1072 70348 1112
rect 70388 1072 70389 1112
rect 70347 1063 70389 1072
rect 70521 1117 70561 1147
rect 70348 978 70388 1063
rect 70521 1061 70561 1077
rect 70635 1112 70677 1121
rect 70635 1072 70636 1112
rect 70676 1109 70677 1112
rect 70732 1112 70772 1121
rect 70676 1072 70732 1109
rect 70635 1069 70772 1072
rect 70635 1063 70677 1069
rect 70732 1063 70772 1069
rect 70443 944 70485 953
rect 70443 904 70444 944
rect 70484 904 70485 944
rect 70443 895 70485 904
rect 70252 820 70388 860
rect 70348 80 70388 820
rect 70444 810 70484 895
rect 70828 860 70868 2500
rect 70923 1532 70965 1541
rect 70923 1492 70924 1532
rect 70964 1492 70965 1532
rect 70923 1483 70965 1492
rect 70732 820 70868 860
rect 70924 1112 70964 1483
rect 71212 1364 71252 3172
rect 71404 3163 71444 3172
rect 71788 3212 71828 3221
rect 71788 1373 71828 3172
rect 72076 2969 72116 3424
rect 72267 3464 72309 3473
rect 72267 3424 72268 3464
rect 72308 3424 72309 3464
rect 72267 3415 72309 3424
rect 72460 3464 72500 3475
rect 72268 3330 72308 3415
rect 72460 3389 72500 3424
rect 72651 3464 72693 3473
rect 72651 3424 72652 3464
rect 72692 3424 72693 3464
rect 72651 3415 72693 3424
rect 72843 3464 72885 3473
rect 72843 3424 72844 3464
rect 72884 3424 72885 3464
rect 72843 3415 72885 3424
rect 73036 3464 73076 3475
rect 72459 3380 72501 3389
rect 72459 3340 72460 3380
rect 72500 3340 72501 3380
rect 72459 3331 72501 3340
rect 72172 3212 72212 3221
rect 72075 2960 72117 2969
rect 72075 2920 72076 2960
rect 72116 2920 72117 2960
rect 72075 2911 72117 2920
rect 70539 188 70581 197
rect 70539 148 70540 188
rect 70580 148 70581 188
rect 70539 139 70581 148
rect 70540 80 70580 139
rect 70732 80 70772 820
rect 70924 692 70964 1072
rect 71020 1324 71252 1364
rect 71787 1364 71829 1373
rect 71787 1324 71788 1364
rect 71828 1324 71829 1364
rect 71020 944 71060 1324
rect 71787 1315 71829 1324
rect 71116 1121 71156 1206
rect 71115 1112 71157 1121
rect 71115 1072 71116 1112
rect 71156 1072 71157 1112
rect 71115 1063 71157 1072
rect 71308 1112 71348 1123
rect 71884 1121 71924 1206
rect 72075 1196 72117 1205
rect 72075 1156 72076 1196
rect 72116 1156 72117 1196
rect 72075 1147 72117 1156
rect 71212 953 71252 1038
rect 71308 1037 71348 1072
rect 71499 1112 71541 1121
rect 71499 1072 71500 1112
rect 71540 1072 71541 1112
rect 71499 1063 71541 1072
rect 71692 1112 71732 1121
rect 71883 1112 71925 1121
rect 71732 1072 71828 1112
rect 71692 1063 71732 1072
rect 71307 1028 71349 1037
rect 71307 988 71308 1028
rect 71348 988 71349 1028
rect 71307 979 71349 988
rect 71500 978 71540 1063
rect 71211 944 71253 953
rect 71020 904 71157 944
rect 71117 860 71157 904
rect 71211 904 71212 944
rect 71252 904 71253 944
rect 71211 895 71253 904
rect 71596 944 71636 953
rect 70828 652 70964 692
rect 71116 820 71157 860
rect 71499 860 71541 869
rect 71499 820 71500 860
rect 71540 820 71541 860
rect 70828 281 70868 652
rect 70923 524 70965 533
rect 70923 484 70924 524
rect 70964 484 70965 524
rect 70923 475 70965 484
rect 70827 272 70869 281
rect 70827 232 70828 272
rect 70868 232 70869 272
rect 70827 223 70869 232
rect 70924 80 70964 475
rect 71116 80 71156 820
rect 71499 811 71541 820
rect 71307 524 71349 533
rect 71307 484 71308 524
rect 71348 484 71349 524
rect 71307 475 71349 484
rect 71308 80 71348 475
rect 71500 80 71540 811
rect 71596 533 71636 904
rect 71691 944 71733 953
rect 71691 904 71692 944
rect 71732 904 71733 944
rect 71691 895 71733 904
rect 71595 524 71637 533
rect 71595 484 71596 524
rect 71636 484 71637 524
rect 71595 475 71637 484
rect 71692 80 71732 895
rect 71788 617 71828 1072
rect 71883 1072 71884 1112
rect 71924 1072 71925 1112
rect 71883 1063 71925 1072
rect 72076 1112 72116 1147
rect 72076 1061 72116 1072
rect 71883 944 71925 953
rect 71980 944 72020 953
rect 71883 904 71884 944
rect 71924 904 71980 944
rect 71883 895 71925 904
rect 71980 895 72020 904
rect 72075 944 72117 953
rect 72075 904 72076 944
rect 72116 904 72117 944
rect 72075 895 72117 904
rect 71883 776 71925 785
rect 71883 736 71884 776
rect 71924 736 71925 776
rect 71883 727 71925 736
rect 71787 608 71829 617
rect 71787 568 71788 608
rect 71828 568 71829 608
rect 71787 559 71829 568
rect 71788 365 71828 559
rect 71787 356 71829 365
rect 71787 316 71788 356
rect 71828 316 71829 356
rect 71787 307 71829 316
rect 71884 80 71924 727
rect 72076 80 72116 895
rect 72172 785 72212 3172
rect 72460 3137 72500 3331
rect 72652 3330 72692 3415
rect 72844 3330 72884 3415
rect 73036 3389 73076 3424
rect 73035 3380 73077 3389
rect 73035 3340 73036 3380
rect 73076 3340 73172 3380
rect 73035 3331 73077 3340
rect 72556 3212 72596 3221
rect 72940 3212 72980 3221
rect 72459 3128 72501 3137
rect 72459 3088 72460 3128
rect 72500 3088 72501 3128
rect 72459 3079 72501 3088
rect 72556 2540 72596 3172
rect 72364 2500 72596 2540
rect 72748 3172 72940 3212
rect 72268 1373 72308 1458
rect 72267 1364 72309 1373
rect 72267 1324 72268 1364
rect 72308 1324 72309 1364
rect 72267 1315 72309 1324
rect 72267 1112 72309 1121
rect 72267 1072 72268 1112
rect 72308 1072 72309 1112
rect 72267 1063 72309 1072
rect 72268 978 72308 1063
rect 72171 776 72213 785
rect 72364 776 72404 2500
rect 72748 1364 72788 3172
rect 72940 3163 72980 3172
rect 73132 2717 73172 3340
rect 72939 2708 72981 2717
rect 72939 2668 72940 2708
rect 72980 2668 72981 2708
rect 72939 2659 72981 2668
rect 73131 2708 73173 2717
rect 73131 2668 73132 2708
rect 73172 2668 73173 2708
rect 73131 2659 73173 2668
rect 72940 2624 72980 2659
rect 72940 2573 72980 2584
rect 73132 2624 73172 2659
rect 73132 2574 73172 2584
rect 73324 2624 73364 3583
rect 73707 3212 73749 3221
rect 73707 3172 73708 3212
rect 73748 3172 73749 3212
rect 73707 3163 73749 3172
rect 73515 2708 73557 2717
rect 73515 2668 73516 2708
rect 73556 2668 73557 2708
rect 73515 2659 73557 2668
rect 73324 2549 73364 2584
rect 73516 2624 73556 2659
rect 73708 2633 73748 3163
rect 73899 2708 73941 2717
rect 73899 2668 73900 2708
rect 73940 2668 73941 2708
rect 73899 2659 73941 2668
rect 73901 2647 73941 2659
rect 73516 2573 73556 2584
rect 73707 2624 73749 2633
rect 73707 2584 73708 2624
rect 73748 2584 73749 2624
rect 73707 2575 73749 2584
rect 73901 2574 73941 2607
rect 73036 2540 73076 2549
rect 73036 1448 73076 2500
rect 73323 2540 73365 2549
rect 73323 2500 73324 2540
rect 73364 2500 73365 2540
rect 73323 2491 73365 2500
rect 73420 2540 73460 2549
rect 73420 1448 73460 2500
rect 73804 2540 73844 2549
rect 73804 1448 73844 2500
rect 73996 1457 74036 3928
rect 74092 3919 74132 3928
rect 74764 3919 74804 3928
rect 74956 3464 74996 3473
rect 74668 3424 74956 3464
rect 75052 3464 75092 4012
rect 80332 4002 80372 4087
rect 80428 4052 80468 4061
rect 77931 3800 77973 3809
rect 77931 3760 77932 3800
rect 77972 3760 77973 3800
rect 77931 3751 77973 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 76011 3716 76053 3725
rect 76011 3676 76012 3716
rect 76052 3676 76053 3716
rect 76011 3667 76053 3676
rect 76779 3716 76821 3725
rect 76779 3676 76780 3716
rect 76820 3676 76821 3716
rect 76779 3667 76821 3676
rect 75147 3464 75189 3473
rect 75052 3424 75148 3464
rect 75188 3424 75189 3464
rect 74091 2708 74133 2717
rect 74091 2668 74092 2708
rect 74132 2668 74133 2708
rect 74091 2659 74133 2668
rect 74092 2624 74132 2659
rect 74092 2573 74132 2584
rect 74284 2603 74324 2635
rect 74284 2549 74324 2563
rect 74188 2540 74228 2549
rect 72556 1324 72788 1364
rect 72940 1408 73076 1448
rect 73324 1408 73460 1448
rect 73708 1408 73844 1448
rect 73995 1448 74037 1457
rect 74188 1448 74228 2500
rect 74283 2540 74325 2549
rect 74283 2500 74284 2540
rect 74324 2500 74325 2540
rect 74283 2491 74325 2500
rect 74668 2213 74708 3424
rect 74956 3415 74996 3424
rect 75147 3415 75189 3424
rect 75340 3464 75380 3473
rect 75148 3330 75188 3415
rect 75052 3212 75092 3221
rect 74763 2792 74805 2801
rect 74763 2752 74764 2792
rect 74804 2752 74805 2792
rect 74763 2743 74805 2752
rect 74764 2624 74804 2743
rect 74955 2708 74997 2717
rect 74955 2668 74956 2708
rect 74996 2668 74997 2708
rect 74955 2659 74997 2668
rect 74667 2204 74709 2213
rect 74667 2164 74668 2204
rect 74708 2164 74709 2204
rect 74667 2155 74709 2164
rect 74764 1961 74804 2584
rect 74956 2624 74996 2659
rect 74956 2573 74996 2584
rect 74860 2540 74900 2549
rect 74763 1952 74805 1961
rect 74763 1912 74764 1952
rect 74804 1912 74805 1952
rect 74763 1903 74805 1912
rect 74860 1532 74900 2500
rect 73995 1408 73996 1448
rect 74036 1408 74037 1448
rect 72459 1196 72501 1205
rect 72459 1156 72460 1196
rect 72500 1156 72501 1196
rect 72459 1147 72501 1156
rect 72460 1112 72500 1147
rect 72460 1061 72500 1072
rect 72556 944 72596 1324
rect 72843 1280 72885 1289
rect 72843 1240 72844 1280
rect 72884 1240 72885 1280
rect 72843 1231 72885 1240
rect 72652 1121 72692 1206
rect 72651 1112 72693 1121
rect 72651 1072 72652 1112
rect 72692 1072 72693 1112
rect 72651 1063 72693 1072
rect 72844 1112 72884 1231
rect 72844 1063 72884 1072
rect 72748 944 72788 953
rect 72556 904 72692 944
rect 72171 736 72172 776
rect 72212 736 72213 776
rect 72171 727 72213 736
rect 72268 736 72404 776
rect 72268 80 72308 736
rect 72459 524 72501 533
rect 72459 484 72460 524
rect 72500 484 72501 524
rect 72459 475 72501 484
rect 72460 80 72500 475
rect 72652 80 72692 904
rect 72748 533 72788 904
rect 72843 944 72885 953
rect 72843 904 72844 944
rect 72884 904 72885 944
rect 72940 944 72980 1408
rect 73036 1121 73076 1206
rect 73035 1112 73077 1121
rect 73035 1072 73036 1112
rect 73076 1072 73077 1112
rect 73035 1063 73077 1072
rect 73228 1112 73268 1121
rect 73131 944 73173 953
rect 72940 904 73076 944
rect 72843 895 72885 904
rect 72747 524 72789 533
rect 72747 484 72748 524
rect 72788 484 72789 524
rect 72747 475 72789 484
rect 72844 80 72884 895
rect 73036 80 73076 904
rect 73131 904 73132 944
rect 73172 904 73173 944
rect 73131 895 73173 904
rect 73132 810 73172 895
rect 73228 701 73268 1072
rect 73324 944 73364 1408
rect 73420 1121 73460 1206
rect 73612 1205 73652 1207
rect 73611 1196 73653 1205
rect 73611 1156 73612 1196
rect 73652 1156 73653 1196
rect 73611 1147 73653 1156
rect 73419 1112 73461 1121
rect 73419 1072 73420 1112
rect 73460 1072 73461 1112
rect 73419 1063 73461 1072
rect 73612 1112 73652 1147
rect 73612 1063 73652 1072
rect 73516 944 73556 953
rect 73324 904 73460 944
rect 73227 692 73269 701
rect 73227 652 73228 692
rect 73268 652 73269 692
rect 73227 643 73269 652
rect 73131 440 73173 449
rect 73228 440 73268 643
rect 73323 524 73365 533
rect 73323 484 73324 524
rect 73364 484 73365 524
rect 73323 475 73365 484
rect 73131 400 73132 440
rect 73172 400 73268 440
rect 73131 391 73173 400
rect 73324 272 73364 475
rect 73228 232 73364 272
rect 73228 80 73268 232
rect 73420 80 73460 904
rect 73516 533 73556 904
rect 73611 944 73653 953
rect 73611 904 73612 944
rect 73652 904 73653 944
rect 73708 944 73748 1408
rect 73995 1399 74037 1408
rect 74092 1408 74228 1448
rect 74476 1492 74900 1532
rect 73804 1121 73844 1206
rect 73995 1196 74037 1205
rect 73995 1156 73996 1196
rect 74036 1156 74037 1196
rect 73995 1147 74037 1156
rect 73803 1112 73845 1121
rect 73803 1072 73804 1112
rect 73844 1072 73845 1112
rect 73803 1063 73845 1072
rect 73996 1112 74036 1147
rect 73996 1061 74036 1072
rect 73899 944 73941 953
rect 73708 904 73844 944
rect 73611 895 73653 904
rect 73515 524 73557 533
rect 73515 484 73516 524
rect 73556 484 73557 524
rect 73515 475 73557 484
rect 73612 80 73652 895
rect 73804 80 73844 904
rect 73899 904 73900 944
rect 73940 904 73941 944
rect 74092 944 74132 1408
rect 74188 1121 74228 1206
rect 74187 1112 74229 1121
rect 74187 1072 74188 1112
rect 74228 1072 74229 1112
rect 74187 1063 74229 1072
rect 74380 1112 74420 1121
rect 74380 953 74420 1072
rect 74284 944 74324 953
rect 74092 904 74228 944
rect 73899 895 73941 904
rect 73900 810 73940 895
rect 73995 272 74037 281
rect 73995 232 73996 272
rect 74036 232 74037 272
rect 73995 223 74037 232
rect 73996 80 74036 223
rect 74188 80 74228 904
rect 74284 281 74324 904
rect 74379 944 74421 953
rect 74379 904 74380 944
rect 74420 904 74421 944
rect 74379 895 74421 904
rect 74476 860 74516 1492
rect 74955 1448 74997 1457
rect 74955 1408 74956 1448
rect 74996 1408 74997 1448
rect 74955 1399 74997 1408
rect 74859 1364 74901 1373
rect 74859 1324 74860 1364
rect 74900 1324 74901 1364
rect 74859 1315 74901 1324
rect 74764 1121 74804 1206
rect 74571 1112 74613 1121
rect 74571 1072 74572 1112
rect 74612 1072 74613 1112
rect 74571 1063 74613 1072
rect 74763 1112 74805 1121
rect 74763 1072 74764 1112
rect 74804 1072 74805 1112
rect 74763 1063 74805 1072
rect 74572 978 74612 1063
rect 74668 944 74708 953
rect 74476 820 74612 860
rect 74379 524 74421 533
rect 74379 484 74380 524
rect 74420 484 74421 524
rect 74379 475 74421 484
rect 74283 272 74325 281
rect 74283 232 74284 272
rect 74324 232 74325 272
rect 74283 223 74325 232
rect 74380 80 74420 475
rect 74572 80 74612 820
rect 74668 533 74708 904
rect 74763 944 74805 953
rect 74763 904 74764 944
rect 74804 904 74805 944
rect 74860 944 74900 1315
rect 74956 1121 74996 1399
rect 75052 1373 75092 3172
rect 75340 2885 75380 3424
rect 75531 3464 75573 3473
rect 75531 3424 75532 3464
rect 75572 3424 75573 3464
rect 75531 3415 75573 3424
rect 75819 3464 75861 3473
rect 75819 3424 75820 3464
rect 75860 3424 75861 3464
rect 75819 3415 75861 3424
rect 76012 3464 76052 3667
rect 75532 3330 75572 3415
rect 75436 3212 75476 3221
rect 75339 2876 75381 2885
rect 75339 2836 75340 2876
rect 75380 2836 75381 2876
rect 75339 2827 75381 2836
rect 75340 2381 75380 2827
rect 75339 2372 75381 2381
rect 75339 2332 75340 2372
rect 75380 2332 75381 2372
rect 75339 2323 75381 2332
rect 75436 1616 75476 3172
rect 75628 2633 75668 2718
rect 75820 2717 75860 3415
rect 76012 3389 76052 3424
rect 76203 3464 76245 3473
rect 76203 3424 76204 3464
rect 76244 3424 76245 3464
rect 76203 3415 76245 3424
rect 76396 3464 76436 3473
rect 76011 3380 76053 3389
rect 76011 3340 76012 3380
rect 76052 3340 76053 3380
rect 76011 3331 76053 3340
rect 76204 3330 76244 3415
rect 76396 3305 76436 3424
rect 76587 3464 76629 3473
rect 76780 3464 76820 3667
rect 77932 3557 77972 3751
rect 77643 3548 77685 3557
rect 77643 3508 77644 3548
rect 77684 3508 77685 3548
rect 77643 3499 77685 3508
rect 77931 3548 77973 3557
rect 77931 3508 77932 3548
rect 77972 3508 77973 3548
rect 77931 3499 77973 3508
rect 76587 3424 76588 3464
rect 76628 3424 76629 3464
rect 76587 3415 76629 3424
rect 76684 3424 76780 3464
rect 76588 3330 76628 3415
rect 76395 3296 76437 3305
rect 76395 3256 76396 3296
rect 76436 3256 76437 3296
rect 76395 3247 76437 3256
rect 76108 3212 76148 3221
rect 75819 2708 75861 2717
rect 75819 2668 75820 2708
rect 75860 2668 75861 2708
rect 75819 2659 75861 2668
rect 75627 2624 75669 2633
rect 75627 2584 75628 2624
rect 75668 2584 75669 2624
rect 75627 2575 75669 2584
rect 75820 2624 75860 2659
rect 75820 2574 75860 2584
rect 75244 1576 75476 1616
rect 75724 2540 75764 2549
rect 76108 2540 76148 3172
rect 76396 2969 76436 3247
rect 76492 3212 76532 3221
rect 76395 2960 76437 2969
rect 76395 2920 76396 2960
rect 76436 2920 76437 2960
rect 76395 2911 76437 2920
rect 75051 1364 75093 1373
rect 75051 1324 75052 1364
rect 75092 1324 75093 1364
rect 75051 1315 75093 1324
rect 74955 1112 74997 1121
rect 74955 1072 74956 1112
rect 74996 1072 74997 1112
rect 74955 1063 74997 1072
rect 75148 1112 75188 1121
rect 75051 944 75093 953
rect 74860 904 74996 944
rect 74763 895 74805 904
rect 74667 524 74709 533
rect 74667 484 74668 524
rect 74708 484 74709 524
rect 74667 475 74709 484
rect 74764 80 74804 895
rect 74956 80 74996 904
rect 75051 904 75052 944
rect 75092 904 75093 944
rect 75051 895 75093 904
rect 75052 810 75092 895
rect 75148 869 75188 1072
rect 75244 944 75284 1576
rect 75724 1364 75764 2500
rect 75628 1324 75764 1364
rect 76012 2500 76148 2540
rect 75531 1280 75573 1289
rect 75531 1240 75532 1280
rect 75572 1240 75573 1280
rect 75531 1231 75573 1240
rect 75340 1121 75380 1207
rect 75339 1113 75381 1121
rect 75339 1072 75340 1113
rect 75380 1072 75381 1113
rect 75339 1063 75381 1072
rect 75532 1112 75572 1231
rect 75532 1063 75572 1072
rect 75436 944 75476 953
rect 75244 904 75380 944
rect 75147 860 75189 869
rect 75147 820 75148 860
rect 75188 820 75189 860
rect 75147 811 75189 820
rect 75147 524 75189 533
rect 75147 484 75148 524
rect 75188 484 75189 524
rect 75147 475 75189 484
rect 75148 80 75188 475
rect 75340 80 75380 904
rect 75436 533 75476 904
rect 75531 944 75573 953
rect 75531 904 75532 944
rect 75572 904 75573 944
rect 75628 944 75668 1324
rect 75724 1121 75764 1206
rect 75723 1112 75765 1121
rect 75723 1072 75724 1112
rect 75764 1072 75765 1112
rect 75723 1063 75765 1072
rect 75915 1112 75957 1121
rect 75915 1072 75916 1112
rect 75956 1072 75957 1112
rect 75915 1063 75957 1072
rect 75916 978 75956 1063
rect 75819 944 75861 953
rect 75628 904 75764 944
rect 75531 895 75573 904
rect 75435 524 75477 533
rect 75435 484 75436 524
rect 75476 484 75477 524
rect 75435 475 75477 484
rect 75532 80 75572 895
rect 75724 80 75764 904
rect 75819 904 75820 944
rect 75860 904 75861 944
rect 76012 944 76052 2500
rect 76492 1280 76532 3172
rect 76684 3053 76724 3424
rect 76780 3415 76820 3424
rect 76971 3464 77013 3473
rect 76971 3424 76972 3464
rect 77012 3424 77013 3464
rect 76971 3415 77013 3424
rect 77451 3464 77493 3473
rect 77451 3424 77452 3464
rect 77492 3424 77493 3464
rect 77451 3415 77493 3424
rect 77644 3464 77684 3499
rect 76876 3212 76916 3221
rect 76780 3172 76876 3212
rect 76683 3044 76725 3053
rect 76683 3004 76684 3044
rect 76724 3004 76725 3044
rect 76683 2995 76725 3004
rect 76396 1240 76532 1280
rect 76108 1121 76148 1206
rect 76300 1121 76340 1206
rect 76396 1196 76436 1240
rect 76396 1156 76437 1196
rect 76107 1112 76149 1121
rect 76107 1072 76108 1112
rect 76148 1072 76149 1112
rect 76107 1063 76149 1072
rect 76299 1112 76341 1121
rect 76299 1072 76300 1112
rect 76340 1072 76341 1112
rect 76397 1101 76437 1156
rect 76299 1063 76341 1072
rect 76396 1061 76437 1101
rect 76492 1101 76532 1123
rect 76204 944 76244 953
rect 76012 904 76148 944
rect 75819 895 75861 904
rect 75820 810 75860 895
rect 75915 524 75957 533
rect 75915 484 75916 524
rect 75956 484 75957 524
rect 75915 475 75957 484
rect 75916 80 75956 475
rect 76108 80 76148 904
rect 76204 533 76244 904
rect 76299 944 76341 953
rect 76299 904 76300 944
rect 76340 904 76341 944
rect 76299 895 76341 904
rect 76203 524 76245 533
rect 76203 484 76204 524
rect 76244 484 76245 524
rect 76203 475 76245 484
rect 76300 80 76340 895
rect 76396 860 76436 1061
rect 76492 1037 76532 1061
rect 76684 1112 76724 1121
rect 76491 1028 76533 1037
rect 76491 988 76492 1028
rect 76532 988 76533 1028
rect 76491 979 76533 988
rect 76587 944 76629 953
rect 76587 904 76588 944
rect 76628 904 76629 944
rect 76587 895 76629 904
rect 76396 820 76532 860
rect 76492 80 76532 820
rect 76588 810 76628 895
rect 76684 869 76724 1072
rect 76683 860 76725 869
rect 76683 820 76684 860
rect 76724 820 76725 860
rect 76780 860 76820 3172
rect 76876 3163 76916 3172
rect 76972 2624 77012 3415
rect 77452 3330 77492 3415
rect 77644 3413 77684 3424
rect 77932 3464 77972 3499
rect 77932 3414 77972 3424
rect 78123 3464 78165 3473
rect 78316 3464 78356 3473
rect 78123 3424 78124 3464
rect 78164 3424 78165 3464
rect 78123 3415 78165 3424
rect 78220 3424 78316 3464
rect 78124 3330 78164 3415
rect 77548 3212 77588 3221
rect 77260 2633 77300 2718
rect 77068 2624 77108 2633
rect 76972 2584 77068 2624
rect 77068 2575 77108 2584
rect 77259 2624 77301 2633
rect 77259 2584 77260 2624
rect 77300 2584 77301 2624
rect 77259 2575 77301 2584
rect 77163 2540 77205 2549
rect 77163 2500 77164 2540
rect 77204 2500 77205 2540
rect 77163 2491 77205 2500
rect 77164 2406 77204 2491
rect 77451 1616 77493 1625
rect 77451 1576 77452 1616
rect 77492 1576 77493 1616
rect 77451 1567 77493 1576
rect 77067 1532 77109 1541
rect 77067 1492 77068 1532
rect 77108 1492 77109 1532
rect 77067 1483 77109 1492
rect 76876 1112 76916 1123
rect 76876 1037 76916 1072
rect 77068 1112 77108 1483
rect 77260 1112 77300 1123
rect 77108 1072 77204 1112
rect 77068 1063 77108 1072
rect 76875 1028 76917 1037
rect 76875 988 76876 1028
rect 76916 988 76917 1028
rect 76875 979 76917 988
rect 76972 944 77012 953
rect 76780 820 76916 860
rect 76683 811 76725 820
rect 76683 524 76725 533
rect 76683 484 76684 524
rect 76724 484 76725 524
rect 76683 475 76725 484
rect 76684 80 76724 475
rect 76876 80 76916 820
rect 76972 533 77012 904
rect 77067 944 77109 953
rect 77067 904 77068 944
rect 77108 904 77109 944
rect 77067 895 77109 904
rect 76971 524 77013 533
rect 76971 484 76972 524
rect 77012 484 77013 524
rect 76971 475 77013 484
rect 77068 80 77108 895
rect 77164 197 77204 1072
rect 77260 1037 77300 1072
rect 77452 1112 77492 1567
rect 77259 1028 77301 1037
rect 77259 988 77260 1028
rect 77300 988 77301 1028
rect 77259 979 77301 988
rect 77356 953 77396 1038
rect 77452 1037 77492 1072
rect 77451 1028 77493 1037
rect 77451 988 77452 1028
rect 77492 988 77493 1028
rect 77451 979 77493 988
rect 77355 944 77397 953
rect 77355 904 77356 944
rect 77396 904 77397 944
rect 77548 944 77588 3172
rect 78028 3212 78068 3221
rect 78028 2540 78068 3172
rect 78220 3137 78260 3424
rect 78316 3415 78356 3424
rect 78507 3464 78549 3473
rect 78987 3464 79029 3473
rect 78507 3424 78508 3464
rect 78548 3424 78644 3464
rect 78507 3415 78549 3424
rect 78508 3330 78548 3415
rect 78412 3212 78452 3221
rect 78219 3128 78261 3137
rect 78219 3088 78220 3128
rect 78260 3088 78261 3128
rect 78219 3079 78261 3088
rect 77932 2500 78068 2540
rect 77644 1121 77684 1206
rect 77643 1112 77685 1121
rect 77643 1072 77644 1112
rect 77684 1072 77685 1112
rect 77643 1063 77685 1072
rect 77836 1112 77876 1121
rect 77836 1028 77876 1072
rect 77833 988 77876 1028
rect 77740 944 77780 953
rect 77548 904 77684 944
rect 77355 895 77397 904
rect 77259 524 77301 533
rect 77259 484 77260 524
rect 77300 484 77301 524
rect 77259 475 77301 484
rect 77451 524 77493 533
rect 77451 484 77452 524
rect 77492 484 77493 524
rect 77451 475 77493 484
rect 77163 188 77205 197
rect 77163 148 77164 188
rect 77204 148 77205 188
rect 77163 139 77205 148
rect 77260 80 77300 475
rect 77452 80 77492 475
rect 77644 80 77684 904
rect 77833 944 77873 988
rect 77932 944 77972 2500
rect 78220 2465 78260 3079
rect 78412 2540 78452 3172
rect 78604 2624 78644 3424
rect 78987 3424 78988 3464
rect 79028 3424 79029 3464
rect 78987 3415 79029 3424
rect 79179 3464 79221 3473
rect 79179 3424 79180 3464
rect 79220 3424 79221 3464
rect 79179 3415 79221 3424
rect 79372 3464 79412 3473
rect 78988 3305 79028 3415
rect 79180 3330 79220 3415
rect 79372 3305 79412 3424
rect 79564 3464 79604 3473
rect 78987 3296 79029 3305
rect 78987 3256 78988 3296
rect 79028 3256 79029 3296
rect 78987 3247 79029 3256
rect 79371 3296 79413 3305
rect 79371 3256 79372 3296
rect 79412 3256 79413 3296
rect 79371 3247 79413 3256
rect 79084 3212 79124 3221
rect 79468 3212 79508 3221
rect 79124 3172 79220 3212
rect 79084 3163 79124 3172
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 78796 2633 78836 2718
rect 78604 2575 78644 2584
rect 78795 2624 78837 2633
rect 78795 2584 78796 2624
rect 78836 2584 78837 2624
rect 78795 2575 78837 2584
rect 78316 2500 78452 2540
rect 78700 2540 78740 2549
rect 78219 2456 78261 2465
rect 78219 2416 78220 2456
rect 78260 2416 78261 2456
rect 78219 2407 78261 2416
rect 78028 1121 78068 1206
rect 78027 1112 78069 1121
rect 78027 1072 78028 1112
rect 78068 1072 78069 1112
rect 78027 1063 78069 1072
rect 78220 1112 78260 1121
rect 78220 953 78260 1072
rect 78124 944 78164 953
rect 77833 904 77876 944
rect 77932 904 78068 944
rect 77740 533 77780 904
rect 77836 617 77876 904
rect 77835 608 77877 617
rect 77835 568 77836 608
rect 77876 568 77877 608
rect 77835 559 77877 568
rect 77739 524 77781 533
rect 77739 484 77740 524
rect 77780 484 77781 524
rect 77739 475 77781 484
rect 77835 440 77877 449
rect 77835 400 77836 440
rect 77876 400 77877 440
rect 77835 391 77877 400
rect 77836 80 77876 391
rect 78028 80 78068 904
rect 78124 449 78164 904
rect 78219 944 78261 953
rect 78219 904 78220 944
rect 78260 904 78261 944
rect 78316 944 78356 2500
rect 78700 1700 78740 2500
rect 78604 1660 78740 1700
rect 78604 1364 78644 1660
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 78604 1324 78740 1364
rect 78412 1121 78452 1206
rect 78411 1112 78453 1121
rect 78411 1072 78412 1112
rect 78452 1072 78453 1112
rect 78411 1063 78453 1072
rect 78604 1112 78644 1123
rect 78604 1037 78644 1072
rect 78603 1028 78645 1037
rect 78603 988 78604 1028
rect 78644 988 78645 1028
rect 78603 979 78645 988
rect 78508 944 78548 953
rect 78316 904 78452 944
rect 78219 895 78261 904
rect 78123 440 78165 449
rect 78315 440 78357 449
rect 78123 400 78124 440
rect 78164 400 78165 440
rect 78123 391 78165 400
rect 78220 400 78316 440
rect 78356 400 78357 440
rect 78220 80 78260 400
rect 78315 391 78357 400
rect 78412 80 78452 904
rect 78700 944 78740 1324
rect 79180 1289 79220 3172
rect 79360 1289 79400 1308
rect 79179 1280 79221 1289
rect 79360 1280 79413 1289
rect 79179 1240 79180 1280
rect 79220 1240 79221 1280
rect 79179 1231 79221 1240
rect 79276 1240 79372 1280
rect 79412 1240 79413 1280
rect 78796 1121 78836 1206
rect 78795 1112 78837 1121
rect 78795 1072 78796 1112
rect 78836 1072 78837 1112
rect 78795 1063 78837 1072
rect 78988 1112 79028 1121
rect 79180 1112 79220 1121
rect 79028 1072 79124 1112
rect 78988 1063 79028 1072
rect 78892 944 78932 953
rect 78700 904 78836 944
rect 78508 449 78548 904
rect 78603 524 78645 533
rect 78603 484 78604 524
rect 78644 484 78645 524
rect 78603 475 78645 484
rect 78507 440 78549 449
rect 78507 400 78508 440
rect 78548 400 78549 440
rect 78507 391 78549 400
rect 78604 80 78644 475
rect 78796 80 78836 904
rect 78892 533 78932 904
rect 78987 944 79029 953
rect 78987 904 78988 944
rect 79028 904 79029 944
rect 78987 895 79029 904
rect 78891 524 78933 533
rect 78891 484 78892 524
rect 78932 484 78933 524
rect 78891 475 78933 484
rect 78988 80 79028 895
rect 79084 365 79124 1072
rect 79220 1109 79221 1112
rect 79276 1109 79316 1240
rect 79371 1231 79413 1240
rect 79220 1072 79316 1109
rect 79180 1069 79316 1072
rect 79372 1112 79412 1121
rect 79180 1063 79220 1069
rect 79275 944 79317 953
rect 79275 904 79276 944
rect 79316 904 79317 944
rect 79275 895 79317 904
rect 79276 810 79316 895
rect 79372 701 79412 1072
rect 79468 944 79508 3172
rect 79564 2801 79604 3424
rect 79756 3464 79796 3473
rect 79756 3305 79796 3424
rect 79948 3464 79988 3473
rect 79755 3296 79797 3305
rect 79755 3256 79756 3296
rect 79796 3256 79797 3296
rect 79755 3247 79797 3256
rect 79948 3221 79988 3424
rect 80140 3464 80180 3473
rect 80140 3305 80180 3424
rect 80331 3464 80373 3473
rect 80331 3424 80332 3464
rect 80372 3424 80373 3464
rect 80331 3415 80373 3424
rect 80332 3330 80372 3415
rect 80139 3296 80181 3305
rect 80139 3256 80140 3296
rect 80180 3256 80181 3296
rect 80139 3247 80181 3256
rect 79852 3212 79892 3221
rect 79563 2792 79605 2801
rect 79563 2752 79564 2792
rect 79604 2752 79605 2792
rect 79563 2743 79605 2752
rect 79852 1625 79892 3172
rect 79947 3212 79989 3221
rect 79947 3172 79948 3212
rect 79988 3172 79989 3212
rect 79947 3163 79989 3172
rect 80235 3212 80277 3221
rect 80235 3172 80236 3212
rect 80276 3172 80277 3212
rect 80235 3163 80277 3172
rect 79948 2717 79988 3163
rect 80236 3078 80276 3163
rect 79947 2708 79989 2717
rect 79947 2668 79948 2708
rect 79988 2668 79989 2708
rect 79947 2659 79989 2668
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 79948 1952 79988 1963
rect 79948 1877 79988 1912
rect 80140 1952 80180 1961
rect 80180 1912 80372 1952
rect 80140 1903 80180 1912
rect 79947 1868 79989 1877
rect 79947 1828 79948 1868
rect 79988 1828 79989 1868
rect 79947 1819 79989 1828
rect 80140 1700 80180 1709
rect 80180 1660 80276 1700
rect 80140 1651 80180 1660
rect 79851 1616 79893 1625
rect 79851 1576 79852 1616
rect 79892 1576 79893 1616
rect 79851 1567 79893 1576
rect 80043 1616 80085 1625
rect 80043 1576 80044 1616
rect 80084 1576 80085 1616
rect 80043 1567 80085 1576
rect 79755 1532 79797 1541
rect 79755 1492 79756 1532
rect 79796 1492 79797 1532
rect 79755 1483 79797 1492
rect 79563 1280 79605 1289
rect 79563 1240 79564 1280
rect 79604 1240 79605 1280
rect 79563 1231 79605 1240
rect 79564 1121 79604 1231
rect 79563 1112 79605 1121
rect 79563 1072 79564 1112
rect 79604 1072 79605 1112
rect 79563 1063 79605 1072
rect 79756 1112 79796 1483
rect 80044 1373 80084 1567
rect 80043 1364 80085 1373
rect 80043 1324 80044 1364
rect 80084 1324 80180 1364
rect 80043 1315 80085 1324
rect 79948 1121 79988 1206
rect 79756 1063 79796 1072
rect 79947 1112 79989 1121
rect 79947 1072 79948 1112
rect 79988 1072 79989 1112
rect 79947 1063 79989 1072
rect 80140 1112 80180 1324
rect 80140 1063 80180 1072
rect 80044 953 80084 1038
rect 80236 953 80276 1660
rect 80332 1121 80372 1912
rect 80428 1289 80468 4012
rect 80716 3968 80756 4096
rect 80811 4096 80812 4136
rect 80852 4096 80853 4136
rect 80811 4087 80853 4096
rect 86571 4136 86613 4145
rect 86571 4096 86572 4136
rect 86612 4096 86613 4136
rect 86571 4087 86613 4096
rect 86668 4136 86708 4171
rect 80812 4002 80852 4087
rect 80716 3919 80756 3928
rect 81004 3968 81044 3977
rect 86572 3968 86612 4087
rect 86668 4085 86708 4096
rect 87051 4136 87093 4145
rect 87051 4096 87052 4136
rect 87092 4096 87093 4136
rect 87051 4087 87093 4096
rect 87243 4136 87285 4145
rect 87243 4096 87244 4136
rect 87284 4096 87285 4136
rect 87243 4087 87285 4096
rect 91563 4136 91605 4145
rect 91563 4096 91564 4136
rect 91604 4096 91605 4136
rect 91563 4087 91605 4096
rect 91756 4136 91796 4759
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 92043 4136 92085 4145
rect 91796 4096 91988 4136
rect 91756 4087 91796 4096
rect 87052 4002 87092 4087
rect 87148 4052 87188 4061
rect 81044 3928 81332 3968
rect 80619 3212 80661 3221
rect 80619 3172 80620 3212
rect 80660 3172 80661 3212
rect 80619 3163 80661 3172
rect 80523 1364 80565 1373
rect 80523 1324 80524 1364
rect 80564 1324 80565 1364
rect 80523 1315 80565 1324
rect 80427 1280 80469 1289
rect 80427 1240 80428 1280
rect 80468 1240 80469 1280
rect 80427 1231 80469 1240
rect 80331 1112 80373 1121
rect 80331 1072 80332 1112
rect 80372 1072 80373 1112
rect 80331 1063 80373 1072
rect 80524 1112 80564 1315
rect 80524 1063 80564 1072
rect 80332 978 80372 1063
rect 79660 944 79700 953
rect 79468 904 79604 944
rect 79371 692 79413 701
rect 79371 652 79372 692
rect 79412 652 79413 692
rect 79371 643 79413 652
rect 79179 524 79221 533
rect 79179 484 79180 524
rect 79220 484 79221 524
rect 79179 475 79221 484
rect 79083 356 79125 365
rect 79083 316 79084 356
rect 79124 316 79125 356
rect 79083 307 79125 316
rect 79180 80 79220 475
rect 79371 356 79413 365
rect 79371 316 79372 356
rect 79412 316 79413 356
rect 79371 307 79413 316
rect 79372 80 79412 307
rect 79564 80 79604 904
rect 79660 365 79700 904
rect 79755 944 79797 953
rect 79755 904 79756 944
rect 79796 904 79797 944
rect 79755 895 79797 904
rect 80043 944 80085 953
rect 80043 904 80044 944
rect 80084 904 80085 944
rect 80043 895 80085 904
rect 80235 944 80277 953
rect 80235 904 80236 944
rect 80276 904 80277 944
rect 80235 895 80277 904
rect 80428 944 80468 953
rect 79659 356 79701 365
rect 79659 316 79660 356
rect 79700 316 79701 356
rect 79659 307 79701 316
rect 79756 80 79796 895
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 79947 608 79989 617
rect 79947 568 79948 608
rect 79988 568 79989 608
rect 79947 559 79989 568
rect 79948 80 79988 559
rect 80428 524 80468 904
rect 80523 944 80565 953
rect 80523 904 80524 944
rect 80564 904 80565 944
rect 80523 895 80565 904
rect 80140 484 80468 524
rect 80140 80 80180 484
rect 80331 356 80373 365
rect 80331 316 80332 356
rect 80372 316 80373 356
rect 80331 307 80373 316
rect 80332 80 80372 307
rect 80524 80 80564 895
rect 80620 365 80660 3163
rect 80811 1952 80853 1961
rect 80811 1912 80812 1952
rect 80852 1912 80853 1952
rect 80811 1903 80853 1912
rect 81004 1952 81044 3928
rect 81292 3473 81332 3928
rect 86572 3919 86612 3928
rect 86860 3968 86900 3977
rect 82923 3716 82965 3725
rect 82923 3676 82924 3716
rect 82964 3676 82965 3716
rect 82923 3667 82965 3676
rect 81100 3464 81140 3473
rect 81100 3137 81140 3424
rect 81291 3464 81333 3473
rect 81291 3424 81292 3464
rect 81332 3424 81333 3464
rect 81291 3415 81333 3424
rect 81484 3464 81524 3473
rect 81292 3330 81332 3415
rect 81484 3305 81524 3424
rect 81675 3464 81717 3473
rect 81675 3424 81676 3464
rect 81716 3424 81717 3464
rect 81675 3415 81717 3424
rect 82156 3464 82196 3475
rect 81483 3296 81525 3305
rect 81483 3256 81484 3296
rect 81524 3256 81525 3296
rect 81483 3247 81525 3256
rect 81196 3212 81236 3221
rect 81099 3128 81141 3137
rect 81099 3088 81100 3128
rect 81140 3088 81141 3128
rect 81099 3079 81141 3088
rect 81100 2213 81140 3079
rect 81099 2204 81141 2213
rect 81099 2164 81100 2204
rect 81140 2164 81141 2204
rect 81099 2155 81141 2164
rect 81004 1903 81044 1912
rect 80812 1818 80852 1903
rect 80908 1700 80948 1709
rect 80716 1660 80908 1700
rect 80619 356 80661 365
rect 80619 316 80620 356
rect 80660 316 80661 356
rect 80619 307 80661 316
rect 80716 80 80756 1660
rect 80908 1651 80948 1660
rect 80907 1280 80949 1289
rect 80907 1240 80908 1280
rect 80948 1240 80949 1280
rect 80907 1231 80949 1240
rect 81099 1280 81141 1289
rect 81099 1240 81100 1280
rect 81140 1240 81141 1280
rect 81099 1231 81141 1240
rect 80908 1112 80948 1231
rect 80908 1063 80948 1072
rect 81100 1112 81140 1231
rect 81100 1063 81140 1072
rect 81004 944 81044 953
rect 81196 944 81236 3172
rect 81484 2381 81524 3247
rect 81580 3212 81620 3221
rect 81483 2372 81525 2381
rect 81483 2332 81484 2372
rect 81524 2332 81525 2372
rect 81483 2323 81525 2332
rect 81483 1448 81525 1457
rect 81483 1408 81484 1448
rect 81524 1408 81525 1448
rect 81483 1399 81525 1408
rect 81291 1196 81333 1205
rect 81291 1156 81292 1196
rect 81332 1156 81333 1196
rect 81291 1147 81333 1156
rect 81292 1112 81332 1147
rect 81292 1061 81332 1072
rect 81484 1112 81524 1399
rect 81484 1063 81524 1072
rect 81388 944 81428 953
rect 81580 944 81620 3172
rect 81676 2624 81716 3415
rect 82156 3389 82196 3424
rect 82347 3464 82389 3473
rect 82347 3424 82348 3464
rect 82388 3424 82389 3464
rect 82347 3415 82389 3424
rect 82540 3464 82580 3473
rect 82155 3380 82197 3389
rect 82155 3340 82156 3380
rect 82196 3340 82197 3380
rect 82155 3331 82197 3340
rect 82348 3330 82388 3415
rect 82252 3212 82292 3221
rect 82292 3172 82388 3212
rect 82252 3163 82292 3172
rect 81868 2633 81908 2718
rect 81676 2575 81716 2584
rect 81867 2624 81909 2633
rect 81867 2584 81868 2624
rect 81908 2584 81909 2624
rect 81867 2575 81909 2584
rect 81772 2540 81812 2549
rect 81772 1364 81812 2500
rect 81772 1324 82004 1364
rect 81675 1196 81717 1205
rect 81675 1156 81676 1196
rect 81716 1156 81717 1196
rect 81675 1147 81717 1156
rect 81676 1112 81716 1147
rect 81868 1121 81908 1206
rect 81676 1061 81716 1072
rect 81867 1112 81909 1121
rect 81867 1072 81868 1112
rect 81908 1072 81909 1112
rect 81867 1063 81909 1072
rect 80908 904 81004 944
rect 80908 80 80948 904
rect 81004 895 81044 904
rect 81100 904 81236 944
rect 81292 904 81388 944
rect 81100 80 81140 904
rect 81292 80 81332 904
rect 81388 895 81428 904
rect 81484 904 81620 944
rect 81772 944 81812 953
rect 81964 944 82004 1324
rect 82059 1196 82101 1205
rect 82059 1156 82060 1196
rect 82100 1156 82101 1196
rect 82059 1147 82101 1156
rect 82060 1112 82100 1147
rect 82252 1121 82292 1206
rect 82060 1061 82100 1072
rect 82251 1112 82293 1121
rect 82251 1072 82252 1112
rect 82292 1072 82293 1112
rect 82251 1063 82293 1072
rect 82156 944 82196 953
rect 82348 944 82388 3172
rect 82540 2969 82580 3424
rect 82731 3464 82773 3473
rect 82731 3424 82732 3464
rect 82772 3424 82773 3464
rect 82731 3415 82773 3424
rect 82924 3464 82964 3667
rect 83787 3632 83829 3641
rect 83787 3592 83788 3632
rect 83828 3592 83829 3632
rect 86860 3632 86900 3928
rect 86860 3592 87092 3632
rect 83787 3583 83829 3592
rect 82924 3415 82964 3424
rect 83115 3464 83157 3473
rect 83595 3464 83637 3473
rect 83115 3424 83116 3464
rect 83156 3424 83252 3464
rect 83115 3415 83157 3424
rect 82732 3330 82772 3415
rect 83116 3330 83156 3415
rect 82636 3212 82676 3221
rect 83020 3212 83060 3221
rect 82676 3172 82772 3212
rect 82636 3163 82676 3172
rect 82539 2960 82581 2969
rect 82539 2920 82540 2960
rect 82580 2920 82581 2960
rect 82539 2911 82581 2920
rect 82443 1196 82485 1205
rect 82443 1156 82444 1196
rect 82484 1156 82485 1196
rect 82443 1147 82485 1156
rect 82444 1112 82484 1147
rect 82636 1121 82676 1206
rect 82444 1061 82484 1072
rect 82635 1112 82677 1121
rect 82635 1072 82636 1112
rect 82676 1072 82677 1112
rect 82635 1063 82677 1072
rect 82540 944 82580 953
rect 82732 944 82772 3172
rect 83060 3172 83156 3212
rect 83020 3163 83060 3172
rect 82828 1373 82868 1458
rect 82827 1364 82869 1373
rect 82827 1324 82828 1364
rect 82868 1324 82869 1364
rect 82827 1315 82869 1324
rect 82827 1196 82869 1205
rect 82827 1156 82828 1196
rect 82868 1156 82869 1196
rect 82827 1147 82869 1156
rect 82828 1112 82868 1147
rect 83020 1121 83060 1206
rect 82828 1061 82868 1072
rect 83019 1112 83061 1121
rect 83019 1072 83020 1112
rect 83060 1072 83061 1112
rect 83019 1063 83061 1072
rect 83116 944 83156 3172
rect 83212 2624 83252 3424
rect 83595 3424 83596 3464
rect 83636 3424 83637 3464
rect 83595 3415 83637 3424
rect 83788 3464 83828 3583
rect 84172 3557 84212 3588
rect 84171 3548 84213 3557
rect 84171 3508 84172 3548
rect 84212 3508 84213 3548
rect 84171 3499 84213 3508
rect 83788 3415 83828 3424
rect 83979 3464 84021 3473
rect 83979 3424 83980 3464
rect 84020 3424 84021 3464
rect 83979 3415 84021 3424
rect 84172 3464 84212 3499
rect 87052 3473 87092 3592
rect 83596 3330 83636 3415
rect 83980 3330 84020 3415
rect 83691 3212 83733 3221
rect 83691 3172 83692 3212
rect 83732 3172 83733 3212
rect 83691 3163 83733 3172
rect 84076 3212 84116 3221
rect 83692 3078 83732 3163
rect 83212 2575 83252 2584
rect 83403 2624 83445 2633
rect 83403 2584 83404 2624
rect 83444 2584 83445 2624
rect 83403 2575 83445 2584
rect 83308 2540 83348 2549
rect 83308 1364 83348 2500
rect 83404 2490 83444 2575
rect 84076 2540 84116 3172
rect 84172 2885 84212 3424
rect 84363 3464 84405 3473
rect 84363 3424 84364 3464
rect 84404 3424 84405 3464
rect 84363 3415 84405 3424
rect 84555 3464 84597 3473
rect 86860 3464 86900 3473
rect 84555 3424 84556 3464
rect 84596 3424 84597 3464
rect 84555 3415 84597 3424
rect 86764 3424 86860 3464
rect 84171 2876 84213 2885
rect 84171 2836 84172 2876
rect 84212 2836 84213 2876
rect 84171 2827 84213 2836
rect 84364 2633 84404 3415
rect 84556 3330 84596 3415
rect 84460 3212 84500 3221
rect 84500 3172 84692 3212
rect 84460 3163 84500 3172
rect 84363 2624 84405 2633
rect 84363 2584 84364 2624
rect 84404 2584 84405 2624
rect 84363 2575 84405 2584
rect 84076 2500 84308 2540
rect 83883 1448 83925 1457
rect 83883 1408 83884 1448
rect 83924 1408 83925 1448
rect 83883 1399 83925 1408
rect 83308 1324 83540 1364
rect 83211 1196 83253 1205
rect 83211 1156 83212 1196
rect 83252 1156 83253 1196
rect 83211 1147 83253 1156
rect 83212 1112 83252 1147
rect 83212 1061 83252 1072
rect 83307 1112 83349 1121
rect 83393 1112 83433 1118
rect 83307 1072 83308 1112
rect 83348 1109 83433 1112
rect 83348 1072 83393 1109
rect 83307 1063 83349 1072
rect 83393 1060 83433 1069
rect 83308 944 83348 953
rect 83500 944 83540 1324
rect 83595 1196 83637 1205
rect 83595 1156 83596 1196
rect 83636 1156 83637 1196
rect 83595 1147 83637 1156
rect 83596 1112 83636 1147
rect 83596 1061 83636 1072
rect 83793 1109 83833 1118
rect 83884 1109 83924 1399
rect 83979 1196 84021 1205
rect 83979 1156 83980 1196
rect 84020 1156 84021 1196
rect 83979 1147 84021 1156
rect 83833 1069 83924 1109
rect 83793 1060 83833 1069
rect 83692 944 83732 953
rect 81484 80 81524 904
rect 81772 524 81812 904
rect 81865 904 82004 944
rect 82060 904 82156 944
rect 81865 776 81905 904
rect 81865 736 81908 776
rect 81676 484 81812 524
rect 81676 80 81716 484
rect 81868 80 81908 736
rect 82060 80 82100 904
rect 82156 895 82196 904
rect 82252 904 82388 944
rect 82444 904 82540 944
rect 82252 80 82292 904
rect 82444 80 82484 904
rect 82540 895 82580 904
rect 82636 904 82772 944
rect 83020 904 83156 944
rect 83212 904 83308 944
rect 82636 80 82676 904
rect 82827 776 82869 785
rect 82827 736 82828 776
rect 82868 736 82869 776
rect 82827 727 82869 736
rect 82828 80 82868 727
rect 83020 80 83060 904
rect 83212 80 83252 904
rect 83308 895 83348 904
rect 83404 904 83540 944
rect 83596 904 83692 944
rect 83404 80 83444 904
rect 83596 80 83636 904
rect 83692 895 83732 904
rect 83787 776 83829 785
rect 83787 736 83788 776
rect 83828 736 83829 776
rect 83787 727 83829 736
rect 83788 80 83828 727
rect 83884 533 83924 1069
rect 83980 1112 84020 1147
rect 84172 1121 84212 1206
rect 83980 1061 84020 1072
rect 84171 1112 84213 1121
rect 84171 1072 84172 1112
rect 84212 1072 84213 1112
rect 84171 1063 84213 1072
rect 84076 944 84116 953
rect 84268 944 84308 2500
rect 84363 1196 84405 1205
rect 84363 1156 84364 1196
rect 84404 1156 84405 1196
rect 84363 1147 84405 1156
rect 84364 1112 84404 1147
rect 84556 1121 84596 1206
rect 84364 1061 84404 1072
rect 84555 1112 84597 1121
rect 84555 1072 84556 1112
rect 84596 1072 84597 1112
rect 84555 1063 84597 1072
rect 84460 944 84500 953
rect 84652 944 84692 3172
rect 84939 2792 84981 2801
rect 84939 2752 84940 2792
rect 84980 2752 84981 2792
rect 84939 2743 84981 2752
rect 86091 2792 86133 2801
rect 86091 2752 86092 2792
rect 86132 2752 86133 2792
rect 86091 2743 86133 2752
rect 84747 2624 84789 2633
rect 84747 2584 84748 2624
rect 84788 2584 84789 2624
rect 84747 2575 84789 2584
rect 84940 2624 84980 2743
rect 85323 2708 85365 2717
rect 85323 2668 85324 2708
rect 85364 2668 85365 2708
rect 85323 2659 85365 2668
rect 84940 2575 84980 2584
rect 85131 2624 85173 2633
rect 85131 2584 85132 2624
rect 85172 2584 85173 2624
rect 85131 2575 85173 2584
rect 85324 2624 85364 2659
rect 85708 2633 85748 2718
rect 85899 2708 85941 2717
rect 85899 2668 85900 2708
rect 85940 2668 85941 2708
rect 85899 2659 85941 2668
rect 84748 2490 84788 2575
rect 84844 2540 84884 2549
rect 84844 1364 84884 2500
rect 85132 2490 85172 2575
rect 85324 2573 85364 2584
rect 85515 2624 85557 2633
rect 85515 2584 85516 2624
rect 85556 2584 85557 2624
rect 85515 2575 85557 2584
rect 85707 2624 85749 2633
rect 85707 2584 85708 2624
rect 85748 2584 85749 2624
rect 85707 2575 85749 2584
rect 85900 2624 85940 2659
rect 85227 2540 85269 2549
rect 85227 2500 85228 2540
rect 85268 2500 85269 2540
rect 85227 2491 85269 2500
rect 85228 2406 85268 2491
rect 85516 2490 85556 2575
rect 85900 2573 85940 2584
rect 86092 2624 86132 2743
rect 86283 2708 86325 2717
rect 86283 2668 86284 2708
rect 86324 2668 86325 2708
rect 86283 2659 86325 2668
rect 86092 2575 86132 2584
rect 86284 2624 86324 2659
rect 86284 2573 86324 2584
rect 86475 2624 86517 2633
rect 86475 2584 86476 2624
rect 86516 2584 86517 2624
rect 86475 2575 86517 2584
rect 85612 2540 85652 2549
rect 85323 1364 85365 1373
rect 85516 1364 85556 1373
rect 84844 1324 85076 1364
rect 84747 1196 84789 1205
rect 84747 1156 84748 1196
rect 84788 1156 84789 1196
rect 84747 1147 84789 1156
rect 84748 1112 84788 1147
rect 84940 1121 84980 1206
rect 84748 1061 84788 1072
rect 84939 1112 84981 1121
rect 84939 1072 84940 1112
rect 84980 1072 84981 1112
rect 84939 1063 84981 1072
rect 84844 944 84884 953
rect 85036 944 85076 1324
rect 85323 1324 85324 1364
rect 85364 1324 85365 1364
rect 85323 1315 85365 1324
rect 85420 1324 85516 1364
rect 85131 1196 85173 1205
rect 85131 1156 85132 1196
rect 85172 1156 85173 1196
rect 85131 1147 85173 1156
rect 85132 1112 85172 1147
rect 85132 1061 85172 1072
rect 85324 1112 85364 1315
rect 85324 1063 85364 1072
rect 85228 944 85268 953
rect 83980 904 84076 944
rect 83883 524 83925 533
rect 83883 484 83884 524
rect 83924 484 83925 524
rect 83883 475 83925 484
rect 83980 80 84020 904
rect 84076 895 84116 904
rect 84172 904 84308 944
rect 84364 904 84460 944
rect 84172 80 84212 904
rect 84364 80 84404 904
rect 84460 895 84500 904
rect 84556 904 84692 944
rect 84748 904 84844 944
rect 84556 80 84596 904
rect 84748 80 84788 904
rect 84844 895 84884 904
rect 84940 904 85076 944
rect 85132 904 85228 944
rect 85420 944 85460 1324
rect 85516 1315 85556 1324
rect 85515 1196 85557 1205
rect 85515 1156 85516 1196
rect 85556 1156 85557 1196
rect 85515 1147 85557 1156
rect 85516 1112 85556 1147
rect 85516 1061 85556 1072
rect 85420 904 85556 944
rect 84940 80 84980 904
rect 85132 80 85172 904
rect 85228 895 85268 904
rect 85323 860 85365 869
rect 85323 820 85324 860
rect 85364 820 85365 860
rect 85323 811 85365 820
rect 85324 80 85364 811
rect 85516 80 85556 904
rect 85612 869 85652 2500
rect 85996 2540 86036 2549
rect 85707 1532 85749 1541
rect 85707 1492 85708 1532
rect 85748 1492 85749 1532
rect 85707 1483 85749 1492
rect 85708 1289 85748 1483
rect 85900 1364 85940 1373
rect 85804 1324 85900 1364
rect 85707 1280 85749 1289
rect 85707 1240 85708 1280
rect 85748 1240 85749 1280
rect 85707 1231 85749 1240
rect 85708 1112 85748 1231
rect 85708 1063 85748 1072
rect 85804 1028 85844 1324
rect 85900 1315 85940 1324
rect 85900 1205 85940 1220
rect 85899 1196 85941 1205
rect 85899 1156 85900 1196
rect 85940 1156 85941 1196
rect 85899 1147 85941 1156
rect 85900 1125 85940 1147
rect 85900 1076 85940 1085
rect 85804 988 85933 1028
rect 85893 944 85933 988
rect 85996 944 86036 2500
rect 86380 2540 86420 2549
rect 86380 2288 86420 2500
rect 86476 2490 86516 2575
rect 86380 2248 86612 2288
rect 86091 1616 86133 1625
rect 86091 1576 86092 1616
rect 86132 1576 86133 1616
rect 86091 1567 86133 1576
rect 86092 1112 86132 1567
rect 86283 1196 86325 1205
rect 86283 1156 86284 1196
rect 86324 1156 86325 1196
rect 86283 1147 86325 1156
rect 86284 1112 86324 1147
rect 86476 1121 86516 1206
rect 86132 1072 86228 1112
rect 86092 1063 86132 1072
rect 85893 904 85940 944
rect 85996 904 86125 944
rect 85611 860 85653 869
rect 85611 820 85612 860
rect 85652 820 85653 860
rect 85611 811 85653 820
rect 85707 776 85749 785
rect 85707 736 85708 776
rect 85748 736 85749 776
rect 85707 727 85749 736
rect 85611 692 85653 701
rect 85611 652 85612 692
rect 85652 652 85653 692
rect 85611 643 85653 652
rect 85612 365 85652 643
rect 85611 356 85653 365
rect 85611 316 85612 356
rect 85652 316 85653 356
rect 85611 307 85653 316
rect 85708 80 85748 727
rect 85900 80 85940 904
rect 86085 860 86125 904
rect 86085 820 86132 860
rect 86092 80 86132 820
rect 86188 365 86228 1072
rect 86284 1061 86324 1072
rect 86475 1112 86517 1121
rect 86475 1072 86476 1112
rect 86516 1072 86517 1112
rect 86475 1063 86517 1072
rect 86380 944 86420 953
rect 86572 944 86612 2248
rect 86764 1961 86804 3424
rect 86860 3415 86900 3424
rect 87051 3464 87093 3473
rect 87051 3424 87052 3464
rect 87092 3424 87093 3464
rect 87051 3415 87093 3424
rect 87052 3330 87092 3415
rect 86956 3212 86996 3221
rect 86860 3172 86956 3212
rect 86763 1952 86805 1961
rect 86763 1912 86764 1952
rect 86804 1912 86805 1952
rect 86763 1903 86805 1912
rect 86860 1364 86900 3172
rect 86956 3163 86996 3172
rect 86860 1324 86996 1364
rect 86667 1196 86709 1205
rect 86667 1156 86668 1196
rect 86708 1156 86709 1196
rect 86667 1147 86709 1156
rect 86668 1112 86708 1147
rect 86860 1121 86900 1206
rect 86668 1061 86708 1072
rect 86859 1112 86901 1121
rect 86859 1072 86860 1112
rect 86900 1072 86901 1112
rect 86859 1063 86901 1072
rect 86764 944 86804 953
rect 86956 944 86996 1324
rect 87046 1196 87088 1205
rect 87046 1156 87047 1196
rect 87087 1156 87092 1196
rect 87046 1147 87092 1156
rect 87052 1112 87092 1147
rect 87148 1112 87188 4012
rect 87244 4002 87284 4087
rect 91564 4002 91604 4087
rect 91659 4052 91701 4061
rect 91659 4012 91660 4052
rect 91700 4012 91701 4052
rect 91659 4003 91701 4012
rect 91660 3918 91700 4003
rect 91948 3968 91988 4096
rect 92043 4096 92044 4136
rect 92084 4096 92085 4136
rect 92043 4087 92085 4096
rect 92044 4002 92084 4087
rect 93579 4052 93621 4061
rect 93579 4012 93580 4052
rect 93620 4012 93621 4052
rect 93579 4003 93621 4012
rect 91948 3919 91988 3928
rect 92236 3968 92276 3977
rect 88779 3800 88821 3809
rect 88779 3760 88780 3800
rect 88820 3760 88821 3800
rect 88779 3751 88821 3760
rect 87627 3548 87669 3557
rect 87627 3508 87628 3548
rect 87668 3508 87669 3548
rect 87627 3499 87669 3508
rect 87244 3464 87284 3473
rect 87244 3137 87284 3424
rect 87435 3464 87477 3473
rect 87435 3424 87436 3464
rect 87476 3424 87477 3464
rect 87435 3415 87477 3424
rect 87628 3464 87668 3499
rect 87436 3330 87476 3415
rect 87628 3305 87668 3424
rect 87819 3464 87861 3473
rect 87819 3424 87820 3464
rect 87860 3424 87861 3464
rect 87819 3415 87861 3424
rect 88012 3464 88052 3473
rect 87820 3330 87860 3415
rect 87627 3296 87669 3305
rect 87627 3256 87628 3296
rect 87668 3256 87669 3296
rect 87627 3247 87669 3256
rect 87340 3212 87380 3221
rect 87243 3128 87285 3137
rect 87243 3088 87244 3128
rect 87284 3088 87285 3128
rect 87243 3079 87285 3088
rect 87244 1121 87284 1206
rect 87243 1112 87285 1121
rect 87148 1072 87244 1112
rect 87284 1072 87285 1112
rect 87052 1063 87092 1072
rect 87243 1063 87285 1072
rect 87148 944 87188 953
rect 87340 944 87380 3172
rect 87724 3212 87764 3221
rect 87627 1280 87669 1289
rect 87627 1240 87628 1280
rect 87668 1240 87669 1280
rect 87627 1231 87669 1240
rect 87436 1121 87476 1206
rect 87435 1112 87477 1121
rect 87435 1072 87436 1112
rect 87476 1072 87477 1112
rect 87435 1063 87477 1072
rect 87628 1112 87668 1231
rect 87628 1063 87668 1072
rect 87532 944 87572 953
rect 87724 944 87764 3172
rect 88012 2717 88052 3424
rect 88203 3464 88245 3473
rect 88203 3424 88204 3464
rect 88244 3424 88245 3464
rect 88203 3415 88245 3424
rect 88396 3464 88436 3475
rect 88204 3330 88244 3415
rect 88396 3389 88436 3424
rect 88587 3464 88629 3473
rect 88587 3424 88588 3464
rect 88628 3424 88629 3464
rect 88587 3415 88629 3424
rect 88780 3464 88820 3751
rect 89163 3716 89205 3725
rect 89163 3676 89164 3716
rect 89204 3676 89205 3716
rect 89163 3667 89205 3676
rect 88395 3380 88437 3389
rect 88395 3340 88396 3380
rect 88436 3340 88437 3380
rect 88395 3331 88437 3340
rect 88588 3330 88628 3415
rect 88108 3212 88148 3221
rect 88011 2708 88053 2717
rect 88011 2668 88012 2708
rect 88052 2668 88053 2708
rect 88011 2659 88053 2668
rect 87820 1121 87860 1206
rect 88011 1196 88053 1205
rect 88011 1156 88012 1196
rect 88052 1156 88053 1196
rect 88011 1147 88053 1156
rect 87819 1112 87861 1121
rect 87819 1072 87820 1112
rect 87860 1072 87861 1112
rect 87819 1063 87861 1072
rect 88012 1112 88052 1147
rect 88012 1061 88052 1072
rect 87916 944 87956 953
rect 88108 944 88148 3172
rect 88492 3212 88532 3221
rect 88395 1448 88437 1457
rect 88395 1408 88396 1448
rect 88436 1408 88437 1448
rect 88395 1399 88437 1408
rect 88204 1121 88244 1206
rect 88396 1125 88436 1399
rect 88203 1112 88245 1121
rect 88203 1072 88204 1112
rect 88244 1072 88245 1112
rect 88396 1076 88436 1085
rect 88203 1063 88245 1072
rect 88300 944 88340 953
rect 88492 944 88532 3172
rect 88780 2969 88820 3424
rect 88971 3464 89013 3473
rect 88971 3424 88972 3464
rect 89012 3424 89013 3464
rect 88971 3415 89013 3424
rect 89164 3464 89204 3667
rect 92236 3641 92276 3928
rect 89931 3632 89973 3641
rect 89931 3592 89932 3632
rect 89972 3592 89973 3632
rect 89931 3583 89973 3592
rect 90699 3632 90741 3641
rect 90699 3592 90700 3632
rect 90740 3592 90741 3632
rect 90699 3583 90741 3592
rect 92235 3632 92277 3641
rect 92235 3592 92236 3632
rect 92276 3592 92277 3632
rect 92235 3583 92277 3592
rect 93099 3632 93141 3641
rect 93099 3592 93100 3632
rect 93140 3592 93141 3632
rect 93099 3583 93141 3592
rect 93483 3632 93525 3641
rect 93483 3592 93484 3632
rect 93524 3592 93525 3632
rect 93483 3583 93525 3592
rect 88972 3330 89012 3415
rect 89164 3305 89204 3424
rect 89355 3464 89397 3473
rect 89355 3424 89356 3464
rect 89396 3424 89397 3464
rect 89355 3415 89397 3424
rect 89548 3464 89588 3473
rect 89356 3330 89396 3415
rect 89163 3296 89205 3305
rect 89163 3256 89164 3296
rect 89204 3256 89205 3296
rect 89163 3247 89205 3256
rect 88876 3212 88916 3221
rect 88779 2960 88821 2969
rect 88779 2920 88780 2960
rect 88820 2920 88821 2960
rect 88779 2911 88821 2920
rect 88779 1364 88821 1373
rect 88779 1324 88780 1364
rect 88820 1324 88821 1364
rect 88779 1315 88821 1324
rect 88588 1121 88628 1206
rect 88587 1112 88629 1121
rect 88587 1072 88588 1112
rect 88628 1072 88629 1112
rect 88587 1063 88629 1072
rect 88780 1112 88820 1315
rect 88780 1063 88820 1072
rect 88684 944 88724 953
rect 88876 944 88916 3172
rect 89260 3212 89300 3221
rect 88972 1121 89012 1206
rect 89163 1196 89205 1205
rect 89163 1156 89164 1196
rect 89204 1156 89205 1196
rect 89163 1147 89205 1156
rect 88971 1112 89013 1121
rect 88971 1072 88972 1112
rect 89012 1072 89013 1112
rect 88971 1063 89013 1072
rect 89164 1112 89204 1147
rect 89164 1061 89204 1072
rect 89068 1028 89108 1037
rect 89068 944 89108 988
rect 86284 904 86380 944
rect 86187 356 86229 365
rect 86187 316 86188 356
rect 86228 316 86229 356
rect 86187 307 86229 316
rect 86284 80 86324 904
rect 86380 895 86420 904
rect 86476 904 86612 944
rect 86668 904 86764 944
rect 86476 80 86516 904
rect 86668 80 86708 904
rect 86764 895 86804 904
rect 86860 904 86996 944
rect 87052 904 87148 944
rect 86860 80 86900 904
rect 87052 80 87092 904
rect 87148 895 87188 904
rect 87244 904 87380 944
rect 87436 904 87532 944
rect 87244 80 87284 904
rect 87436 80 87476 904
rect 87532 895 87572 904
rect 87628 904 87764 944
rect 87820 904 87916 944
rect 87628 80 87668 904
rect 87820 80 87860 904
rect 87916 895 87956 904
rect 88012 904 88148 944
rect 88204 904 88300 944
rect 88012 80 88052 904
rect 88204 80 88244 904
rect 88300 895 88340 904
rect 88396 904 88532 944
rect 88588 904 88684 944
rect 88396 80 88436 904
rect 88588 80 88628 904
rect 88684 895 88724 904
rect 88780 904 88916 944
rect 88972 904 89108 944
rect 88780 80 88820 904
rect 88972 80 89012 904
rect 89260 776 89300 3172
rect 89548 2633 89588 3424
rect 89739 3464 89781 3473
rect 89739 3424 89740 3464
rect 89780 3424 89781 3464
rect 89739 3415 89781 3424
rect 89932 3464 89972 3583
rect 89740 3330 89780 3415
rect 89932 3221 89972 3424
rect 90123 3464 90165 3473
rect 90123 3424 90124 3464
rect 90164 3424 90165 3464
rect 90123 3415 90165 3424
rect 90316 3464 90356 3473
rect 90124 3330 90164 3415
rect 89644 3212 89684 3221
rect 89547 2624 89589 2633
rect 89547 2584 89548 2624
rect 89588 2584 89589 2624
rect 89547 2575 89589 2584
rect 89355 1364 89397 1373
rect 89355 1324 89356 1364
rect 89396 1324 89397 1364
rect 89355 1315 89397 1324
rect 89356 1121 89396 1315
rect 89547 1196 89589 1205
rect 89547 1156 89548 1196
rect 89588 1156 89589 1196
rect 89547 1147 89589 1156
rect 89355 1112 89397 1121
rect 89355 1072 89356 1112
rect 89396 1072 89397 1112
rect 89355 1063 89397 1072
rect 89548 1112 89588 1147
rect 89548 1061 89588 1072
rect 89452 944 89492 953
rect 89644 944 89684 3172
rect 89931 3212 89973 3221
rect 89931 3172 89932 3212
rect 89972 3172 89973 3212
rect 89931 3163 89973 3172
rect 90028 3212 90068 3221
rect 89739 1364 89781 1373
rect 89739 1324 89740 1364
rect 89780 1324 89781 1364
rect 89739 1315 89781 1324
rect 89740 1112 89780 1315
rect 89931 1280 89973 1289
rect 89931 1240 89932 1280
rect 89972 1240 89973 1280
rect 89931 1231 89973 1240
rect 89740 1063 89780 1072
rect 89932 1112 89972 1231
rect 89932 1063 89972 1072
rect 89836 944 89876 953
rect 90028 944 90068 3172
rect 90316 3053 90356 3424
rect 90507 3464 90549 3473
rect 90507 3424 90508 3464
rect 90548 3424 90549 3464
rect 90507 3415 90549 3424
rect 90700 3464 90740 3583
rect 90700 3415 90740 3424
rect 90891 3464 90933 3473
rect 90891 3424 90892 3464
rect 90932 3424 90933 3464
rect 90891 3415 90933 3424
rect 91084 3464 91124 3473
rect 90508 3330 90548 3415
rect 90892 3330 90932 3415
rect 90412 3212 90452 3221
rect 90315 3044 90357 3053
rect 90315 3004 90316 3044
rect 90356 3004 90357 3044
rect 90315 2995 90357 3004
rect 90316 2885 90356 2995
rect 90315 2876 90357 2885
rect 90315 2836 90316 2876
rect 90356 2836 90357 2876
rect 90315 2827 90357 2836
rect 90123 1364 90165 1373
rect 90123 1324 90124 1364
rect 90164 1324 90165 1364
rect 90123 1315 90165 1324
rect 90124 1112 90164 1315
rect 90315 1280 90357 1289
rect 90315 1240 90316 1280
rect 90356 1240 90357 1280
rect 90315 1231 90357 1240
rect 90124 1063 90164 1072
rect 90316 1112 90356 1231
rect 90316 1063 90356 1072
rect 90220 944 90260 953
rect 90412 944 90452 3172
rect 90796 3212 90836 3221
rect 90507 1364 90549 1373
rect 90507 1324 90508 1364
rect 90548 1324 90549 1364
rect 90507 1315 90549 1324
rect 90508 1112 90548 1315
rect 90508 1063 90548 1072
rect 90700 1101 90740 1123
rect 90700 1037 90740 1061
rect 90699 1028 90741 1037
rect 90699 988 90700 1028
rect 90740 988 90741 1028
rect 90699 979 90741 988
rect 90604 944 90644 953
rect 89164 736 89300 776
rect 89356 904 89452 944
rect 89164 80 89204 736
rect 89356 80 89396 904
rect 89452 895 89492 904
rect 89548 904 89684 944
rect 89740 904 89836 944
rect 89548 80 89588 904
rect 89740 80 89780 904
rect 89836 895 89876 904
rect 89932 904 90068 944
rect 90124 904 90220 944
rect 89932 80 89972 904
rect 90124 80 90164 904
rect 90220 895 90260 904
rect 90316 904 90452 944
rect 90508 904 90604 944
rect 90316 80 90356 904
rect 90508 80 90548 904
rect 90604 895 90644 904
rect 90796 440 90836 3172
rect 91084 2549 91124 3424
rect 91275 3464 91317 3473
rect 91275 3424 91276 3464
rect 91316 3424 91317 3464
rect 91275 3415 91317 3424
rect 91468 3464 91508 3473
rect 91276 3330 91316 3415
rect 91180 3212 91220 3221
rect 91083 2540 91125 2549
rect 91083 2500 91084 2540
rect 91124 2500 91125 2540
rect 91083 2491 91125 2500
rect 91084 2381 91124 2491
rect 91083 2372 91125 2381
rect 91083 2332 91084 2372
rect 91124 2332 91125 2372
rect 91083 2323 91125 2332
rect 90891 1364 90933 1373
rect 90891 1324 90892 1364
rect 90932 1324 90933 1364
rect 90891 1315 90933 1324
rect 90892 1112 90932 1315
rect 91084 1121 91124 1206
rect 90892 1063 90932 1072
rect 91083 1112 91125 1121
rect 91083 1072 91084 1112
rect 91124 1072 91125 1112
rect 91083 1063 91125 1072
rect 90988 944 91028 953
rect 91180 944 91220 3172
rect 91468 2885 91508 3424
rect 91659 3464 91701 3473
rect 91659 3424 91660 3464
rect 91700 3424 91701 3464
rect 91659 3415 91701 3424
rect 91852 3464 91892 3473
rect 91660 3330 91700 3415
rect 91564 3212 91604 3221
rect 91467 2876 91509 2885
rect 91467 2836 91468 2876
rect 91508 2836 91509 2876
rect 91467 2827 91509 2836
rect 91275 1364 91317 1373
rect 91275 1324 91276 1364
rect 91316 1324 91317 1364
rect 91275 1315 91317 1324
rect 91276 1112 91316 1315
rect 91468 1121 91508 1206
rect 91276 1063 91316 1072
rect 91467 1112 91509 1121
rect 91467 1072 91468 1112
rect 91508 1072 91509 1112
rect 91467 1063 91509 1072
rect 91372 1028 91412 1037
rect 91372 944 91412 988
rect 91564 944 91604 3172
rect 91852 2717 91892 3424
rect 92043 3464 92085 3473
rect 92043 3424 92044 3464
rect 92084 3424 92085 3464
rect 92043 3415 92085 3424
rect 92236 3464 92276 3473
rect 92044 3330 92084 3415
rect 91948 3212 91988 3221
rect 91851 2708 91893 2717
rect 91851 2668 91852 2708
rect 91892 2668 91893 2708
rect 91851 2659 91893 2668
rect 91659 1364 91701 1373
rect 91659 1324 91660 1364
rect 91700 1324 91701 1364
rect 91659 1315 91701 1324
rect 91660 1112 91700 1315
rect 91852 1121 91892 1206
rect 91660 1063 91700 1072
rect 91851 1112 91893 1121
rect 91851 1072 91852 1112
rect 91892 1072 91893 1112
rect 91851 1063 91893 1072
rect 90700 400 90836 440
rect 90892 904 90988 944
rect 90700 80 90740 400
rect 90892 80 90932 904
rect 90988 895 91028 904
rect 91084 904 91220 944
rect 91276 904 91412 944
rect 91473 904 91604 944
rect 91756 944 91796 953
rect 91948 944 91988 3172
rect 92236 2969 92276 3424
rect 92427 3464 92469 3473
rect 92427 3424 92428 3464
rect 92468 3424 92469 3464
rect 92427 3415 92469 3424
rect 92619 3464 92661 3473
rect 92619 3424 92620 3464
rect 92660 3424 92661 3464
rect 92619 3415 92661 3424
rect 92811 3464 92853 3473
rect 92811 3424 92812 3464
rect 92852 3424 92853 3464
rect 92811 3415 92853 3424
rect 92428 3330 92468 3415
rect 92620 3330 92660 3415
rect 92812 3330 92852 3415
rect 92332 3212 92372 3221
rect 92235 2960 92277 2969
rect 92235 2920 92236 2960
rect 92276 2920 92277 2960
rect 92235 2911 92277 2920
rect 92043 1364 92085 1373
rect 92043 1324 92044 1364
rect 92084 1324 92085 1364
rect 92043 1315 92085 1324
rect 92044 1112 92084 1315
rect 92044 1063 92084 1072
rect 92236 1112 92276 1121
rect 92140 1028 92180 1037
rect 92140 944 92180 988
rect 92236 944 92276 1072
rect 90987 692 91029 701
rect 90987 652 90988 692
rect 91028 652 91029 692
rect 90987 643 91029 652
rect 90988 533 91028 643
rect 90987 524 91029 533
rect 90987 484 90988 524
rect 91028 484 91029 524
rect 90987 475 91029 484
rect 91084 80 91124 904
rect 91276 80 91316 904
rect 91473 860 91513 904
rect 91468 820 91513 860
rect 91468 80 91508 820
rect 91756 524 91796 904
rect 91660 484 91796 524
rect 91852 904 91988 944
rect 92044 904 92180 944
rect 92233 904 92276 944
rect 91660 80 91700 484
rect 91852 80 91892 904
rect 92044 80 92084 904
rect 92233 860 92273 904
rect 92140 820 92273 860
rect 92140 281 92180 820
rect 92332 692 92372 3172
rect 92716 3212 92756 3221
rect 92756 3172 92852 3212
rect 92716 3163 92756 3172
rect 92715 2624 92757 2633
rect 92715 2584 92716 2624
rect 92756 2584 92757 2624
rect 92715 2575 92757 2584
rect 92523 1952 92565 1961
rect 92523 1912 92524 1952
rect 92564 1912 92565 1952
rect 92523 1903 92565 1912
rect 92716 1952 92756 2575
rect 92716 1903 92756 1912
rect 92524 1818 92564 1903
rect 92619 1700 92661 1709
rect 92619 1660 92620 1700
rect 92660 1660 92661 1700
rect 92619 1651 92661 1660
rect 92620 1566 92660 1651
rect 92812 1448 92852 3172
rect 92907 3128 92949 3137
rect 92907 3088 92908 3128
rect 92948 3088 92949 3128
rect 92907 3079 92949 3088
rect 92908 2624 92948 3079
rect 93100 2633 93140 3583
rect 93291 3464 93333 3473
rect 93291 3424 93292 3464
rect 93332 3424 93333 3464
rect 93291 3415 93333 3424
rect 93484 3464 93524 3583
rect 93484 3415 93524 3424
rect 93292 3330 93332 3415
rect 93388 3212 93428 3221
rect 93292 3172 93388 3212
rect 92908 2575 92948 2584
rect 93099 2624 93141 2633
rect 93099 2584 93100 2624
rect 93140 2584 93141 2624
rect 93099 2575 93141 2584
rect 93004 2540 93044 2549
rect 93004 2465 93044 2500
rect 93100 2490 93140 2575
rect 93003 2456 93045 2465
rect 93003 2416 93004 2456
rect 93044 2416 93045 2456
rect 93003 2407 93045 2416
rect 93004 2405 93044 2407
rect 93099 1700 93141 1709
rect 93099 1660 93100 1700
rect 93140 1660 93141 1700
rect 93099 1651 93141 1660
rect 92716 1408 92852 1448
rect 92427 1364 92469 1373
rect 92427 1324 92428 1364
rect 92468 1324 92469 1364
rect 92427 1315 92469 1324
rect 92428 1121 92468 1315
rect 92619 1280 92661 1289
rect 92619 1240 92620 1280
rect 92660 1240 92661 1280
rect 92619 1231 92661 1240
rect 92427 1112 92469 1121
rect 92427 1072 92428 1112
rect 92468 1072 92469 1112
rect 92427 1063 92469 1072
rect 92620 1112 92660 1231
rect 92620 1063 92660 1072
rect 92524 944 92564 953
rect 92716 944 92756 1408
rect 92812 1121 92852 1206
rect 92811 1112 92853 1121
rect 92811 1072 92812 1112
rect 92852 1072 92853 1112
rect 92811 1063 92853 1072
rect 93003 1112 93045 1121
rect 93003 1072 93004 1112
rect 93044 1072 93045 1112
rect 93003 1063 93045 1072
rect 93004 978 93044 1063
rect 92908 944 92948 953
rect 92236 652 92372 692
rect 92428 904 92524 944
rect 92139 272 92181 281
rect 92139 232 92140 272
rect 92180 232 92181 272
rect 92139 223 92181 232
rect 92236 80 92276 652
rect 92428 80 92468 904
rect 92524 895 92564 904
rect 92620 904 92756 944
rect 92812 904 92908 944
rect 92620 80 92660 904
rect 92812 80 92852 904
rect 92908 895 92948 904
rect 93100 860 93140 1651
rect 93195 1280 93237 1289
rect 93195 1240 93196 1280
rect 93236 1240 93237 1280
rect 93195 1231 93237 1240
rect 93196 1112 93236 1231
rect 93292 1121 93332 3172
rect 93388 3163 93428 3172
rect 93580 2792 93620 4003
rect 94443 3800 94485 3809
rect 94443 3760 94444 3800
rect 94484 3760 94485 3800
rect 94443 3751 94485 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 94251 3632 94293 3641
rect 94251 3592 94252 3632
rect 94292 3592 94293 3632
rect 94251 3583 94293 3592
rect 94059 3464 94101 3473
rect 94059 3424 94060 3464
rect 94100 3424 94101 3464
rect 94059 3415 94101 3424
rect 94252 3464 94292 3583
rect 94252 3415 94292 3424
rect 94444 3464 94484 3751
rect 94635 3716 94677 3725
rect 94635 3676 94636 3716
rect 94676 3676 94677 3716
rect 94635 3667 94677 3676
rect 94636 3557 94676 3667
rect 94635 3548 94677 3557
rect 94635 3508 94636 3548
rect 94676 3508 94677 3548
rect 94635 3499 94677 3508
rect 95019 3548 95061 3557
rect 95019 3508 95020 3548
rect 95060 3508 95061 3548
rect 95019 3499 95061 3508
rect 95307 3548 95349 3557
rect 95307 3508 95308 3548
rect 95348 3508 95349 3548
rect 95307 3499 95349 3508
rect 95691 3548 95733 3557
rect 95691 3508 95692 3548
rect 95732 3508 95733 3548
rect 95691 3499 95733 3508
rect 96171 3548 96213 3557
rect 96171 3508 96172 3548
rect 96212 3508 96213 3548
rect 96171 3499 96213 3508
rect 96555 3548 96597 3557
rect 96555 3508 96556 3548
rect 96596 3508 96597 3548
rect 96555 3499 96597 3508
rect 94444 3415 94484 3424
rect 94636 3464 94676 3499
rect 94060 3330 94100 3415
rect 94636 3414 94676 3424
rect 94827 3464 94869 3473
rect 94827 3424 94828 3464
rect 94868 3424 94869 3464
rect 94827 3415 94869 3424
rect 95020 3464 95060 3499
rect 94347 3380 94389 3389
rect 94347 3340 94348 3380
rect 94388 3340 94389 3380
rect 94347 3331 94389 3340
rect 94156 3212 94196 3221
rect 94196 3172 94292 3212
rect 94156 3163 94196 3172
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 93388 2752 93620 2792
rect 93388 1229 93428 2752
rect 93675 2708 93717 2717
rect 93580 2668 93676 2708
rect 93716 2668 93717 2708
rect 93580 2624 93620 2668
rect 93675 2659 93717 2668
rect 93580 2575 93620 2584
rect 93771 2624 93813 2633
rect 93771 2584 93772 2624
rect 93812 2584 93813 2624
rect 93771 2575 93813 2584
rect 93676 2540 93716 2549
rect 93483 2456 93525 2465
rect 93483 2416 93484 2456
rect 93524 2416 93525 2456
rect 93483 2407 93525 2416
rect 93388 1121 93435 1229
rect 93196 1063 93236 1072
rect 93291 1112 93333 1121
rect 93291 1072 93292 1112
rect 93332 1072 93333 1112
rect 93291 1063 93333 1072
rect 93388 1112 93436 1121
rect 93435 1072 93436 1112
rect 93388 1063 93436 1072
rect 93292 944 93332 953
rect 93484 944 93524 2407
rect 93676 1280 93716 2500
rect 93772 2490 93812 2575
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 94252 1289 94292 3172
rect 94348 2885 94388 3331
rect 94828 3330 94868 3415
rect 95020 3413 95060 3424
rect 94540 3212 94580 3221
rect 94924 3212 94964 3221
rect 94580 3172 94676 3212
rect 94540 3163 94580 3172
rect 94347 2876 94389 2885
rect 94347 2836 94348 2876
rect 94388 2836 94389 2876
rect 94347 2827 94389 2836
rect 94636 1541 94676 3172
rect 94635 1532 94677 1541
rect 94635 1492 94636 1532
rect 94676 1492 94677 1532
rect 94635 1483 94677 1492
rect 94924 1457 94964 3172
rect 95115 2624 95157 2633
rect 95115 2584 95116 2624
rect 95156 2584 95157 2624
rect 95115 2575 95157 2584
rect 95308 2624 95348 3499
rect 95500 3464 95540 3473
rect 95500 3221 95540 3424
rect 95692 3464 95732 3499
rect 95692 3413 95732 3424
rect 95980 3464 96020 3473
rect 95499 3212 95541 3221
rect 95499 3172 95500 3212
rect 95540 3172 95541 3212
rect 95499 3163 95541 3172
rect 95596 3212 95636 3221
rect 95308 2575 95348 2584
rect 95116 2490 95156 2575
rect 95212 2540 95252 2549
rect 95212 2456 95252 2500
rect 95212 2416 95540 2456
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 95500 2120 95540 2416
rect 95404 2080 95540 2120
rect 94347 1448 94389 1457
rect 94347 1408 94348 1448
rect 94388 1408 94389 1448
rect 94347 1399 94389 1408
rect 94923 1448 94965 1457
rect 94923 1408 94924 1448
rect 94964 1408 94965 1448
rect 94923 1399 94965 1408
rect 94251 1280 94293 1289
rect 93676 1240 93908 1280
rect 93580 1121 93620 1206
rect 93579 1112 93621 1121
rect 93579 1072 93580 1112
rect 93620 1072 93621 1112
rect 93579 1063 93621 1072
rect 93772 1112 93812 1123
rect 93772 1037 93812 1072
rect 93771 1028 93813 1037
rect 93771 988 93772 1028
rect 93812 988 93813 1028
rect 93771 979 93813 988
rect 93868 953 93908 1240
rect 94251 1240 94252 1280
rect 94292 1240 94293 1280
rect 94251 1231 94293 1240
rect 93964 1121 94004 1206
rect 94156 1121 94196 1206
rect 93963 1112 94005 1121
rect 93963 1072 93964 1112
rect 94004 1072 94005 1112
rect 93963 1063 94005 1072
rect 94155 1112 94197 1121
rect 94155 1072 94156 1112
rect 94196 1072 94197 1112
rect 94155 1063 94197 1072
rect 94348 1112 94388 1399
rect 94348 1063 94388 1072
rect 94540 1101 94580 1123
rect 94732 1121 94772 1204
rect 94731 1112 94773 1121
rect 94731 1069 94732 1112
rect 94772 1069 94773 1112
rect 94731 1063 94773 1069
rect 94924 1101 94964 1123
rect 94540 1037 94580 1061
rect 94732 1060 94772 1063
rect 94539 1028 94581 1037
rect 94539 988 94540 1028
rect 94580 988 94581 1028
rect 94539 979 94581 988
rect 94828 953 94868 1038
rect 94924 1037 94964 1061
rect 95116 1101 95156 1118
rect 95116 1037 95156 1061
rect 95308 1101 95348 1123
rect 94923 1028 94965 1037
rect 94923 988 94924 1028
rect 94964 988 94965 1028
rect 94923 979 94965 988
rect 95110 1028 95156 1037
rect 95110 988 95111 1028
rect 95151 988 95156 1028
rect 95110 979 95152 988
rect 95212 953 95252 1038
rect 95308 1037 95348 1061
rect 95307 1028 95349 1037
rect 95307 988 95308 1028
rect 95348 988 95349 1028
rect 95307 979 95349 988
rect 95404 953 95444 2080
rect 95596 1289 95636 3172
rect 95980 3137 96020 3424
rect 96172 3464 96212 3499
rect 96172 3413 96212 3424
rect 96076 3212 96116 3221
rect 96116 3172 96212 3212
rect 96076 3163 96116 3172
rect 95979 3128 96021 3137
rect 95979 3088 95980 3128
rect 96020 3088 96021 3128
rect 95979 3079 96021 3088
rect 96172 2540 96212 3172
rect 96556 2717 96596 3499
rect 98187 3380 98229 3389
rect 98187 3340 98188 3380
rect 98228 3340 98229 3380
rect 98187 3331 98229 3340
rect 98091 2960 98133 2969
rect 98091 2920 98092 2960
rect 98132 2920 98133 2960
rect 98091 2911 98133 2920
rect 97515 2792 97557 2801
rect 97515 2752 97516 2792
rect 97556 2752 97557 2792
rect 97515 2743 97557 2752
rect 96555 2708 96597 2717
rect 96555 2668 96556 2708
rect 96596 2668 96597 2708
rect 96555 2659 96597 2668
rect 96939 2708 96981 2717
rect 96939 2668 96940 2708
rect 96980 2668 96981 2708
rect 96939 2659 96981 2668
rect 97323 2708 97365 2717
rect 97323 2668 97324 2708
rect 97364 2668 97365 2708
rect 97323 2659 97365 2668
rect 96363 2624 96405 2633
rect 96363 2584 96364 2624
rect 96404 2584 96405 2624
rect 96363 2575 96405 2584
rect 96556 2624 96596 2659
rect 96172 2500 96308 2540
rect 96268 1364 96308 2500
rect 96364 2490 96404 2575
rect 96556 2574 96596 2584
rect 96747 2624 96789 2633
rect 96747 2584 96748 2624
rect 96788 2584 96789 2624
rect 96747 2575 96789 2584
rect 96940 2624 96980 2659
rect 96460 2540 96500 2549
rect 96460 1448 96500 2500
rect 96748 2490 96788 2575
rect 96940 2573 96980 2584
rect 97131 2624 97173 2633
rect 97131 2584 97132 2624
rect 97172 2584 97173 2624
rect 97131 2575 97173 2584
rect 97324 2624 97364 2659
rect 96844 2540 96884 2549
rect 96844 1532 96884 2500
rect 97132 2490 97172 2575
rect 97324 2573 97364 2584
rect 97516 2624 97556 2743
rect 97707 2708 97749 2717
rect 97707 2668 97708 2708
rect 97748 2668 97749 2708
rect 97707 2659 97749 2668
rect 97899 2708 97941 2717
rect 97899 2668 97900 2708
rect 97940 2668 97941 2708
rect 97899 2659 97941 2668
rect 97516 2575 97556 2584
rect 97709 2647 97749 2659
rect 97709 2574 97749 2607
rect 97900 2624 97940 2659
rect 97228 2540 97268 2549
rect 97035 1532 97077 1541
rect 96844 1492 97036 1532
rect 97076 1492 97077 1532
rect 97035 1483 97077 1492
rect 96460 1408 96980 1448
rect 96268 1324 96596 1364
rect 95595 1280 95637 1289
rect 95595 1240 95596 1280
rect 95636 1240 95637 1280
rect 95595 1231 95637 1240
rect 96171 1280 96213 1289
rect 96171 1240 96172 1280
rect 96212 1240 96213 1280
rect 96171 1231 96213 1240
rect 95500 1121 95540 1206
rect 95884 1121 95924 1206
rect 96075 1196 96117 1205
rect 96075 1156 96076 1196
rect 96116 1156 96117 1196
rect 96075 1147 96117 1156
rect 95499 1112 95541 1121
rect 95499 1072 95500 1112
rect 95540 1072 95541 1112
rect 95499 1063 95541 1072
rect 95699 1112 95739 1118
rect 95883 1112 95925 1121
rect 95699 1109 95828 1112
rect 95739 1072 95828 1109
rect 95699 1060 95739 1069
rect 93676 944 93716 953
rect 93004 820 93140 860
rect 93196 904 93292 944
rect 93004 80 93044 820
rect 93196 80 93236 904
rect 93292 895 93332 904
rect 93388 904 93524 944
rect 93580 904 93676 944
rect 93388 80 93428 904
rect 93580 80 93620 904
rect 93676 895 93716 904
rect 93867 944 93909 953
rect 94060 944 94100 953
rect 93867 904 93868 944
rect 93908 904 93909 944
rect 93867 895 93909 904
rect 93964 904 94060 944
rect 93771 860 93813 869
rect 93771 820 93772 860
rect 93812 820 93813 860
rect 93771 811 93813 820
rect 93772 80 93812 811
rect 93964 80 94004 904
rect 94060 895 94100 904
rect 94155 944 94197 953
rect 94444 944 94484 953
rect 94155 904 94156 944
rect 94196 904 94197 944
rect 94155 895 94197 904
rect 94348 904 94444 944
rect 94156 80 94196 895
rect 94348 80 94388 904
rect 94444 895 94484 904
rect 94731 944 94773 953
rect 94731 904 94732 944
rect 94772 904 94773 944
rect 94731 895 94773 904
rect 94827 944 94869 953
rect 94827 904 94828 944
rect 94868 904 94869 944
rect 94827 895 94869 904
rect 95211 944 95253 953
rect 95211 904 95212 944
rect 95252 904 95253 944
rect 95211 895 95253 904
rect 95403 944 95445 953
rect 95596 944 95636 953
rect 95403 904 95404 944
rect 95444 904 95445 944
rect 95403 895 95445 904
rect 95500 904 95596 944
rect 94539 860 94581 869
rect 94539 820 94540 860
rect 94580 820 94581 860
rect 94539 811 94581 820
rect 94540 80 94580 811
rect 94635 776 94677 785
rect 94635 736 94636 776
rect 94676 736 94677 776
rect 94635 727 94677 736
rect 94636 617 94676 727
rect 94635 608 94677 617
rect 94635 568 94636 608
rect 94676 568 94677 608
rect 94635 559 94677 568
rect 94732 80 94772 895
rect 94827 776 94869 785
rect 94827 736 94828 776
rect 94868 736 94869 776
rect 94827 727 94869 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
rect 94828 440 94868 727
rect 95307 608 95349 617
rect 95307 568 95308 608
rect 95348 568 95349 608
rect 95307 559 95349 568
rect 94828 400 94964 440
rect 94924 80 94964 400
rect 95115 104 95157 113
rect 95115 80 95116 104
rect 64244 64 64264 80
rect 64184 0 64264 64
rect 64376 0 64456 80
rect 64568 0 64648 80
rect 64760 0 64840 80
rect 64952 0 65032 80
rect 65144 0 65224 80
rect 65336 0 65416 80
rect 65528 0 65608 80
rect 65720 0 65800 80
rect 65912 0 65992 80
rect 66104 0 66184 80
rect 66296 0 66376 80
rect 66488 0 66568 80
rect 66680 0 66760 80
rect 66872 0 66952 80
rect 67064 0 67144 80
rect 67256 0 67336 80
rect 67448 0 67528 80
rect 67640 0 67720 80
rect 67832 0 67912 80
rect 68024 0 68104 80
rect 68216 0 68296 80
rect 68408 0 68488 80
rect 68600 0 68680 80
rect 68792 0 68872 80
rect 68984 0 69064 80
rect 69176 0 69256 80
rect 69368 0 69448 80
rect 69560 0 69640 80
rect 69752 0 69832 80
rect 69944 0 70024 80
rect 70136 0 70216 80
rect 70328 0 70408 80
rect 70520 0 70600 80
rect 70712 0 70792 80
rect 70904 0 70984 80
rect 71096 0 71176 80
rect 71288 0 71368 80
rect 71480 0 71560 80
rect 71672 0 71752 80
rect 71864 0 71944 80
rect 72056 0 72136 80
rect 72248 0 72328 80
rect 72440 0 72520 80
rect 72632 0 72712 80
rect 72824 0 72904 80
rect 73016 0 73096 80
rect 73208 0 73288 80
rect 73400 0 73480 80
rect 73592 0 73672 80
rect 73784 0 73864 80
rect 73976 0 74056 80
rect 74168 0 74248 80
rect 74360 0 74440 80
rect 74552 0 74632 80
rect 74744 0 74824 80
rect 74936 0 75016 80
rect 75128 0 75208 80
rect 75320 0 75400 80
rect 75512 0 75592 80
rect 75704 0 75784 80
rect 75896 0 75976 80
rect 76088 0 76168 80
rect 76280 0 76360 80
rect 76472 0 76552 80
rect 76664 0 76744 80
rect 76856 0 76936 80
rect 77048 0 77128 80
rect 77240 0 77320 80
rect 77432 0 77512 80
rect 77624 0 77704 80
rect 77816 0 77896 80
rect 78008 0 78088 80
rect 78200 0 78280 80
rect 78392 0 78472 80
rect 78584 0 78664 80
rect 78776 0 78856 80
rect 78968 0 79048 80
rect 79160 0 79240 80
rect 79352 0 79432 80
rect 79544 0 79624 80
rect 79736 0 79816 80
rect 79928 0 80008 80
rect 80120 0 80200 80
rect 80312 0 80392 80
rect 80504 0 80584 80
rect 80696 0 80776 80
rect 80888 0 80968 80
rect 81080 0 81160 80
rect 81272 0 81352 80
rect 81464 0 81544 80
rect 81656 0 81736 80
rect 81848 0 81928 80
rect 82040 0 82120 80
rect 82232 0 82312 80
rect 82424 0 82504 80
rect 82616 0 82696 80
rect 82808 0 82888 80
rect 83000 0 83080 80
rect 83192 0 83272 80
rect 83384 0 83464 80
rect 83576 0 83656 80
rect 83768 0 83848 80
rect 83960 0 84040 80
rect 84152 0 84232 80
rect 84344 0 84424 80
rect 84536 0 84616 80
rect 84728 0 84808 80
rect 84920 0 85000 80
rect 85112 0 85192 80
rect 85304 0 85384 80
rect 85496 0 85576 80
rect 85688 0 85768 80
rect 85880 0 85960 80
rect 86072 0 86152 80
rect 86264 0 86344 80
rect 86456 0 86536 80
rect 86648 0 86728 80
rect 86840 0 86920 80
rect 87032 0 87112 80
rect 87224 0 87304 80
rect 87416 0 87496 80
rect 87608 0 87688 80
rect 87800 0 87880 80
rect 87992 0 88072 80
rect 88184 0 88264 80
rect 88376 0 88456 80
rect 88568 0 88648 80
rect 88760 0 88840 80
rect 88952 0 89032 80
rect 89144 0 89224 80
rect 89336 0 89416 80
rect 89528 0 89608 80
rect 89720 0 89800 80
rect 89912 0 89992 80
rect 90104 0 90184 80
rect 90296 0 90376 80
rect 90488 0 90568 80
rect 90680 0 90760 80
rect 90872 0 90952 80
rect 91064 0 91144 80
rect 91256 0 91336 80
rect 91448 0 91528 80
rect 91640 0 91720 80
rect 91832 0 91912 80
rect 92024 0 92104 80
rect 92216 0 92296 80
rect 92408 0 92488 80
rect 92600 0 92680 80
rect 92792 0 92872 80
rect 92984 0 93064 80
rect 93176 0 93256 80
rect 93368 0 93448 80
rect 93560 0 93640 80
rect 93752 0 93832 80
rect 93944 0 94024 80
rect 94136 0 94216 80
rect 94328 0 94408 80
rect 94520 0 94600 80
rect 94712 0 94792 80
rect 94904 0 94984 80
rect 95096 64 95116 80
rect 95156 80 95157 104
rect 95308 80 95348 559
rect 95500 80 95540 904
rect 95596 895 95636 904
rect 95691 944 95733 953
rect 95691 904 95692 944
rect 95732 904 95733 944
rect 95691 895 95733 904
rect 95692 80 95732 895
rect 95788 869 95828 1072
rect 95883 1072 95884 1112
rect 95924 1072 95925 1112
rect 95883 1063 95925 1072
rect 96076 1112 96116 1147
rect 96076 1061 96116 1072
rect 95980 944 96020 953
rect 96172 944 96212 1231
rect 96268 1121 96308 1206
rect 96459 1196 96501 1205
rect 96459 1156 96460 1196
rect 96500 1156 96501 1196
rect 96459 1147 96501 1156
rect 96267 1112 96309 1121
rect 96267 1072 96268 1112
rect 96308 1072 96309 1112
rect 96267 1063 96309 1072
rect 96460 1112 96500 1147
rect 96460 1061 96500 1072
rect 96364 944 96404 953
rect 96556 944 96596 1324
rect 96652 1121 96692 1206
rect 96843 1196 96885 1205
rect 96843 1156 96844 1196
rect 96884 1156 96885 1196
rect 96843 1147 96885 1156
rect 96651 1112 96693 1121
rect 96651 1072 96652 1112
rect 96692 1072 96693 1112
rect 96651 1063 96693 1072
rect 96844 1112 96884 1147
rect 96844 1061 96884 1072
rect 96748 944 96788 953
rect 96940 944 96980 1408
rect 97228 1364 97268 2500
rect 97611 2540 97653 2549
rect 97611 2500 97612 2540
rect 97652 2500 97653 2540
rect 97611 2491 97653 2500
rect 97612 2406 97652 2491
rect 97900 1952 97940 2584
rect 98092 2624 98132 2911
rect 98092 2575 98132 2584
rect 97900 1903 97940 1912
rect 97996 2540 98036 2549
rect 97996 1868 98036 2500
rect 98188 2288 98228 3331
rect 98092 2248 98228 2288
rect 98092 1973 98132 2248
rect 98092 1924 98132 1933
rect 97996 1828 98132 1868
rect 97996 1700 98036 1709
rect 97996 1373 98036 1660
rect 97995 1364 98037 1373
rect 97228 1324 97748 1364
rect 97036 1121 97076 1206
rect 97227 1196 97269 1205
rect 97227 1156 97228 1196
rect 97268 1156 97269 1196
rect 97227 1147 97269 1156
rect 97611 1196 97653 1205
rect 97611 1156 97612 1196
rect 97652 1156 97653 1196
rect 97611 1147 97653 1156
rect 97227 1125 97267 1147
rect 97035 1112 97077 1121
rect 97035 1072 97036 1112
rect 97076 1072 97077 1112
rect 97035 1063 97077 1072
rect 97227 1062 97267 1085
rect 97420 1112 97460 1121
rect 97132 944 97172 953
rect 95884 904 95980 944
rect 95787 860 95829 869
rect 95787 820 95788 860
rect 95828 820 95829 860
rect 95787 811 95829 820
rect 95884 80 95924 904
rect 95980 895 96020 904
rect 96076 904 96212 944
rect 96268 904 96364 944
rect 96076 80 96116 904
rect 96268 80 96308 904
rect 96364 895 96404 904
rect 96460 904 96596 944
rect 96652 904 96748 944
rect 96460 80 96500 904
rect 96652 80 96692 904
rect 96748 895 96788 904
rect 96844 904 96980 944
rect 97036 904 97132 944
rect 96844 80 96884 904
rect 97036 80 97076 904
rect 97132 895 97172 904
rect 97227 776 97269 785
rect 97227 736 97228 776
rect 97268 736 97269 776
rect 97227 727 97269 736
rect 97228 80 97268 727
rect 97420 608 97460 1072
rect 97612 1112 97652 1147
rect 97612 1061 97652 1072
rect 97324 568 97460 608
rect 97516 944 97556 953
rect 97708 944 97748 1324
rect 97995 1324 97996 1364
rect 98036 1324 98037 1364
rect 98092 1364 98132 1828
rect 98380 1364 98420 1373
rect 98092 1324 98324 1364
rect 97995 1315 98037 1324
rect 97995 1196 98037 1205
rect 97995 1156 97996 1196
rect 98036 1156 98037 1196
rect 97995 1147 98037 1156
rect 97995 1125 98035 1147
rect 97324 449 97364 568
rect 97516 524 97556 904
rect 97420 484 97556 524
rect 97612 904 97748 944
rect 97804 1112 97844 1121
rect 97323 440 97365 449
rect 97323 400 97324 440
rect 97364 400 97365 440
rect 97323 391 97365 400
rect 97420 80 97460 484
rect 97612 80 97652 904
rect 97804 860 97844 1072
rect 97995 1062 98035 1085
rect 98188 1112 98228 1121
rect 97900 1028 97940 1037
rect 98188 1028 98228 1072
rect 97708 820 97844 860
rect 97891 988 97900 1028
rect 97891 979 97940 988
rect 98092 988 98228 1028
rect 97708 197 97748 820
rect 97891 776 97931 979
rect 97995 944 98037 953
rect 97995 904 97996 944
rect 98036 904 98037 944
rect 97995 895 98037 904
rect 97804 736 97931 776
rect 97707 188 97749 197
rect 97707 148 97708 188
rect 97748 148 97749 188
rect 97707 139 97749 148
rect 97804 80 97844 736
rect 97996 80 98036 895
rect 98092 281 98132 988
rect 98284 944 98324 1324
rect 98420 1324 98516 1364
rect 98380 1315 98420 1324
rect 98476 1280 98516 1324
rect 98859 1280 98901 1289
rect 98476 1240 98708 1280
rect 98379 1196 98421 1205
rect 98379 1156 98380 1196
rect 98420 1156 98421 1196
rect 98379 1147 98421 1156
rect 98380 1112 98420 1147
rect 98668 1121 98708 1240
rect 98859 1240 98860 1280
rect 98900 1240 98901 1280
rect 98859 1231 98901 1240
rect 98763 1196 98805 1205
rect 98763 1156 98764 1196
rect 98804 1156 98805 1196
rect 98763 1147 98805 1156
rect 98572 1112 98612 1121
rect 98380 1061 98420 1072
rect 98476 1072 98572 1112
rect 98284 904 98420 944
rect 98187 860 98229 869
rect 98187 820 98188 860
rect 98228 820 98229 860
rect 98187 811 98229 820
rect 98091 272 98133 281
rect 98091 232 98092 272
rect 98132 232 98133 272
rect 98091 223 98133 232
rect 98188 80 98228 811
rect 98380 80 98420 904
rect 98476 365 98516 1072
rect 98572 1063 98612 1072
rect 98667 1112 98709 1121
rect 98667 1072 98668 1112
rect 98708 1072 98709 1112
rect 98667 1063 98709 1072
rect 98764 1112 98804 1147
rect 98764 1061 98804 1072
rect 98668 944 98708 953
rect 98572 904 98668 944
rect 98475 356 98517 365
rect 98475 316 98476 356
rect 98516 316 98517 356
rect 98475 307 98517 316
rect 98572 80 98612 904
rect 98668 895 98708 904
rect 98860 860 98900 1231
rect 98955 1196 98997 1205
rect 98955 1156 98956 1196
rect 98996 1156 98997 1196
rect 98955 1147 98997 1156
rect 98956 1112 98996 1147
rect 98956 1061 98996 1072
rect 99147 1112 99189 1121
rect 99147 1072 99148 1112
rect 99188 1072 99189 1112
rect 99147 1063 99189 1072
rect 99148 978 99188 1063
rect 99052 944 99092 953
rect 98764 820 98900 860
rect 98956 904 99052 944
rect 98764 80 98804 820
rect 98956 80 98996 904
rect 99052 895 99092 904
rect 95156 64 95176 80
rect 95096 0 95176 64
rect 95288 0 95368 80
rect 95480 0 95560 80
rect 95672 0 95752 80
rect 95864 0 95944 80
rect 96056 0 96136 80
rect 96248 0 96328 80
rect 96440 0 96520 80
rect 96632 0 96712 80
rect 96824 0 96904 80
rect 97016 0 97096 80
rect 97208 0 97288 80
rect 97400 0 97480 80
rect 97592 0 97672 80
rect 97784 0 97864 80
rect 97976 0 98056 80
rect 98168 0 98248 80
rect 98360 0 98440 80
rect 98552 0 98632 80
rect 98744 0 98824 80
rect 98936 0 99016 80
<< via2 >>
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 6220 6952 6260 6992
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 24556 6952 24596 6992
rect 28108 6952 28148 6992
rect 17164 6868 17204 6908
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 41068 6952 41108 6992
rect 41740 6952 41780 6992
rect 39052 6616 39092 6656
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 24556 5608 24596 5648
rect 41356 6868 41396 6908
rect 42028 6868 42068 6908
rect 41740 6532 41780 6572
rect 46732 6616 46772 6656
rect 47596 6616 47636 6656
rect 48460 6616 48500 6656
rect 44716 6532 44756 6572
rect 45772 6532 45812 6572
rect 46348 6532 46388 6572
rect 42028 6448 42068 6488
rect 44524 6448 44564 6488
rect 45868 6448 45908 6488
rect 46540 6532 46580 6572
rect 46636 6448 46676 6488
rect 41452 5608 41492 5648
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 18892 4516 18932 4556
rect 19468 4516 19508 4556
rect 20044 4516 20084 4556
rect 18508 4348 18548 4388
rect 6988 4264 7028 4304
rect 7564 4264 7604 4304
rect 7180 4096 7220 4136
rect 7564 4096 7604 4136
rect 18316 4096 18356 4136
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 4396 3592 4436 3632
rect 1612 3088 1652 3128
rect 2092 3424 2132 3464
rect 3724 3424 3764 3464
rect 4204 3424 4244 3464
rect 6412 3508 6452 3548
rect 4588 3424 4628 3464
rect 2668 3256 2708 3296
rect 1804 2416 1844 2456
rect 1036 1240 1076 1280
rect 844 1156 884 1196
rect 1228 1072 1268 1112
rect 1516 1912 1556 1952
rect 1420 1240 1460 1280
rect 2284 2584 2324 2624
rect 2092 2416 2132 2456
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 3148 2752 3188 2792
rect 2476 2416 2516 2456
rect 1516 1156 1556 1196
rect 1612 1072 1652 1112
rect 1804 1156 1844 1196
rect 1996 1072 2036 1112
rect 2860 2500 2900 2540
rect 3532 2584 3572 2624
rect 4972 3424 5012 3464
rect 5164 3424 5204 3464
rect 3244 2500 3284 2540
rect 3916 2584 3956 2624
rect 3628 2500 3668 2540
rect 4684 3172 4724 3212
rect 4876 3172 4916 3212
rect 4972 3004 5012 3044
rect 2188 1072 2228 1112
rect 2380 652 2420 692
rect 2572 1156 2612 1196
rect 2764 1072 2804 1112
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 2956 1156 2996 1196
rect 3148 1072 3188 1112
rect 3340 1156 3380 1196
rect 3532 1072 3572 1112
rect 3724 1240 3764 1280
rect 3916 1072 3956 1112
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 5932 3424 5972 3464
rect 5740 3004 5780 3044
rect 5356 2584 5396 2624
rect 5740 2584 5780 2624
rect 5548 2248 5588 2288
rect 4108 1240 4148 1280
rect 5068 1240 5108 1280
rect 4492 1156 4532 1196
rect 4300 1072 4340 1112
rect 4876 1156 4916 1196
rect 4684 1072 4724 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 4300 568 4340 608
rect 4684 316 4724 356
rect 5068 568 5108 608
rect 6700 3424 6740 3464
rect 6892 3424 6932 3464
rect 7084 3424 7124 3464
rect 6412 3088 6452 3128
rect 6316 3004 6356 3044
rect 6124 2584 6164 2624
rect 6796 3088 6836 3128
rect 6700 2920 6740 2960
rect 6604 2584 6644 2624
rect 6412 2416 6452 2456
rect 6412 1996 6452 2036
rect 6220 1324 6260 1364
rect 5260 1156 5300 1196
rect 6796 1996 6836 2036
rect 6796 1408 6836 1448
rect 6700 1240 6740 1280
rect 5644 1156 5684 1196
rect 6124 1156 6164 1196
rect 6412 1156 6452 1196
rect 5356 652 5396 692
rect 5836 484 5876 524
rect 6508 1072 6548 1112
rect 5932 232 5972 272
rect 7276 3508 7316 3548
rect 9196 3760 9236 3800
rect 15244 3760 15284 3800
rect 8428 3676 8468 3716
rect 7468 3424 7508 3464
rect 6988 2584 7028 2624
rect 7180 2584 7220 2624
rect 7084 2500 7124 2540
rect 6988 2080 7028 2120
rect 7276 1996 7316 2036
rect 6988 1156 7028 1196
rect 6412 904 6452 944
rect 6220 736 6260 776
rect 6220 484 6260 524
rect 6807 904 6847 944
rect 6508 316 6548 356
rect 6796 316 6836 356
rect 6604 148 6644 188
rect 7180 1156 7220 1196
rect 7372 1156 7412 1196
rect 7852 3424 7892 3464
rect 8236 3424 8276 3464
rect 7660 2920 7700 2960
rect 7564 1156 7604 1196
rect 7756 1072 7796 1112
rect 7276 904 7316 944
rect 7564 904 7604 944
rect 8044 2584 8084 2624
rect 8620 3424 8660 3464
rect 8428 3256 8468 3296
rect 7660 484 7700 524
rect 8140 1072 8180 1112
rect 8332 1156 8372 1196
rect 8524 1156 8564 1196
rect 8044 904 8084 944
rect 8332 904 8372 944
rect 7948 484 7988 524
rect 7852 232 7892 272
rect 9004 3424 9044 3464
rect 12076 3676 12116 3716
rect 12460 3676 12500 3716
rect 10156 3592 10196 3632
rect 10540 3592 10580 3632
rect 10924 3592 10964 3632
rect 11308 3592 11348 3632
rect 11692 3592 11732 3632
rect 9580 3508 9620 3548
rect 9964 3508 10004 3548
rect 8812 2752 8852 2792
rect 8908 1156 8948 1196
rect 8428 484 8468 524
rect 9388 3424 9428 3464
rect 9772 3424 9812 3464
rect 10156 3424 10196 3464
rect 11116 3424 11156 3464
rect 11500 3424 11540 3464
rect 11692 3424 11732 3464
rect 10732 3340 10772 3380
rect 10348 3256 10388 3296
rect 9196 2668 9236 2708
rect 9100 1240 9140 1280
rect 9292 1156 9332 1196
rect 9100 1072 9140 1112
rect 8812 904 8852 944
rect 9100 904 9140 944
rect 8716 484 8756 524
rect 8620 400 8660 440
rect 9676 1156 9716 1196
rect 9484 988 9524 1028
rect 9196 484 9236 524
rect 10060 1156 10100 1196
rect 9868 1072 9908 1112
rect 9580 904 9620 944
rect 9868 904 9908 944
rect 9484 820 9524 860
rect 9484 484 9524 524
rect 10444 1156 10484 1196
rect 10252 1072 10292 1112
rect 10828 1156 10868 1196
rect 10636 1072 10676 1112
rect 10348 904 10388 944
rect 9964 484 10004 524
rect 10636 904 10676 944
rect 10252 484 10292 524
rect 11692 3256 11732 3296
rect 11116 2248 11156 2288
rect 11212 1156 11252 1196
rect 10732 232 10772 272
rect 12076 3424 12116 3464
rect 16780 3676 16820 3716
rect 14476 3592 14516 3632
rect 15244 3592 15284 3632
rect 13228 3508 13268 3548
rect 13612 3508 13652 3548
rect 13996 3508 14036 3548
rect 14284 3508 14324 3548
rect 12268 3256 12308 3296
rect 11884 3172 11924 3212
rect 11692 2836 11732 2876
rect 12268 3088 12308 3128
rect 13036 3424 13076 3464
rect 12748 2584 12788 2624
rect 11596 1156 11636 1196
rect 11500 1072 11540 1112
rect 11980 1156 12020 1196
rect 11116 904 11156 944
rect 11404 904 11444 944
rect 11020 652 11060 692
rect 11020 400 11060 440
rect 11020 232 11060 272
rect 11500 148 11540 188
rect 12172 2080 12212 2120
rect 12364 1156 12404 1196
rect 12172 1072 12212 1112
rect 11692 820 11732 860
rect 13036 1576 13076 1616
rect 12652 1156 12692 1196
rect 12556 1072 12596 1112
rect 12268 904 12308 944
rect 11884 484 11924 524
rect 11788 400 11828 440
rect 11788 148 11828 188
rect 12556 904 12596 944
rect 12172 484 12212 524
rect 13036 1156 13076 1196
rect 12940 1072 12980 1112
rect 13132 1072 13172 1112
rect 13804 2920 13844 2960
rect 13420 2416 13460 2456
rect 13324 1156 13364 1196
rect 13516 1072 13556 1112
rect 13036 904 13076 944
rect 12652 484 12692 524
rect 13324 904 13364 944
rect 12940 484 12980 524
rect 14668 3508 14708 3548
rect 15052 3508 15092 3548
rect 14284 2668 14324 2708
rect 13804 2416 13844 2456
rect 13420 484 13460 524
rect 13900 1072 13940 1112
rect 14092 1156 14132 1196
rect 13804 904 13844 944
rect 14092 904 14132 944
rect 13708 736 13748 776
rect 13708 484 13748 524
rect 14476 2668 14516 2708
rect 15436 3508 15476 3548
rect 15820 3508 15860 3548
rect 16204 3508 16244 3548
rect 16588 3508 16628 3548
rect 16012 3424 16052 3464
rect 15820 3256 15860 3296
rect 14860 2752 14900 2792
rect 14284 2332 14324 2372
rect 14284 1324 14324 1364
rect 14284 1072 14324 1112
rect 14668 1072 14708 1112
rect 14860 1156 14900 1196
rect 15052 1156 15092 1196
rect 14572 904 14612 944
rect 14860 904 14900 944
rect 14380 820 14420 860
rect 14572 736 14612 776
rect 14476 652 14516 692
rect 14572 232 14612 272
rect 15244 1240 15284 1280
rect 15436 1156 15476 1196
rect 14956 232 14996 272
rect 15244 652 15284 692
rect 15820 1156 15860 1196
rect 15628 988 15668 1028
rect 16972 3508 17012 3548
rect 17356 3508 17396 3548
rect 17932 3508 17972 3548
rect 17164 3424 17204 3464
rect 17548 3424 17588 3464
rect 17740 3424 17780 3464
rect 18412 3928 18452 3968
rect 18508 3844 18548 3884
rect 19084 4348 19124 4388
rect 19756 4348 19796 4388
rect 18988 4012 19028 4052
rect 19180 4012 19220 4052
rect 18892 3928 18932 3968
rect 19084 3928 19124 3968
rect 18796 3760 18836 3800
rect 16780 3256 16820 3296
rect 18124 3424 18164 3464
rect 18508 3424 18548 3464
rect 18700 3424 18740 3464
rect 19084 3760 19124 3800
rect 19756 4096 19796 4136
rect 19948 4096 19988 4136
rect 16396 2836 16436 2876
rect 16204 1156 16244 1196
rect 16012 1072 16052 1112
rect 15724 904 15764 944
rect 16012 904 16052 944
rect 15148 232 15188 272
rect 15340 232 15380 272
rect 15628 232 15668 272
rect 16396 1240 16436 1280
rect 16396 988 16436 1028
rect 16588 1156 16628 1196
rect 16780 1240 16820 1280
rect 16972 1156 17012 1196
rect 16108 232 16148 272
rect 16396 232 16436 272
rect 16684 820 16724 860
rect 16684 232 16724 272
rect 17356 1156 17396 1196
rect 17164 1072 17204 1112
rect 16876 904 16916 944
rect 17164 904 17204 944
rect 17932 3172 17972 3212
rect 18316 3172 18356 3212
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 17644 1072 17684 1112
rect 17836 1072 17876 1112
rect 18028 1072 18068 1112
rect 17932 988 17972 1028
rect 17548 904 17588 944
rect 17260 484 17300 524
rect 17740 904 17780 944
rect 18988 3088 19028 3128
rect 18988 2752 19028 2792
rect 19660 3928 19700 3968
rect 19948 3928 19988 3968
rect 22348 4180 22388 4220
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 38668 4516 38708 4556
rect 37324 4348 37364 4388
rect 38188 4348 38228 4388
rect 38956 4432 38996 4472
rect 25900 4264 25940 4304
rect 28012 4264 28052 4304
rect 24460 4180 24500 4220
rect 25132 4180 25172 4220
rect 22444 4012 22484 4052
rect 24268 4012 24308 4052
rect 20236 3928 20276 3968
rect 24364 3928 24404 3968
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 21100 3760 21140 3800
rect 19372 3508 19412 3548
rect 20716 3508 20756 3548
rect 19948 3424 19988 3464
rect 20149 3449 20189 3464
rect 20149 3424 20189 3449
rect 19372 3172 19412 3212
rect 20044 2836 20084 2876
rect 19852 2752 19892 2792
rect 19468 2584 19508 2624
rect 19660 2584 19700 2624
rect 20908 3424 20948 3464
rect 21676 3676 21716 3716
rect 21388 3592 21428 3632
rect 20716 2668 20756 2708
rect 18892 1576 18932 1616
rect 18316 1156 18356 1196
rect 18508 1072 18548 1112
rect 18028 904 18068 944
rect 18316 904 18356 944
rect 17932 820 17972 860
rect 17740 736 17780 776
rect 17548 484 17588 524
rect 18892 1072 18932 1112
rect 18700 988 18740 1028
rect 18796 904 18836 944
rect 18700 820 18740 860
rect 18412 484 18452 524
rect 19084 1240 19124 1280
rect 20236 2584 20276 2624
rect 20428 2584 20468 2624
rect 19372 2248 19412 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 19372 1912 19412 1952
rect 19564 1912 19604 1952
rect 19276 1156 19316 1196
rect 19180 1072 19220 1112
rect 19084 904 19124 944
rect 18700 484 18740 524
rect 18796 400 18836 440
rect 19468 1408 19508 1448
rect 19468 1240 19508 1280
rect 19852 1240 19892 1280
rect 19660 1072 19700 1112
rect 21292 3424 21332 3464
rect 23116 3592 23156 3632
rect 21676 3424 21716 3464
rect 22060 3424 22100 3464
rect 21100 3088 21140 3128
rect 21868 2584 21908 2624
rect 22540 3424 22580 3464
rect 22348 3340 22388 3380
rect 20044 1912 20084 1952
rect 19948 1156 19988 1196
rect 20236 1156 20276 1196
rect 20044 1072 20084 1112
rect 19852 988 19892 1028
rect 19564 904 19604 944
rect 19948 904 19988 944
rect 20236 904 20276 944
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 19180 484 19220 524
rect 19468 484 19508 524
rect 19948 484 19988 524
rect 19852 64 19892 104
rect 20044 64 20084 104
rect 20428 1492 20468 1532
rect 20428 1072 20468 1112
rect 20812 1072 20852 1112
rect 20620 988 20660 1028
rect 21004 1156 21044 1196
rect 21196 1156 21236 1196
rect 20716 904 20756 944
rect 21004 904 21044 944
rect 20620 484 20660 524
rect 21580 1156 21620 1196
rect 21100 484 21140 524
rect 22924 3424 22964 3464
rect 22732 2920 22772 2960
rect 21964 1156 22004 1196
rect 21388 820 21428 860
rect 21388 484 21428 524
rect 22156 1072 22196 1112
rect 22348 1072 22388 1112
rect 21484 316 21524 356
rect 21772 316 21812 356
rect 21676 148 21716 188
rect 22252 904 22292 944
rect 21868 232 21908 272
rect 22540 1156 22580 1196
rect 22732 1072 22772 1112
rect 22540 904 22580 944
rect 22156 232 22196 272
rect 23596 3424 23636 3464
rect 23788 3424 23828 3464
rect 24172 3256 24212 3296
rect 23596 3172 23636 3212
rect 23116 2668 23156 2708
rect 23404 2584 23444 2624
rect 23116 1072 23156 1112
rect 22924 988 22964 1028
rect 23020 904 23060 944
rect 23980 3172 24020 3212
rect 24364 3172 24404 3212
rect 27916 4096 27956 4136
rect 25036 4012 25076 4052
rect 26092 4012 26132 4052
rect 24652 3172 24692 3212
rect 24556 3004 24596 3044
rect 24556 2836 24596 2876
rect 23692 1492 23732 1532
rect 23308 1156 23348 1196
rect 23500 1072 23540 1112
rect 23308 904 23348 944
rect 23788 1072 23828 1112
rect 23884 988 23924 1028
rect 22636 484 22676 524
rect 22924 484 22964 524
rect 23788 904 23828 944
rect 23404 232 23444 272
rect 23884 484 23924 524
rect 23692 232 23732 272
rect 24268 1072 24308 1112
rect 24071 904 24111 944
rect 24172 904 24212 944
rect 23980 400 24020 440
rect 24460 1156 24500 1196
rect 24460 904 24500 944
rect 24940 3928 24980 3968
rect 25324 3424 25364 3464
rect 25516 3424 25556 3464
rect 24844 1912 24884 1952
rect 24748 1660 24788 1700
rect 24652 1156 24692 1196
rect 25132 1660 25172 1700
rect 25036 1156 25076 1196
rect 24844 1072 24884 1112
rect 24940 904 24980 944
rect 25228 904 25268 944
rect 27340 3760 27380 3800
rect 26956 3508 26996 3548
rect 25900 3424 25940 3464
rect 25708 2416 25748 2456
rect 25516 1408 25556 1448
rect 25708 1240 25748 1280
rect 25516 1072 25556 1112
rect 25708 904 25748 944
rect 25612 484 25652 524
rect 26284 3424 26324 3464
rect 26764 3424 26804 3464
rect 26092 3088 26132 3128
rect 26092 2164 26132 2204
rect 25900 1240 25940 1280
rect 26092 1828 26132 1868
rect 26092 1324 26132 1364
rect 25996 1072 26036 1112
rect 25900 988 25940 1028
rect 26092 988 26132 1028
rect 25996 652 26036 692
rect 25996 484 26036 524
rect 26572 2584 26612 2624
rect 27148 3424 27188 3464
rect 27628 3676 27668 3716
rect 27820 3424 27860 3464
rect 26956 3004 26996 3044
rect 28108 2584 28148 2624
rect 26476 1072 26516 1112
rect 26380 904 26420 944
rect 26284 736 26324 776
rect 26380 652 26420 692
rect 26668 1156 26708 1196
rect 26860 1072 26900 1112
rect 26668 904 26708 944
rect 26764 652 26804 692
rect 27244 1072 27284 1112
rect 27148 904 27188 944
rect 27148 652 27188 692
rect 27052 568 27092 608
rect 27052 232 27092 272
rect 27436 1240 27476 1280
rect 27628 1072 27668 1112
rect 27436 904 27476 944
rect 27532 652 27572 692
rect 28012 1072 28052 1112
rect 27916 904 27956 944
rect 27820 820 27860 860
rect 27916 652 27956 692
rect 27820 484 27860 524
rect 28204 1156 28244 1196
rect 28396 3508 28436 3548
rect 28396 3340 28436 3380
rect 28588 3340 28628 3380
rect 28300 1072 28340 1112
rect 28204 904 28244 944
rect 28300 652 28340 692
rect 28972 3340 29012 3380
rect 28780 2920 28820 2960
rect 28780 1072 28820 1112
rect 28684 904 28724 944
rect 28684 652 28724 692
rect 28588 568 28628 608
rect 28780 568 28820 608
rect 28780 148 28820 188
rect 29836 3424 29876 3464
rect 29356 3340 29396 3380
rect 29644 3340 29684 3380
rect 29164 2668 29204 2708
rect 28972 1492 29012 1532
rect 29164 1156 29204 1196
rect 28972 1072 29012 1112
rect 28972 904 29012 944
rect 29068 484 29108 524
rect 30220 3424 30260 3464
rect 30028 3340 30068 3380
rect 30412 3340 30452 3380
rect 29548 2584 29588 2624
rect 29740 2584 29780 2624
rect 29548 1156 29588 1196
rect 29452 652 29492 692
rect 29356 568 29396 608
rect 29452 484 29492 524
rect 29356 148 29396 188
rect 29932 1156 29972 1196
rect 29740 1072 29780 1112
rect 29836 904 29876 944
rect 29836 652 29876 692
rect 30316 1156 30356 1196
rect 30124 1072 30164 1112
rect 30124 904 30164 944
rect 30220 652 30260 692
rect 30508 904 30548 944
rect 30700 2836 30740 2876
rect 30700 2584 30740 2624
rect 30892 2584 30932 2624
rect 30700 1324 30740 1364
rect 31468 3424 31508 3464
rect 31180 2164 31220 2204
rect 31180 1660 31220 1700
rect 30700 1072 30740 1112
rect 30892 1072 30932 1112
rect 31084 1072 31124 1112
rect 30604 652 30644 692
rect 30988 904 31028 944
rect 30988 568 31028 608
rect 31660 3424 31700 3464
rect 32236 4096 32276 4136
rect 32812 4096 32852 4136
rect 32236 3928 32276 3968
rect 32524 3928 32564 3968
rect 32140 3844 32180 3884
rect 32236 3592 32276 3632
rect 32044 3424 32084 3464
rect 32428 3424 32468 3464
rect 31564 3088 31604 3128
rect 31756 3172 31796 3212
rect 31660 2584 31700 2624
rect 31564 2080 31604 2120
rect 31948 1912 31988 1952
rect 31468 1576 31508 1616
rect 31468 1072 31508 1112
rect 31372 904 31412 944
rect 31276 652 31316 692
rect 31660 1240 31700 1280
rect 31660 1072 31700 1112
rect 31852 1324 31892 1364
rect 31852 1156 31892 1196
rect 32140 1828 32180 1868
rect 32140 1240 32180 1280
rect 32620 3004 32660 3044
rect 37228 4096 37268 4136
rect 37708 4180 37748 4220
rect 37804 4096 37844 4136
rect 37228 3928 37268 3968
rect 32908 3844 32948 3884
rect 33004 3760 33044 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 35692 3760 35732 3800
rect 33388 3676 33428 3716
rect 33004 3592 33044 3632
rect 32812 3424 32852 3464
rect 33196 3424 33236 3464
rect 33580 3424 33620 3464
rect 32716 1912 32756 1952
rect 32620 1744 32660 1784
rect 32524 1408 32564 1448
rect 32044 1072 32084 1112
rect 31948 652 31988 692
rect 32044 400 32084 440
rect 32236 1156 32276 1196
rect 32428 1072 32468 1112
rect 32236 904 32276 944
rect 32620 1240 32660 1280
rect 32812 1072 32852 1112
rect 32716 904 32756 944
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 33772 2584 33812 2624
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 33196 1072 33236 1112
rect 33580 1072 33620 1112
rect 33388 988 33428 1028
rect 32332 484 32372 524
rect 32524 400 32564 440
rect 32908 652 32948 692
rect 32908 484 32948 524
rect 33100 568 33140 608
rect 33004 232 33044 272
rect 33292 904 33332 944
rect 33196 484 33236 524
rect 33484 652 33524 692
rect 34156 3508 34196 3548
rect 33964 3424 34004 3464
rect 34348 3424 34388 3464
rect 34444 3172 34484 3212
rect 34732 3424 34772 3464
rect 34540 2920 34580 2960
rect 33868 1240 33908 1280
rect 33964 1072 34004 1112
rect 35116 3424 35156 3464
rect 35500 3424 35540 3464
rect 37708 3928 37748 3968
rect 35884 3424 35924 3464
rect 36268 3424 36308 3464
rect 36076 3340 36116 3380
rect 35308 3004 35348 3044
rect 34924 2668 34964 2708
rect 34828 2416 34868 2456
rect 35308 2416 35348 2456
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 34924 1408 34964 1448
rect 35308 1408 35348 1448
rect 34444 1240 34484 1280
rect 34156 1156 34196 1196
rect 34252 1072 34292 1112
rect 33772 820 33812 860
rect 33676 484 33716 524
rect 33580 400 33620 440
rect 34156 568 34196 608
rect 33868 484 33908 524
rect 34732 1156 34772 1196
rect 34540 1072 34580 1112
rect 35116 1156 35156 1196
rect 35500 1156 35540 1196
rect 35404 1072 35444 1112
rect 34636 904 34676 944
rect 35212 904 35252 944
rect 35404 904 35444 944
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 34060 400 34100 440
rect 34252 400 34292 440
rect 34636 568 34676 608
rect 34444 484 34484 524
rect 34732 484 34772 524
rect 34828 400 34868 440
rect 35020 400 35060 440
rect 34732 148 34772 188
rect 35116 148 35156 188
rect 35404 400 35444 440
rect 35692 2164 35732 2204
rect 35692 1660 35732 1700
rect 36076 3004 36116 3044
rect 35980 1492 36020 1532
rect 36652 3424 36692 3464
rect 36844 3424 36884 3464
rect 37516 3424 37556 3464
rect 37708 3424 37748 3464
rect 38092 4012 38132 4052
rect 37996 3760 38036 3800
rect 38476 4180 38516 4220
rect 38380 4096 38420 4136
rect 38956 4012 38996 4052
rect 38380 3928 38420 3968
rect 38284 3676 38324 3716
rect 41452 5440 41492 5480
rect 41548 5188 41588 5228
rect 41548 5020 41588 5060
rect 41356 4936 41396 4976
rect 41260 4348 41300 4388
rect 41452 4264 41492 4304
rect 47884 6448 47924 6488
rect 49036 6616 49076 6656
rect 48556 6448 48596 6488
rect 48748 6448 48788 6488
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 49420 6448 49460 6488
rect 46828 6280 46868 6320
rect 41836 5440 41876 5480
rect 41740 5020 41780 5060
rect 41644 4936 41684 4976
rect 41452 4096 41492 4136
rect 41740 4348 41780 4388
rect 41260 3928 41300 3968
rect 41644 3928 41684 3968
rect 41740 3676 41780 3716
rect 38380 3592 38420 3632
rect 38572 3592 38612 3632
rect 40972 3592 41012 3632
rect 36460 2836 36500 2876
rect 36460 2248 36500 2288
rect 36748 1492 36788 1532
rect 36364 1408 36404 1448
rect 35884 1156 35924 1196
rect 36268 1156 36308 1196
rect 35980 1072 36020 1112
rect 35692 820 35732 860
rect 35980 904 36020 944
rect 35788 484 35828 524
rect 35596 148 35636 188
rect 36364 1072 36404 1112
rect 36172 904 36212 944
rect 36652 1072 36692 1112
rect 37132 1408 37172 1448
rect 36844 1072 36884 1112
rect 37036 1072 37076 1112
rect 36460 820 36500 860
rect 36076 316 36116 356
rect 36364 484 36404 524
rect 36556 484 36596 524
rect 36844 820 36884 860
rect 38476 3424 38516 3464
rect 38380 3340 38420 3380
rect 37804 2584 37844 2624
rect 37612 2332 37652 2372
rect 37612 1912 37652 1952
rect 37804 1576 37844 1616
rect 37324 1072 37364 1112
rect 37516 1072 37556 1112
rect 36940 400 36980 440
rect 37132 484 37172 524
rect 37420 904 37460 944
rect 37996 2836 38036 2876
rect 37900 1072 37940 1112
rect 37516 400 37556 440
rect 37900 904 37940 944
rect 40492 3508 40532 3548
rect 41356 3508 41396 3548
rect 38860 3424 38900 3464
rect 39244 3424 39284 3464
rect 39052 3340 39092 3380
rect 38284 2836 38324 2876
rect 38188 2500 38228 2540
rect 38092 2164 38132 2204
rect 38092 1324 38132 1364
rect 38572 2584 38612 2624
rect 38764 2584 38804 2624
rect 38380 2080 38420 2120
rect 38284 1072 38324 1112
rect 37804 484 37844 524
rect 38188 904 38228 944
rect 38476 1156 38516 1196
rect 38668 1072 38708 1112
rect 38284 484 38324 524
rect 38668 904 38708 944
rect 39628 3424 39668 3464
rect 39436 3256 39476 3296
rect 40012 3424 40052 3464
rect 40300 3424 40340 3464
rect 39436 3088 39476 3128
rect 39820 3172 39860 3212
rect 40780 3424 40820 3464
rect 40492 3256 40532 3296
rect 40204 2584 40244 2624
rect 39052 1744 39092 1784
rect 38860 1156 38900 1196
rect 39052 1072 39092 1112
rect 38572 484 38612 524
rect 38956 904 38996 944
rect 39244 1156 39284 1196
rect 39436 1072 39476 1112
rect 39052 484 39092 524
rect 39436 904 39476 944
rect 39628 1240 39668 1280
rect 39820 1072 39860 1112
rect 39340 400 39380 440
rect 39724 904 39764 944
rect 41164 3424 41204 3464
rect 40972 2920 41012 2960
rect 40972 2752 41012 2792
rect 40012 1156 40052 1196
rect 40204 1072 40244 1112
rect 39820 400 39860 440
rect 40204 904 40244 944
rect 40396 1156 40436 1196
rect 40588 1072 40628 1112
rect 40108 484 40148 524
rect 40492 904 40532 944
rect 40972 1156 41012 1196
rect 40780 1072 40820 1112
rect 40588 484 40628 524
rect 40972 904 41012 944
rect 41644 3424 41684 3464
rect 42124 5440 42164 5480
rect 42028 5020 42068 5060
rect 42700 5020 42740 5060
rect 42124 4936 42164 4976
rect 41932 4348 41972 4388
rect 42124 4264 42164 4304
rect 42604 4264 42644 4304
rect 42028 4180 42068 4220
rect 41932 4096 41972 4136
rect 43948 4516 43988 4556
rect 42796 4348 42836 4388
rect 42508 4012 42548 4052
rect 42028 3928 42068 3968
rect 42316 3928 42356 3968
rect 41932 3424 41972 3464
rect 42124 3340 42164 3380
rect 41836 3172 41876 3212
rect 42028 3172 42068 3212
rect 42124 3088 42164 3128
rect 41836 2920 41876 2960
rect 41356 2668 41396 2708
rect 41644 2668 41684 2708
rect 42028 2668 42068 2708
rect 41836 2584 41876 2624
rect 42220 2584 42260 2624
rect 41740 2500 41780 2540
rect 42028 2416 42068 2456
rect 41164 1072 41204 1112
rect 41356 1072 41396 1112
rect 40876 484 40916 524
rect 41260 904 41300 944
rect 42316 2500 42356 2540
rect 43180 4180 43220 4220
rect 43084 4012 43124 4052
rect 42892 3928 42932 3968
rect 42604 3172 42644 3212
rect 42412 2416 42452 2456
rect 42028 1240 42068 1280
rect 41548 1072 41588 1112
rect 41740 1072 41780 1112
rect 42124 1156 42164 1196
rect 42028 1072 42068 1112
rect 41943 988 41983 1028
rect 41356 484 41396 524
rect 41740 904 41780 944
rect 42028 904 42068 944
rect 42316 1240 42356 1280
rect 42508 1156 42548 1196
rect 42316 1072 42356 1112
rect 41644 400 41684 440
rect 41932 568 41972 608
rect 42124 400 42164 440
rect 42508 904 42548 944
rect 42796 2668 42836 2708
rect 42988 2584 43028 2624
rect 42892 1996 42932 2036
rect 43180 3172 43220 3212
rect 43180 2248 43220 2288
rect 43564 3760 43604 3800
rect 43468 1996 43508 2036
rect 43372 1324 43412 1364
rect 42700 1156 42740 1196
rect 42892 1072 42932 1112
rect 42412 400 42452 440
rect 42796 904 42836 944
rect 43372 1156 43412 1196
rect 43084 1072 43124 1112
rect 43276 1072 43316 1112
rect 42892 400 42932 440
rect 43276 904 43316 944
rect 43180 316 43220 356
rect 43948 3508 43988 3548
rect 44332 5608 44372 5648
rect 44524 5608 44564 5648
rect 45004 5608 45044 5648
rect 44620 5524 44660 5564
rect 44332 5104 44372 5144
rect 44236 4180 44276 4220
rect 44620 5020 44660 5060
rect 44332 4096 44372 4136
rect 44908 5524 44948 5564
rect 44812 5104 44852 5144
rect 45004 5104 45044 5144
rect 45868 5104 45908 5144
rect 45964 4936 46004 4976
rect 45868 4852 45908 4892
rect 46348 5524 46388 5564
rect 46540 5524 46580 5564
rect 47596 5524 47636 5564
rect 46156 5104 46196 5144
rect 46636 5104 46676 5144
rect 48076 5104 48116 5144
rect 46636 4936 46676 4976
rect 46252 4852 46292 4892
rect 45100 4180 45140 4220
rect 44428 4012 44468 4052
rect 45004 4012 45044 4052
rect 44236 3676 44276 3716
rect 44044 2836 44084 2876
rect 43852 1912 43892 1952
rect 43564 1072 43604 1112
rect 43756 1072 43796 1112
rect 43660 484 43700 524
rect 43660 316 43700 356
rect 44236 2416 44276 2456
rect 44620 3760 44660 3800
rect 44620 3592 44660 3632
rect 44428 3508 44468 3548
rect 44620 3088 44660 3128
rect 44332 1408 44372 1448
rect 44140 1072 44180 1112
rect 44140 652 44180 692
rect 43948 568 43988 608
rect 44044 484 44084 524
rect 44343 1156 44383 1196
rect 44428 1072 44468 1112
rect 44332 736 44372 776
rect 44428 652 44468 692
rect 44332 400 44372 440
rect 44524 232 44564 272
rect 44812 3508 44852 3548
rect 45196 3508 45236 3548
rect 45580 3508 45620 3548
rect 45388 3424 45428 3464
rect 45004 2836 45044 2876
rect 45484 2164 45524 2204
rect 45772 3004 45812 3044
rect 46060 4096 46100 4136
rect 46060 3760 46100 3800
rect 46252 4180 46292 4220
rect 46348 4096 46388 4136
rect 45964 3508 46004 3548
rect 46156 3004 46196 3044
rect 45772 2080 45812 2120
rect 44908 1072 44948 1112
rect 44812 652 44852 692
rect 44716 484 44756 524
rect 44812 232 44852 272
rect 45100 1156 45140 1196
rect 45292 1072 45332 1112
rect 45100 736 45140 776
rect 45196 652 45236 692
rect 45292 568 45332 608
rect 45676 1072 45716 1112
rect 45484 904 45524 944
rect 45580 652 45620 692
rect 45484 568 45524 608
rect 45868 1324 45908 1364
rect 45964 1156 46004 1196
rect 46060 1072 46100 1112
rect 45868 988 45908 1028
rect 45964 904 46004 944
rect 45964 652 46004 692
rect 46348 3508 46388 3548
rect 47788 4264 47828 4304
rect 46636 4180 46676 4220
rect 48172 4936 48212 4976
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 56428 6280 56468 6320
rect 49516 5608 49556 5648
rect 48844 5104 48884 5144
rect 49324 5104 49364 5144
rect 48748 4936 48788 4976
rect 48268 4852 48308 4892
rect 49036 4936 49076 4976
rect 48556 4768 48596 4808
rect 48844 4768 48884 4808
rect 48076 4348 48116 4388
rect 48172 4264 48212 4304
rect 47788 3928 47828 3968
rect 47596 3676 47636 3716
rect 47212 3508 47252 3548
rect 46444 3424 46484 3464
rect 47020 3424 47060 3464
rect 46828 3256 46868 3296
rect 46540 2584 46580 2624
rect 46252 1912 46292 1952
rect 46252 1156 46292 1196
rect 46444 1072 46484 1112
rect 46252 904 46292 944
rect 46348 652 46388 692
rect 46636 1156 46676 1196
rect 46828 1072 46868 1112
rect 46636 988 46676 1028
rect 46732 904 46772 944
rect 46732 652 46772 692
rect 47404 3424 47444 3464
rect 47788 3424 47828 3464
rect 47212 2752 47252 2792
rect 47020 1072 47060 1112
rect 47212 988 47252 1028
rect 47020 904 47060 944
rect 47116 652 47156 692
rect 47596 988 47636 1028
rect 47500 904 47540 944
rect 47404 820 47444 860
rect 47500 652 47540 692
rect 48076 3340 48116 3380
rect 48076 2836 48116 2876
rect 47788 2752 47828 2792
rect 48076 2668 48116 2708
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 49612 5020 49652 5060
rect 49324 4768 49364 4808
rect 48652 4264 48692 4304
rect 49036 4264 49076 4304
rect 48364 4096 48404 4136
rect 48556 4096 48596 4136
rect 48844 4180 48884 4220
rect 48940 4096 48980 4136
rect 48748 4012 48788 4052
rect 48268 3508 48308 3548
rect 48268 2752 48308 2792
rect 49132 3592 49172 3632
rect 48748 3508 48788 3548
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 48844 2836 48884 2876
rect 48652 2752 48692 2792
rect 48364 2668 48404 2708
rect 48460 2584 48500 2624
rect 48940 2752 48980 2792
rect 47788 1072 47828 1112
rect 47980 988 48020 1028
rect 47788 904 47828 944
rect 47884 652 47924 692
rect 49132 3172 49172 3212
rect 49132 2752 49172 2792
rect 49324 2584 49364 2624
rect 50380 4936 50420 4976
rect 51244 5272 51284 5312
rect 50668 5104 50708 5144
rect 50860 5020 50900 5060
rect 50476 4852 50516 4892
rect 49612 4180 49652 4220
rect 50380 4684 50420 4724
rect 50188 4516 50228 4556
rect 50188 4096 50228 4136
rect 50668 4684 50708 4724
rect 50668 4348 50708 4388
rect 51532 4936 51572 4976
rect 51244 4768 51284 4808
rect 51532 4768 51572 4808
rect 50572 4096 50612 4136
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 50092 3424 50132 3464
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 48167 1156 48207 1196
rect 48268 1156 48308 1196
rect 48364 988 48404 1028
rect 48268 904 48308 944
rect 48268 652 48308 692
rect 48556 1240 48596 1280
rect 48748 1156 48788 1196
rect 48748 988 48788 1028
rect 48556 904 48596 944
rect 48652 652 48692 692
rect 49132 1156 49172 1196
rect 48940 1072 48980 1112
rect 49036 652 49076 692
rect 49132 148 49172 188
rect 49516 1240 49556 1280
rect 49324 1156 49364 1196
rect 49420 484 49460 524
rect 49420 148 49460 188
rect 49804 1324 49844 1364
rect 49708 1156 49748 1196
rect 49804 988 49844 1028
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 50284 3340 50324 3380
rect 50668 3424 50708 3464
rect 50764 3256 50804 3296
rect 50380 3004 50420 3044
rect 50284 1576 50324 1616
rect 50572 3004 50612 3044
rect 50668 1576 50708 1616
rect 50572 1240 50612 1280
rect 50380 1156 50420 1196
rect 50284 736 50324 776
rect 49804 484 49844 524
rect 50476 904 50516 944
rect 50956 4096 50996 4136
rect 51436 4348 51476 4388
rect 51916 5524 51956 5564
rect 52012 5020 52052 5060
rect 52780 5524 52820 5564
rect 52588 5272 52628 5312
rect 52300 5020 52340 5060
rect 52204 4936 52244 4976
rect 51820 4516 51860 4556
rect 51532 4264 51572 4304
rect 51436 4096 51476 4136
rect 51244 3928 51284 3968
rect 51148 3508 51188 3548
rect 52684 5020 52724 5060
rect 52396 4936 52436 4976
rect 52012 3424 52052 3464
rect 52012 3172 52052 3212
rect 51820 2248 51860 2288
rect 51052 1996 51092 2036
rect 51052 1324 51092 1364
rect 50956 1240 50996 1280
rect 51436 1996 51476 2036
rect 51244 1912 51284 1952
rect 52204 4348 52244 4388
rect 52588 4348 52628 4388
rect 53740 5608 53780 5648
rect 53740 5272 53780 5312
rect 52972 4936 53012 4976
rect 53548 4936 53588 4976
rect 52876 4852 52916 4892
rect 53836 4852 53876 4892
rect 53452 4768 53492 4808
rect 53740 4768 53780 4808
rect 52204 4180 52244 4220
rect 52780 4096 52820 4136
rect 52972 4264 53012 4304
rect 53356 4264 53396 4304
rect 53356 4096 53396 4136
rect 52780 3508 52820 3548
rect 52300 2248 52340 2288
rect 51724 1912 51764 1952
rect 51916 1912 51956 1952
rect 52108 1912 52148 1952
rect 51436 1828 51476 1868
rect 51148 1072 51188 1112
rect 50956 904 50996 944
rect 50860 736 50900 776
rect 51436 1072 51476 1112
rect 52204 1240 52244 1280
rect 52204 1072 52244 1112
rect 52108 904 52148 944
rect 52876 2248 52916 2288
rect 53836 4600 53876 4640
rect 53644 4264 53684 4304
rect 53836 4096 53876 4136
rect 53452 3760 53492 3800
rect 53260 3508 53300 3548
rect 53356 3172 53396 3212
rect 54508 5608 54548 5648
rect 54316 4936 54356 4976
rect 55084 5272 55124 5312
rect 54412 4852 54452 4892
rect 53932 3340 53972 3380
rect 54220 3172 54260 3212
rect 53356 2248 53396 2288
rect 52972 1912 53012 1952
rect 53164 1912 53204 1952
rect 52588 1240 52628 1280
rect 52684 1072 52724 1112
rect 52588 904 52628 944
rect 52492 736 52532 776
rect 54028 1660 54068 1700
rect 53740 1576 53780 1616
rect 53548 1072 53588 1112
rect 53452 904 53492 944
rect 53548 484 53588 524
rect 53548 148 53588 188
rect 53932 904 53972 944
rect 53836 484 53876 524
rect 54124 1576 54164 1616
rect 54508 3004 54548 3044
rect 54316 2248 54356 2288
rect 54508 1660 54548 1700
rect 54412 1408 54452 1448
rect 54892 4768 54932 4808
rect 54796 4600 54836 4640
rect 54892 4180 54932 4220
rect 54796 4096 54836 4136
rect 54700 2248 54740 2288
rect 54220 1324 54260 1364
rect 54124 1072 54164 1112
rect 54508 1072 54548 1112
rect 54412 316 54452 356
rect 55372 5104 55412 5144
rect 55180 4852 55220 4892
rect 55372 4600 55412 4640
rect 55276 4516 55316 4556
rect 55180 4096 55220 4136
rect 55564 5272 55604 5312
rect 56332 5608 56372 5648
rect 55660 4516 55700 4556
rect 54892 3844 54932 3884
rect 55084 3760 55124 3800
rect 54988 3172 55028 3212
rect 55372 3760 55412 3800
rect 55660 3760 55700 3800
rect 55564 3676 55604 3716
rect 55372 3004 55412 3044
rect 55180 2920 55220 2960
rect 54892 2613 54932 2616
rect 54892 2576 54932 2613
rect 54892 484 54932 524
rect 55084 1408 55124 1448
rect 55084 1072 55124 1112
rect 55276 2766 55316 2792
rect 55276 2752 55316 2766
rect 55564 2752 55604 2792
rect 55372 2584 55412 2624
rect 55276 2248 55316 2288
rect 55372 1744 55412 1784
rect 55276 1492 55316 1532
rect 55564 1660 55604 1700
rect 55372 1324 55412 1364
rect 55756 2752 55796 2792
rect 55756 2584 55796 2624
rect 56812 5608 56852 5648
rect 56428 5188 56468 5228
rect 55948 4768 55988 4808
rect 55852 1660 55892 1700
rect 55756 1324 55796 1364
rect 55660 1240 55700 1280
rect 55564 1072 55604 1112
rect 55564 736 55604 776
rect 55468 316 55508 356
rect 56428 4936 56468 4976
rect 56332 4768 56372 4808
rect 58060 5272 58100 5312
rect 56140 3424 56180 3464
rect 56044 2752 56084 2792
rect 56236 2584 56276 2624
rect 55948 1072 55988 1112
rect 55852 484 55892 524
rect 56236 1660 56276 1700
rect 56140 1240 56180 1280
rect 56044 736 56084 776
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 58156 5020 58196 5060
rect 57100 4096 57140 4136
rect 56620 3760 56660 3800
rect 56620 3424 56660 3464
rect 58060 4768 58100 4808
rect 57964 4516 58004 4556
rect 57676 3592 57716 3632
rect 57868 3592 57908 3632
rect 57100 3424 57140 3464
rect 56908 3340 56948 3380
rect 56620 3256 56660 3296
rect 56332 1324 56372 1364
rect 56428 1156 56468 1196
rect 56332 736 56372 776
rect 56332 484 56372 524
rect 56716 1240 56756 1280
rect 56620 1072 56660 1112
rect 57964 3424 58004 3464
rect 58156 4096 58196 4136
rect 58828 5524 58868 5564
rect 58732 5272 58772 5312
rect 58540 4768 58580 4808
rect 58444 4684 58484 4724
rect 58348 4096 58388 4136
rect 61132 5524 61172 5564
rect 58924 5272 58964 5312
rect 58732 4768 58772 4808
rect 58348 3760 58388 3800
rect 58732 3844 58772 3884
rect 58636 3676 58676 3716
rect 60460 5104 60500 5144
rect 59116 4684 59156 4724
rect 59020 4264 59060 4304
rect 59020 4096 59060 4136
rect 59020 3844 59060 3884
rect 58348 3424 58388 3464
rect 58924 3424 58964 3464
rect 59404 4264 59444 4304
rect 60844 4936 60884 4976
rect 60460 4768 60500 4808
rect 59596 4096 59636 4136
rect 60364 4096 60404 4136
rect 59116 3592 59156 3632
rect 58252 3340 58292 3380
rect 58636 3340 58676 3380
rect 59116 3340 59156 3380
rect 57676 2920 57716 2960
rect 58540 3256 58580 3296
rect 57964 2836 58004 2876
rect 58252 2752 58292 2792
rect 58636 2584 58676 2624
rect 58924 2584 58964 2624
rect 57004 2080 57044 2120
rect 57484 2080 57524 2120
rect 58060 2080 58100 2120
rect 57388 1996 57428 2036
rect 57196 1828 57236 1868
rect 57004 1660 57044 1700
rect 57868 1996 57908 2036
rect 58444 1996 58484 2036
rect 57100 1072 57140 1112
rect 57100 736 57140 776
rect 57772 1408 57812 1448
rect 57772 1072 57812 1112
rect 58156 1408 58196 1448
rect 58348 1072 58388 1112
rect 58732 1912 58772 1952
rect 58732 1660 58772 1700
rect 59116 2416 59156 2456
rect 59020 2080 59060 2120
rect 58924 1912 58964 1952
rect 59020 1660 59060 1700
rect 59116 1072 59156 1112
rect 59308 3424 59348 3464
rect 59308 1660 59348 1700
rect 59308 1240 59348 1280
rect 59308 904 59348 944
rect 60652 3676 60692 3716
rect 60652 2836 60692 2876
rect 60460 2584 60500 2624
rect 60556 2416 60596 2456
rect 59980 1912 60020 1952
rect 59500 1576 59540 1616
rect 59884 1240 59924 1280
rect 59596 1072 59636 1112
rect 59500 904 59540 944
rect 60460 1912 60500 1952
rect 60652 1744 60692 1784
rect 60268 1660 60308 1700
rect 60172 1492 60212 1532
rect 60172 1072 60212 1112
rect 60652 1240 60692 1280
rect 60652 1072 60692 1112
rect 60268 148 60308 188
rect 60556 904 60596 944
rect 61036 5440 61076 5480
rect 61228 5272 61268 5312
rect 61036 5104 61076 5144
rect 61516 5608 61556 5648
rect 61516 5272 61556 5312
rect 61420 5188 61460 5228
rect 61324 4936 61364 4976
rect 61228 4852 61268 4892
rect 61036 4684 61076 4724
rect 60940 4600 60980 4640
rect 61324 4684 61364 4724
rect 61900 5608 61940 5648
rect 62572 5608 62612 5648
rect 71884 5608 71924 5648
rect 73324 5608 73364 5648
rect 61996 5440 62036 5480
rect 62380 5440 62420 5480
rect 61900 5272 61940 5312
rect 61804 5020 61844 5060
rect 62188 5020 62228 5060
rect 61228 4012 61268 4052
rect 60940 2836 60980 2876
rect 61516 3928 61556 3968
rect 61708 4936 61748 4976
rect 61900 4936 61940 4976
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 62092 4852 62132 4892
rect 61900 4096 61940 4136
rect 62380 4684 62420 4724
rect 62092 4516 62132 4556
rect 62668 4936 62708 4976
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 62668 4432 62708 4472
rect 67180 4936 67220 4976
rect 73324 4936 73364 4976
rect 69100 4768 69140 4808
rect 66892 4348 66932 4388
rect 62476 4264 62516 4304
rect 62476 4096 62516 4136
rect 66508 4096 66548 4136
rect 62284 4012 62324 4052
rect 61804 3928 61844 3968
rect 61996 3928 62036 3968
rect 61420 2752 61460 2792
rect 61324 2668 61364 2708
rect 61804 2752 61844 2792
rect 60940 2584 60980 2624
rect 61420 2584 61460 2624
rect 61708 2584 61748 2624
rect 61996 2668 62036 2708
rect 60940 1240 60980 1280
rect 61132 1072 61172 1112
rect 61324 2416 61364 2456
rect 61036 904 61076 944
rect 61900 1828 61940 1868
rect 66988 4096 67028 4136
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 64012 3676 64052 3716
rect 63148 3424 63188 3464
rect 63436 3424 63476 3464
rect 63820 3424 63860 3464
rect 66604 3928 66644 3968
rect 66796 3928 66836 3968
rect 66412 3844 66452 3884
rect 65452 3508 65492 3548
rect 65644 3508 65684 3548
rect 66028 3508 66068 3548
rect 66316 3508 66356 3548
rect 63340 3256 63380 3296
rect 62860 2752 62900 2792
rect 63052 2584 63092 2624
rect 62572 1912 62612 1952
rect 62380 1828 62420 1868
rect 63052 1324 63092 1364
rect 62476 904 62516 944
rect 63052 1156 63092 1196
rect 62668 1072 62708 1112
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 63340 2752 63380 2792
rect 63532 2584 63572 2624
rect 64204 3424 64244 3464
rect 64204 2920 64244 2960
rect 64204 2584 64244 2624
rect 64108 2248 64148 2288
rect 64012 1660 64052 1700
rect 64588 3424 64628 3464
rect 65260 3424 65300 3464
rect 64780 3340 64820 3380
rect 64396 3004 64436 3044
rect 64396 2164 64436 2204
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 65836 3424 65876 3464
rect 65452 3340 65492 3380
rect 66220 3424 66260 3464
rect 65356 3172 65396 3212
rect 65068 1912 65108 1952
rect 64204 1324 64244 1364
rect 64684 1324 64724 1364
rect 63724 1240 63764 1280
rect 62764 904 62804 944
rect 62865 904 62905 944
rect 63244 1072 63284 1112
rect 63244 904 63284 944
rect 64876 1240 64916 1280
rect 63532 1156 63572 1196
rect 63628 1072 63668 1112
rect 64012 1156 64052 1196
rect 64396 1156 64436 1196
rect 62860 484 62900 524
rect 63532 904 63572 944
rect 64300 1072 64340 1112
rect 64780 1156 64820 1196
rect 64588 1072 64628 1112
rect 65164 1156 65204 1196
rect 64972 988 65012 1028
rect 63820 904 63860 944
rect 63724 736 63764 776
rect 63628 484 63668 524
rect 64204 904 64244 944
rect 64300 904 64340 944
rect 64876 904 64916 944
rect 65068 904 65108 944
rect 63916 484 63956 524
rect 64204 64 64244 104
rect 64684 736 64724 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 64588 484 64628 524
rect 65548 1156 65588 1196
rect 65452 1072 65492 1112
rect 65356 904 65396 944
rect 65164 400 65204 440
rect 65548 904 65588 944
rect 65932 1156 65972 1196
rect 65740 1072 65780 1112
rect 65452 400 65492 440
rect 65836 904 65876 944
rect 68524 4180 68564 4220
rect 69100 4180 69140 4220
rect 73804 4936 73844 4976
rect 74284 4936 74324 4976
rect 73612 4264 73652 4304
rect 74188 4600 74228 4640
rect 74092 4432 74132 4472
rect 74092 4264 74132 4304
rect 73324 4096 73364 4136
rect 74380 4768 74420 4808
rect 82156 4936 82196 4976
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 80524 4432 80564 4472
rect 74476 4264 74516 4304
rect 74668 4264 74708 4304
rect 74284 4180 74324 4220
rect 74188 4096 74228 4136
rect 74380 4096 74420 4136
rect 67180 3928 67220 3968
rect 68428 3928 68468 3968
rect 66796 3424 66836 3464
rect 66988 3256 67028 3296
rect 66796 2500 66836 2540
rect 66604 2332 66644 2372
rect 66316 1156 66356 1196
rect 66124 1072 66164 1112
rect 65932 484 65972 524
rect 66892 1324 66932 1364
rect 66508 1240 66548 1280
rect 66700 1156 66740 1196
rect 66220 484 66260 524
rect 66316 400 66356 440
rect 66700 904 66740 944
rect 66604 400 66644 440
rect 67372 3592 67412 3632
rect 67180 3424 67220 3464
rect 68620 3508 68660 3548
rect 68908 3928 68948 3968
rect 74764 4180 74804 4220
rect 74860 4096 74900 4136
rect 80332 4096 80372 4136
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 82828 4936 82868 4976
rect 93676 4936 93716 4976
rect 82348 4852 82388 4892
rect 91756 4768 91796 4808
rect 82060 4348 82100 4388
rect 86572 4600 86612 4640
rect 82156 4180 82196 4220
rect 86668 4180 86708 4220
rect 72076 3760 72116 3800
rect 70156 3676 70196 3716
rect 68812 3424 68852 3464
rect 67372 3256 67412 3296
rect 67084 1156 67124 1196
rect 67084 904 67124 944
rect 67372 3004 67412 3044
rect 67372 2584 67412 2624
rect 67564 2416 67604 2456
rect 67852 1912 67892 1952
rect 67276 1156 67316 1196
rect 67468 1072 67508 1112
rect 66796 568 66836 608
rect 66796 400 66836 440
rect 67372 904 67412 944
rect 67852 1072 67892 1112
rect 67468 652 67508 692
rect 68044 1156 68084 1196
rect 68236 1072 68276 1112
rect 67852 652 67892 692
rect 67756 568 67796 608
rect 67852 484 67892 524
rect 67756 148 67796 188
rect 68236 904 68276 944
rect 68716 1576 68756 1616
rect 68428 1072 68468 1112
rect 68620 1072 68660 1112
rect 68140 484 68180 524
rect 68524 904 68564 944
rect 68812 1072 68852 1112
rect 69772 3508 69812 3548
rect 69196 3424 69236 3464
rect 69004 2668 69044 2708
rect 69004 2164 69044 2204
rect 69580 3424 69620 3464
rect 69964 3424 70004 3464
rect 71308 3508 71348 3548
rect 71692 3508 71732 3548
rect 70348 3424 70388 3464
rect 70732 3424 70772 3464
rect 70540 3256 70580 3296
rect 69388 3088 69428 3128
rect 69388 2836 69428 2876
rect 69100 1576 69140 1616
rect 69388 1408 69428 1448
rect 69004 1072 69044 1112
rect 68620 652 68660 692
rect 69196 1072 69236 1112
rect 68908 652 68948 692
rect 69004 484 69044 524
rect 69388 904 69428 944
rect 69772 1156 69812 1196
rect 69676 1072 69716 1112
rect 69292 484 69332 524
rect 69676 904 69716 944
rect 71116 3424 71156 3464
rect 71500 3424 71540 3464
rect 71884 3424 71924 3464
rect 73324 3592 73364 3632
rect 71692 3340 71732 3380
rect 70924 3004 70964 3044
rect 70924 2752 70964 2792
rect 70732 1492 70772 1532
rect 70252 1240 70292 1280
rect 70636 1240 70676 1280
rect 70156 1156 70196 1196
rect 69964 1072 70004 1112
rect 69772 484 69812 524
rect 70156 904 70196 944
rect 70060 484 70100 524
rect 70521 1156 70561 1196
rect 70348 1072 70388 1112
rect 70636 1072 70676 1112
rect 70444 904 70484 944
rect 70924 1492 70964 1532
rect 72268 3424 72308 3464
rect 72652 3424 72692 3464
rect 72844 3424 72884 3464
rect 72460 3340 72500 3380
rect 72076 2920 72116 2960
rect 70540 148 70580 188
rect 71788 1324 71828 1364
rect 71116 1072 71156 1112
rect 72076 1156 72116 1196
rect 71500 1072 71540 1112
rect 71308 988 71348 1028
rect 71212 904 71252 944
rect 71500 820 71540 860
rect 70924 484 70964 524
rect 70828 232 70868 272
rect 71308 484 71348 524
rect 71692 904 71732 944
rect 71596 484 71636 524
rect 71884 1072 71924 1112
rect 71884 904 71924 944
rect 72076 904 72116 944
rect 71884 736 71924 776
rect 71788 568 71828 608
rect 71788 316 71828 356
rect 73036 3340 73076 3380
rect 72460 3088 72500 3128
rect 72268 1324 72308 1364
rect 72268 1072 72308 1112
rect 72940 2668 72980 2708
rect 73132 2668 73172 2708
rect 73708 3172 73748 3212
rect 73516 2668 73556 2708
rect 73900 2668 73940 2708
rect 73708 2584 73748 2624
rect 73324 2500 73364 2540
rect 77932 3760 77972 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 76012 3676 76052 3716
rect 76780 3676 76820 3716
rect 75148 3424 75188 3464
rect 74092 2668 74132 2708
rect 74284 2500 74324 2540
rect 74764 2752 74804 2792
rect 74956 2668 74996 2708
rect 74668 2164 74708 2204
rect 74764 1912 74804 1952
rect 73996 1408 74036 1448
rect 72460 1156 72500 1196
rect 72844 1240 72884 1280
rect 72652 1072 72692 1112
rect 72172 736 72212 776
rect 72460 484 72500 524
rect 72844 904 72884 944
rect 73036 1072 73076 1112
rect 72748 484 72788 524
rect 73132 904 73172 944
rect 73612 1156 73652 1196
rect 73420 1072 73460 1112
rect 73228 652 73268 692
rect 73324 484 73364 524
rect 73132 400 73172 440
rect 73612 904 73652 944
rect 73996 1156 74036 1196
rect 73804 1072 73844 1112
rect 73516 484 73556 524
rect 73900 904 73940 944
rect 74188 1072 74228 1112
rect 73996 232 74036 272
rect 74380 904 74420 944
rect 74956 1408 74996 1448
rect 74860 1324 74900 1364
rect 74572 1072 74612 1112
rect 74764 1072 74804 1112
rect 74380 484 74420 524
rect 74284 232 74324 272
rect 74764 904 74804 944
rect 75532 3424 75572 3464
rect 75820 3424 75860 3464
rect 75340 2836 75380 2876
rect 75340 2332 75380 2372
rect 76204 3424 76244 3464
rect 76012 3340 76052 3380
rect 77644 3508 77684 3548
rect 77932 3508 77972 3548
rect 76588 3424 76628 3464
rect 76396 3256 76436 3296
rect 75820 2668 75860 2708
rect 75628 2584 75668 2624
rect 76396 2920 76436 2960
rect 75052 1324 75092 1364
rect 74956 1072 74996 1112
rect 74668 484 74708 524
rect 75052 904 75092 944
rect 75532 1240 75572 1280
rect 75340 1073 75380 1112
rect 75340 1072 75380 1073
rect 75148 820 75188 860
rect 75148 484 75188 524
rect 75532 904 75572 944
rect 75724 1072 75764 1112
rect 75916 1072 75956 1112
rect 75436 484 75476 524
rect 75820 904 75860 944
rect 76972 3424 77012 3464
rect 77452 3424 77492 3464
rect 76684 3004 76724 3044
rect 76108 1072 76148 1112
rect 76300 1072 76340 1112
rect 75916 484 75956 524
rect 76300 904 76340 944
rect 76204 484 76244 524
rect 76492 988 76532 1028
rect 76588 904 76628 944
rect 76684 820 76724 860
rect 78124 3424 78164 3464
rect 77260 2584 77300 2624
rect 77164 2500 77204 2540
rect 77452 1576 77492 1616
rect 77068 1492 77108 1532
rect 76876 988 76916 1028
rect 76684 484 76724 524
rect 77068 904 77108 944
rect 76972 484 77012 524
rect 77260 988 77300 1028
rect 77452 988 77492 1028
rect 77356 904 77396 944
rect 78508 3424 78548 3464
rect 78220 3088 78260 3128
rect 77644 1072 77684 1112
rect 77260 484 77300 524
rect 77452 484 77492 524
rect 77164 148 77204 188
rect 78988 3424 79028 3464
rect 79180 3424 79220 3464
rect 78988 3256 79028 3296
rect 79372 3256 79412 3296
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 78796 2584 78836 2624
rect 78220 2416 78260 2456
rect 78028 1072 78068 1112
rect 77836 568 77876 608
rect 77740 484 77780 524
rect 77836 400 77876 440
rect 78220 904 78260 944
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 78412 1072 78452 1112
rect 78604 988 78644 1028
rect 78124 400 78164 440
rect 78316 400 78356 440
rect 79180 1240 79220 1280
rect 79372 1240 79412 1280
rect 78796 1072 78836 1112
rect 78604 484 78644 524
rect 78508 400 78548 440
rect 78988 904 79028 944
rect 78892 484 78932 524
rect 79276 904 79316 944
rect 79756 3256 79796 3296
rect 80332 3424 80372 3464
rect 80140 3256 80180 3296
rect 79564 2752 79604 2792
rect 79948 3172 79988 3212
rect 80236 3172 80276 3212
rect 79948 2668 79988 2708
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 79948 1828 79988 1868
rect 79852 1576 79892 1616
rect 80044 1576 80084 1616
rect 79756 1492 79796 1532
rect 79564 1240 79604 1280
rect 79564 1072 79604 1112
rect 80044 1324 80084 1364
rect 79948 1072 79988 1112
rect 80812 4096 80852 4136
rect 86572 4096 86612 4136
rect 87052 4096 87092 4136
rect 87244 4096 87284 4136
rect 91564 4096 91604 4136
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 80620 3172 80660 3212
rect 80524 1324 80564 1364
rect 80428 1240 80468 1280
rect 80332 1072 80372 1112
rect 79372 652 79412 692
rect 79180 484 79220 524
rect 79084 316 79124 356
rect 79372 316 79412 356
rect 79756 904 79796 944
rect 80044 904 80084 944
rect 80236 904 80276 944
rect 79660 316 79700 356
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 79948 568 79988 608
rect 80524 904 80564 944
rect 80332 316 80372 356
rect 80812 1912 80852 1952
rect 82924 3676 82964 3716
rect 81292 3424 81332 3464
rect 81676 3424 81716 3464
rect 81484 3256 81524 3296
rect 81100 3088 81140 3128
rect 81100 2164 81140 2204
rect 80620 316 80660 356
rect 80908 1240 80948 1280
rect 81100 1240 81140 1280
rect 81484 2332 81524 2372
rect 81484 1408 81524 1448
rect 81292 1156 81332 1196
rect 82348 3424 82388 3464
rect 82156 3340 82196 3380
rect 81868 2584 81908 2624
rect 81676 1156 81716 1196
rect 81868 1072 81908 1112
rect 82060 1156 82100 1196
rect 82252 1072 82292 1112
rect 82732 3424 82772 3464
rect 83788 3592 83828 3632
rect 83116 3424 83156 3464
rect 82540 2920 82580 2960
rect 82444 1156 82484 1196
rect 82636 1072 82676 1112
rect 82828 1324 82868 1364
rect 82828 1156 82868 1196
rect 83020 1072 83060 1112
rect 83596 3424 83636 3464
rect 84172 3508 84212 3548
rect 83980 3424 84020 3464
rect 83692 3172 83732 3212
rect 83404 2584 83444 2624
rect 84364 3424 84404 3464
rect 84556 3424 84596 3464
rect 84172 2836 84212 2876
rect 84364 2584 84404 2624
rect 83884 1408 83924 1448
rect 83212 1156 83252 1196
rect 83308 1072 83348 1112
rect 83596 1156 83636 1196
rect 83980 1156 84020 1196
rect 82828 736 82868 776
rect 83788 736 83828 776
rect 84172 1072 84212 1112
rect 84364 1156 84404 1196
rect 84556 1072 84596 1112
rect 84940 2752 84980 2792
rect 86092 2752 86132 2792
rect 84748 2584 84788 2624
rect 85324 2668 85364 2708
rect 85132 2584 85172 2624
rect 85900 2668 85940 2708
rect 85516 2584 85556 2624
rect 85708 2584 85748 2624
rect 85228 2500 85268 2540
rect 86284 2668 86324 2708
rect 86476 2584 86516 2624
rect 84748 1156 84788 1196
rect 84940 1072 84980 1112
rect 85324 1324 85364 1364
rect 85132 1156 85172 1196
rect 83884 484 83924 524
rect 85516 1156 85556 1196
rect 85324 820 85364 860
rect 85708 1492 85748 1532
rect 85708 1240 85748 1280
rect 85900 1156 85940 1196
rect 86092 1576 86132 1616
rect 86284 1156 86324 1196
rect 85612 820 85652 860
rect 85708 736 85748 776
rect 85612 652 85652 692
rect 85612 316 85652 356
rect 86476 1072 86516 1112
rect 87052 3424 87092 3464
rect 86764 1912 86804 1952
rect 86668 1156 86708 1196
rect 86860 1072 86900 1112
rect 87047 1156 87087 1196
rect 91660 4012 91700 4052
rect 92044 4096 92084 4136
rect 93580 4012 93620 4052
rect 88780 3760 88820 3800
rect 87628 3508 87668 3548
rect 87436 3424 87476 3464
rect 87820 3424 87860 3464
rect 87628 3256 87668 3296
rect 87244 3088 87284 3128
rect 87244 1072 87284 1112
rect 87628 1240 87668 1280
rect 87436 1072 87476 1112
rect 88204 3424 88244 3464
rect 88588 3424 88628 3464
rect 89164 3676 89204 3716
rect 88396 3340 88436 3380
rect 88012 2668 88052 2708
rect 88012 1156 88052 1196
rect 87820 1072 87860 1112
rect 88396 1408 88436 1448
rect 88204 1072 88244 1112
rect 88972 3424 89012 3464
rect 89932 3592 89972 3632
rect 90700 3592 90740 3632
rect 92236 3592 92276 3632
rect 93100 3592 93140 3632
rect 93484 3592 93524 3632
rect 89356 3424 89396 3464
rect 89164 3256 89204 3296
rect 88780 2920 88820 2960
rect 88780 1324 88820 1364
rect 88588 1072 88628 1112
rect 89164 1156 89204 1196
rect 88972 1072 89012 1112
rect 86188 316 86228 356
rect 89740 3424 89780 3464
rect 90124 3424 90164 3464
rect 89548 2584 89588 2624
rect 89356 1324 89396 1364
rect 89548 1156 89588 1196
rect 89356 1072 89396 1112
rect 89932 3172 89972 3212
rect 89740 1324 89780 1364
rect 89932 1240 89972 1280
rect 90508 3424 90548 3464
rect 90892 3424 90932 3464
rect 90316 3004 90356 3044
rect 90316 2836 90356 2876
rect 90124 1324 90164 1364
rect 90316 1240 90356 1280
rect 90508 1324 90548 1364
rect 90700 988 90740 1028
rect 91276 3424 91316 3464
rect 91084 2500 91124 2540
rect 91084 2332 91124 2372
rect 90892 1324 90932 1364
rect 91084 1072 91124 1112
rect 91660 3424 91700 3464
rect 91468 2836 91508 2876
rect 91276 1324 91316 1364
rect 91468 1072 91508 1112
rect 92044 3424 92084 3464
rect 91852 2668 91892 2708
rect 91660 1324 91700 1364
rect 91852 1072 91892 1112
rect 92428 3424 92468 3464
rect 92620 3424 92660 3464
rect 92812 3424 92852 3464
rect 92236 2920 92276 2960
rect 92044 1324 92084 1364
rect 90988 652 91028 692
rect 90988 484 91028 524
rect 92716 2584 92756 2624
rect 92524 1912 92564 1952
rect 92620 1660 92660 1700
rect 92908 3088 92948 3128
rect 93292 3424 93332 3464
rect 93100 2584 93140 2624
rect 93004 2416 93044 2456
rect 93100 1660 93140 1700
rect 92428 1324 92468 1364
rect 92620 1240 92660 1280
rect 92428 1072 92468 1112
rect 92812 1072 92852 1112
rect 93004 1072 93044 1112
rect 92140 232 92180 272
rect 93196 1240 93236 1280
rect 94444 3760 94484 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 94252 3592 94292 3632
rect 94060 3424 94100 3464
rect 94636 3676 94676 3716
rect 94636 3508 94676 3548
rect 95020 3508 95060 3548
rect 95308 3508 95348 3548
rect 95692 3508 95732 3548
rect 96172 3508 96212 3548
rect 96556 3508 96596 3548
rect 94828 3424 94868 3464
rect 94348 3340 94388 3380
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 93676 2668 93716 2708
rect 93772 2584 93812 2624
rect 93484 2416 93524 2456
rect 93292 1072 93332 1112
rect 93395 1072 93428 1112
rect 93428 1072 93435 1112
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 94348 2836 94388 2876
rect 94636 1492 94676 1532
rect 95116 2584 95156 2624
rect 95500 3172 95540 3212
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 94348 1408 94388 1448
rect 94924 1408 94964 1448
rect 93580 1072 93620 1112
rect 93772 988 93812 1028
rect 94252 1240 94292 1280
rect 93964 1072 94004 1112
rect 94156 1072 94196 1112
rect 94732 1109 94772 1112
rect 94732 1072 94772 1109
rect 94540 988 94580 1028
rect 94924 988 94964 1028
rect 95111 988 95151 1028
rect 95308 988 95348 1028
rect 95980 3088 96020 3128
rect 98188 3340 98228 3380
rect 98092 2920 98132 2960
rect 97516 2752 97556 2792
rect 96556 2668 96596 2708
rect 96940 2668 96980 2708
rect 97324 2668 97364 2708
rect 96364 2584 96404 2624
rect 96748 2584 96788 2624
rect 97132 2584 97172 2624
rect 97708 2668 97748 2708
rect 97900 2668 97940 2708
rect 97036 1492 97076 1532
rect 95596 1240 95636 1280
rect 96172 1240 96212 1280
rect 96076 1156 96116 1196
rect 95500 1072 95540 1112
rect 93868 904 93908 944
rect 93772 820 93812 860
rect 94156 904 94196 944
rect 94732 904 94772 944
rect 94828 904 94868 944
rect 95212 904 95252 944
rect 95404 904 95444 944
rect 94540 820 94580 860
rect 94636 736 94676 776
rect 94636 568 94676 608
rect 94828 736 94868 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
rect 95308 568 95348 608
rect 95116 64 95156 104
rect 95692 904 95732 944
rect 95884 1072 95924 1112
rect 96460 1156 96500 1196
rect 96268 1072 96308 1112
rect 96844 1156 96884 1196
rect 96652 1072 96692 1112
rect 97612 2500 97652 2540
rect 97228 1156 97268 1196
rect 97612 1156 97652 1196
rect 97036 1072 97076 1112
rect 95788 820 95828 860
rect 97228 736 97268 776
rect 97996 1324 98036 1364
rect 97996 1156 98036 1196
rect 97324 400 97364 440
rect 97996 904 98036 944
rect 97708 148 97748 188
rect 98380 1156 98420 1196
rect 98860 1240 98900 1280
rect 98764 1156 98804 1196
rect 98188 820 98228 860
rect 98092 232 98132 272
rect 98668 1072 98708 1112
rect 98476 316 98516 356
rect 98956 1156 98996 1196
rect 99148 1072 99188 1112
<< metal3 >>
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 6211 6952 6220 6992
rect 6260 6952 24556 6992
rect 24596 6952 24605 6992
rect 28099 6952 28108 6992
rect 28148 6952 41068 6992
rect 41108 6952 41740 6992
rect 41780 6952 41789 6992
rect 17155 6868 17164 6908
rect 17204 6868 41356 6908
rect 41396 6868 42028 6908
rect 42068 6868 42077 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 39043 6616 39052 6656
rect 39092 6616 46732 6656
rect 46772 6616 47596 6656
rect 47636 6616 48460 6656
rect 48500 6616 49036 6656
rect 49076 6616 49085 6656
rect 41731 6532 41740 6572
rect 41780 6532 44716 6572
rect 44756 6532 45772 6572
rect 45812 6532 46348 6572
rect 46388 6532 46397 6572
rect 46531 6532 46540 6572
rect 46580 6532 46589 6572
rect 46540 6488 46580 6532
rect 42019 6448 42028 6488
rect 42068 6448 44524 6488
rect 44564 6448 45868 6488
rect 45908 6448 46580 6488
rect 46627 6448 46636 6488
rect 46676 6448 47884 6488
rect 47924 6448 48556 6488
rect 48596 6448 48748 6488
rect 48788 6448 49420 6488
rect 49460 6448 49469 6488
rect 46819 6280 46828 6320
rect 46868 6280 56428 6320
rect 56468 6280 56477 6320
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 24547 5608 24556 5648
rect 24596 5608 41452 5648
rect 41492 5608 41501 5648
rect 44323 5608 44332 5648
rect 44372 5608 44524 5648
rect 44564 5608 45004 5648
rect 45044 5608 45053 5648
rect 49507 5608 49516 5648
rect 49556 5608 53740 5648
rect 53780 5608 54508 5648
rect 54548 5608 55460 5648
rect 56323 5608 56332 5648
rect 56372 5608 56812 5648
rect 56852 5608 61516 5648
rect 61556 5608 61565 5648
rect 61891 5608 61900 5648
rect 61940 5608 62572 5648
rect 62612 5608 71884 5648
rect 71924 5608 73324 5648
rect 73364 5608 73373 5648
rect 55420 5564 55460 5608
rect 61900 5564 61940 5608
rect 44611 5524 44620 5564
rect 44660 5524 44908 5564
rect 44948 5524 46348 5564
rect 46388 5524 46540 5564
rect 46580 5524 47596 5564
rect 47636 5524 51916 5564
rect 51956 5524 52780 5564
rect 52820 5524 52829 5564
rect 55420 5524 58828 5564
rect 58868 5524 58877 5564
rect 61123 5524 61132 5564
rect 61172 5524 61940 5564
rect 41443 5440 41452 5480
rect 41492 5440 41836 5480
rect 41876 5440 42124 5480
rect 42164 5440 42173 5480
rect 61027 5440 61036 5480
rect 61076 5440 61996 5480
rect 62036 5440 62380 5480
rect 62420 5440 62429 5480
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 51235 5272 51244 5312
rect 51284 5272 52588 5312
rect 52628 5272 53740 5312
rect 53780 5272 55084 5312
rect 55124 5272 55564 5312
rect 55604 5272 58060 5312
rect 58100 5272 58732 5312
rect 58772 5272 58924 5312
rect 58964 5272 61228 5312
rect 61268 5272 61516 5312
rect 61556 5272 61900 5312
rect 61940 5272 61949 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 42211 5228 42269 5229
rect 41539 5188 41548 5228
rect 41588 5188 42220 5228
rect 42260 5188 42269 5228
rect 56419 5188 56428 5228
rect 56468 5188 61420 5228
rect 61460 5188 61469 5228
rect 42211 5187 42269 5188
rect 46051 5144 46109 5145
rect 55363 5144 55421 5145
rect 44323 5104 44332 5144
rect 44372 5104 44812 5144
rect 44852 5104 45004 5144
rect 45044 5104 45868 5144
rect 45908 5104 46060 5144
rect 46100 5104 46156 5144
rect 46196 5104 46636 5144
rect 46676 5104 48076 5144
rect 48116 5104 48844 5144
rect 48884 5104 49324 5144
rect 49364 5104 49373 5144
rect 50659 5104 50668 5144
rect 50708 5104 50717 5144
rect 55278 5104 55372 5144
rect 55412 5104 55421 5144
rect 60451 5104 60460 5144
rect 60500 5104 61036 5144
rect 61076 5104 61085 5144
rect 46051 5103 46109 5104
rect 50668 5060 50708 5104
rect 55363 5103 55421 5104
rect 41539 5020 41548 5060
rect 41588 5020 41740 5060
rect 41780 5020 42028 5060
rect 42068 5020 42700 5060
rect 42740 5020 44620 5060
rect 44660 5020 44669 5060
rect 49603 5020 49612 5060
rect 49652 5020 50708 5060
rect 50851 5020 50860 5060
rect 50900 5020 50909 5060
rect 52003 5020 52012 5060
rect 52052 5020 52300 5060
rect 52340 5020 52684 5060
rect 52724 5020 58156 5060
rect 58196 5020 58205 5060
rect 60748 5020 61804 5060
rect 61844 5020 62188 5060
rect 62228 5020 62237 5060
rect 50371 4976 50429 4977
rect 50860 4976 50900 5020
rect 60748 4976 60788 5020
rect 41347 4936 41356 4976
rect 41396 4936 41644 4976
rect 41684 4936 42124 4976
rect 42164 4936 42173 4976
rect 45955 4936 45964 4976
rect 46004 4936 46636 4976
rect 46676 4936 46685 4976
rect 48163 4936 48172 4976
rect 48212 4936 48748 4976
rect 48788 4936 49036 4976
rect 49076 4936 49085 4976
rect 50286 4936 50380 4976
rect 50420 4936 50900 4976
rect 51523 4936 51532 4976
rect 51572 4936 52204 4976
rect 52244 4936 52253 4976
rect 52387 4936 52396 4976
rect 52436 4936 52445 4976
rect 52963 4936 52972 4976
rect 53012 4936 53548 4976
rect 53588 4936 54316 4976
rect 54356 4936 54365 4976
rect 56419 4936 56428 4976
rect 56468 4936 60788 4976
rect 60835 4936 60844 4976
rect 60884 4936 60893 4976
rect 61315 4936 61324 4976
rect 61364 4936 61708 4976
rect 61748 4936 61900 4976
rect 61940 4936 61949 4976
rect 62659 4936 62668 4976
rect 62708 4936 67180 4976
rect 67220 4936 68060 4976
rect 73315 4936 73324 4976
rect 73364 4936 73804 4976
rect 73844 4936 74284 4976
rect 74324 4936 74333 4976
rect 82147 4936 82156 4976
rect 82196 4936 82828 4976
rect 82868 4936 82877 4976
rect 85660 4936 93676 4976
rect 93716 4936 93725 4976
rect 50371 4935 50429 4936
rect 50860 4892 50900 4936
rect 52396 4892 52436 4936
rect 45859 4852 45868 4892
rect 45908 4852 46252 4892
rect 46292 4852 48268 4892
rect 48308 4852 50476 4892
rect 50516 4852 50525 4892
rect 50860 4852 52876 4892
rect 52916 4852 53836 4892
rect 53876 4852 53885 4892
rect 54403 4852 54412 4892
rect 54452 4852 55180 4892
rect 55220 4852 60500 4892
rect 48355 4808 48413 4809
rect 48931 4808 48989 4809
rect 54892 4808 54932 4852
rect 60460 4808 60500 4852
rect 60844 4808 60884 4936
rect 68020 4892 68060 4936
rect 85660 4892 85700 4936
rect 61219 4852 61228 4892
rect 61268 4852 62092 4892
rect 62132 4852 62141 4892
rect 68020 4852 82348 4892
rect 82388 4852 85700 4892
rect 48355 4768 48364 4808
rect 48404 4768 48556 4808
rect 48596 4768 48605 4808
rect 48835 4768 48844 4808
rect 48884 4768 48940 4808
rect 48980 4768 48989 4808
rect 49315 4768 49324 4808
rect 49364 4768 51244 4808
rect 51284 4768 51293 4808
rect 51523 4768 51532 4808
rect 51572 4768 53452 4808
rect 53492 4768 53740 4808
rect 53780 4768 53789 4808
rect 54883 4768 54892 4808
rect 54932 4768 54941 4808
rect 55276 4768 55948 4808
rect 55988 4768 56332 4808
rect 56372 4768 56381 4808
rect 58051 4768 58060 4808
rect 58100 4768 58540 4808
rect 58580 4768 58732 4808
rect 58772 4768 58781 4808
rect 60451 4768 60460 4808
rect 60500 4768 60884 4808
rect 69091 4768 69100 4808
rect 69140 4768 74380 4808
rect 74420 4768 91756 4808
rect 91796 4768 91805 4808
rect 48355 4767 48413 4768
rect 48931 4767 48989 4768
rect 55276 4724 55316 4768
rect 62371 4724 62429 4725
rect 50371 4684 50380 4724
rect 50420 4684 50668 4724
rect 50708 4684 55316 4724
rect 58435 4684 58444 4724
rect 58484 4684 59116 4724
rect 59156 4684 59165 4724
rect 61027 4684 61036 4724
rect 61076 4684 61324 4724
rect 61364 4684 61373 4724
rect 62286 4684 62380 4724
rect 62420 4684 62429 4724
rect 62371 4683 62429 4684
rect 53827 4600 53836 4640
rect 53876 4600 54796 4640
rect 54836 4600 55372 4640
rect 55412 4600 60940 4640
rect 60980 4600 60989 4640
rect 74179 4600 74188 4640
rect 74228 4600 86572 4640
rect 86612 4600 86621 4640
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 18883 4516 18892 4556
rect 18932 4516 19468 4556
rect 19508 4516 20044 4556
rect 20084 4516 20093 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 38659 4516 38668 4556
rect 38708 4516 43948 4556
rect 43988 4516 43997 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 50179 4516 50188 4556
rect 50228 4516 51820 4556
rect 51860 4516 55276 4556
rect 55316 4516 55660 4556
rect 55700 4516 57964 4556
rect 58004 4516 58013 4556
rect 62083 4516 62092 4556
rect 62132 4516 62804 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 62764 4472 62804 4516
rect 38947 4432 38956 4472
rect 38996 4432 62668 4472
rect 62708 4432 62717 4472
rect 62764 4432 74092 4472
rect 74132 4432 80524 4472
rect 80564 4432 80573 4472
rect 38659 4388 38717 4389
rect 52099 4388 52157 4389
rect 52483 4388 52541 4389
rect 66787 4388 66845 4389
rect 18499 4348 18508 4388
rect 18548 4348 19084 4388
rect 19124 4348 19133 4388
rect 19747 4348 19756 4388
rect 19796 4348 37324 4388
rect 37364 4348 38188 4388
rect 38228 4348 38668 4388
rect 38708 4348 38717 4388
rect 41251 4348 41260 4388
rect 41300 4348 41740 4388
rect 41780 4348 41789 4388
rect 41923 4348 41932 4388
rect 41972 4348 42796 4388
rect 42836 4348 48076 4388
rect 48116 4348 50668 4388
rect 50708 4348 51436 4388
rect 51476 4348 51485 4388
rect 52099 4348 52108 4388
rect 52148 4348 52204 4388
rect 52244 4348 52253 4388
rect 52483 4348 52492 4388
rect 52532 4348 52588 4388
rect 52628 4348 52637 4388
rect 66787 4348 66796 4388
rect 66836 4348 66892 4388
rect 66932 4348 82060 4388
rect 82100 4348 82109 4388
rect 38659 4347 38717 4348
rect 52099 4347 52157 4348
rect 52483 4347 52541 4348
rect 66787 4347 66845 4348
rect 28003 4304 28061 4305
rect 6979 4264 6988 4304
rect 7028 4264 7564 4304
rect 7604 4264 25900 4304
rect 25940 4264 28012 4304
rect 28052 4264 28061 4304
rect 41443 4264 41452 4304
rect 41492 4264 41501 4304
rect 42115 4264 42124 4304
rect 42164 4264 42604 4304
rect 42644 4264 47788 4304
rect 47828 4264 47837 4304
rect 48163 4264 48172 4304
rect 48212 4264 48652 4304
rect 48692 4264 48701 4304
rect 49027 4264 49036 4304
rect 49076 4264 51532 4304
rect 51572 4264 51581 4304
rect 52204 4264 52972 4304
rect 53012 4264 53021 4304
rect 53347 4264 53356 4304
rect 53396 4264 53644 4304
rect 53684 4264 59020 4304
rect 59060 4264 59404 4304
rect 59444 4264 59453 4304
rect 62467 4264 62476 4304
rect 62516 4264 73612 4304
rect 73652 4264 74092 4304
rect 74132 4264 74476 4304
rect 74516 4264 74668 4304
rect 74708 4264 74717 4304
rect 28003 4263 28061 4264
rect 38947 4220 39005 4221
rect 7564 4180 22348 4220
rect 22388 4180 22397 4220
rect 24451 4180 24460 4220
rect 24500 4180 25132 4220
rect 25172 4180 37708 4220
rect 37748 4180 38476 4220
rect 38516 4180 38956 4220
rect 38996 4180 39005 4220
rect 41452 4220 41492 4264
rect 43180 4220 43220 4264
rect 52204 4220 52244 4264
rect 68515 4220 68573 4221
rect 41452 4180 42028 4220
rect 42068 4180 42077 4220
rect 43171 4180 43180 4220
rect 43220 4180 43229 4220
rect 44227 4180 44236 4220
rect 44276 4180 45100 4220
rect 45140 4180 46252 4220
rect 46292 4180 46301 4220
rect 46348 4180 46636 4220
rect 46676 4180 48844 4220
rect 48884 4180 49612 4220
rect 49652 4180 52204 4220
rect 52244 4180 52253 4220
rect 52780 4180 54892 4220
rect 54932 4180 54941 4220
rect 68430 4180 68524 4220
rect 68564 4180 69100 4220
rect 69140 4180 69149 4220
rect 74275 4180 74284 4220
rect 74324 4180 74764 4220
rect 74804 4180 74813 4220
rect 80812 4180 82156 4220
rect 82196 4180 86668 4220
rect 86708 4180 87284 4220
rect 7564 4136 7604 4180
rect 22348 4136 22388 4180
rect 38947 4179 39005 4180
rect 7171 4096 7180 4136
rect 7220 4096 7564 4136
rect 7604 4096 7613 4136
rect 18307 4096 18316 4136
rect 18356 4096 19756 4136
rect 19796 4096 19805 4136
rect 19939 4096 19948 4136
rect 19988 4096 22292 4136
rect 22348 4096 27916 4136
rect 27956 4096 32236 4136
rect 32276 4096 32812 4136
rect 32852 4096 37228 4136
rect 37268 4096 37804 4136
rect 37844 4096 38380 4136
rect 38420 4096 38429 4136
rect 41443 4096 41452 4136
rect 41492 4096 41932 4136
rect 41972 4096 41981 4136
rect 22252 4052 22292 4096
rect 26083 4052 26141 4053
rect 42028 4052 42068 4180
rect 44236 4052 44276 4180
rect 46051 4136 46109 4137
rect 46348 4136 46388 4180
rect 52780 4136 52820 4180
rect 68515 4179 68573 4180
rect 58627 4136 58685 4137
rect 66499 4136 66557 4137
rect 80812 4136 80852 4180
rect 87244 4136 87284 4180
rect 44323 4096 44332 4136
rect 44372 4096 44381 4136
rect 45966 4096 46060 4136
rect 46100 4096 46109 4136
rect 46339 4096 46348 4136
rect 46388 4096 46397 4136
rect 48355 4096 48364 4136
rect 48404 4096 48413 4136
rect 48547 4096 48556 4136
rect 48596 4096 48940 4136
rect 48980 4096 48989 4136
rect 50092 4096 50188 4136
rect 50228 4096 50237 4136
rect 50563 4096 50572 4136
rect 50612 4096 50956 4136
rect 50996 4096 51005 4136
rect 51427 4096 51436 4136
rect 51476 4096 52780 4136
rect 52820 4096 52829 4136
rect 53347 4096 53356 4136
rect 53396 4096 53836 4136
rect 53876 4096 53885 4136
rect 54787 4096 54796 4136
rect 54836 4096 55180 4136
rect 55220 4096 55229 4136
rect 57091 4096 57100 4136
rect 57140 4096 58156 4136
rect 58196 4096 58348 4136
rect 58388 4096 58636 4136
rect 58676 4096 59020 4136
rect 59060 4096 59596 4136
rect 59636 4096 60364 4136
rect 60404 4096 60413 4136
rect 61891 4096 61900 4136
rect 61940 4096 62476 4136
rect 62516 4096 62525 4136
rect 66414 4096 66508 4136
rect 66548 4096 66988 4136
rect 67028 4096 73324 4136
rect 73364 4096 74188 4136
rect 74228 4096 74237 4136
rect 74371 4096 74380 4136
rect 74420 4096 74860 4136
rect 74900 4096 80332 4136
rect 80372 4096 80812 4136
rect 80852 4096 80861 4136
rect 86563 4096 86572 4136
rect 86612 4096 87052 4136
rect 87092 4096 87101 4136
rect 87235 4096 87244 4136
rect 87284 4096 91564 4136
rect 91604 4096 92044 4136
rect 92084 4096 92093 4136
rect 18979 4012 18988 4052
rect 19028 4012 19180 4052
rect 19220 4012 20180 4052
rect 22252 4012 22444 4052
rect 22484 4012 24268 4052
rect 24308 4012 25036 4052
rect 25076 4012 26092 4052
rect 26132 4012 26141 4052
rect 18403 3928 18412 3968
rect 18452 3928 18892 3968
rect 18932 3928 19084 3968
rect 19124 3928 19133 3968
rect 19651 3928 19660 3968
rect 19700 3928 19948 3968
rect 19988 3928 19997 3968
rect 19660 3884 19700 3928
rect 18499 3844 18508 3884
rect 18548 3844 19700 3884
rect 20140 3884 20180 4012
rect 26083 4011 26141 4012
rect 37228 4012 38092 4052
rect 38132 4012 38956 4052
rect 38996 4012 39005 4052
rect 42028 4012 42508 4052
rect 42548 4012 43084 4052
rect 43124 4012 44276 4052
rect 37228 3968 37268 4012
rect 37708 3968 37748 4012
rect 38380 3968 38420 4012
rect 39235 3968 39293 3969
rect 44332 3968 44372 4096
rect 46051 4095 46109 4096
rect 48364 4052 48404 4096
rect 48931 4052 48989 4053
rect 44419 4012 44428 4052
rect 44468 4012 45004 4052
rect 45044 4012 48748 4052
rect 48788 4012 48940 4052
rect 48980 4012 48989 4052
rect 48931 4011 48989 4012
rect 50092 3968 50132 4096
rect 58627 4095 58685 4096
rect 66499 4095 66557 4096
rect 20227 3928 20236 3968
rect 20276 3928 24364 3968
rect 24404 3928 24940 3968
rect 24980 3928 32236 3968
rect 32276 3928 32524 3968
rect 32564 3928 37228 3968
rect 37268 3928 37277 3968
rect 37699 3928 37708 3968
rect 37748 3928 37788 3968
rect 38371 3928 38380 3968
rect 38420 3928 38460 3968
rect 39235 3928 39244 3968
rect 39284 3928 41260 3968
rect 41300 3928 41309 3968
rect 41635 3928 41644 3968
rect 41684 3928 42028 3968
rect 42068 3928 42316 3968
rect 42356 3928 42892 3968
rect 42932 3928 44372 3968
rect 47779 3928 47788 3968
rect 47828 3928 50132 3968
rect 51052 4012 61228 4052
rect 61268 4012 61277 4052
rect 61804 4012 62284 4052
rect 62324 4012 62333 4052
rect 91651 4012 91660 4052
rect 91700 4012 93580 4052
rect 93620 4012 93629 4052
rect 39235 3927 39293 3928
rect 51052 3884 51092 4012
rect 61804 3968 61844 4012
rect 51235 3928 51244 3968
rect 51284 3928 59828 3968
rect 61507 3928 61516 3968
rect 61556 3928 61804 3968
rect 61844 3928 61853 3968
rect 61987 3928 61996 3968
rect 62036 3928 66604 3968
rect 66644 3928 66796 3968
rect 66836 3928 67180 3968
rect 67220 3928 68428 3968
rect 68468 3928 68908 3968
rect 68948 3928 68957 3968
rect 59788 3884 59828 3928
rect 20140 3844 32140 3884
rect 32180 3844 32908 3884
rect 32948 3844 51092 3884
rect 54883 3844 54892 3884
rect 54932 3844 58732 3884
rect 58772 3844 59020 3884
rect 59060 3844 59069 3884
rect 59788 3844 66412 3884
rect 66452 3844 66461 3884
rect 19084 3800 19124 3844
rect 35683 3800 35741 3801
rect 44611 3800 44669 3801
rect 46051 3800 46109 3801
rect 58435 3800 58493 3801
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 9187 3760 9196 3800
rect 9236 3760 15244 3800
rect 15284 3760 15293 3800
rect 15340 3760 18796 3800
rect 18836 3760 18845 3800
rect 19075 3760 19084 3800
rect 19124 3760 19133 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 21091 3760 21100 3800
rect 21140 3760 27340 3800
rect 27380 3760 33004 3800
rect 33044 3760 33053 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 35598 3760 35692 3800
rect 35732 3760 35741 3800
rect 37987 3760 37996 3800
rect 38036 3760 43564 3800
rect 43604 3760 43613 3800
rect 44526 3760 44620 3800
rect 44660 3760 44669 3800
rect 45966 3760 46060 3800
rect 46100 3760 46109 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 53443 3760 53452 3800
rect 53492 3760 55084 3800
rect 55124 3760 55372 3800
rect 55412 3760 55421 3800
rect 55651 3760 55660 3800
rect 55700 3760 56620 3800
rect 56660 3760 56669 3800
rect 58339 3760 58348 3800
rect 58388 3760 58444 3800
rect 58484 3760 58493 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 72067 3760 72076 3800
rect 72116 3760 77932 3800
rect 77972 3760 77981 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 88771 3760 88780 3800
rect 88820 3760 94444 3800
rect 94484 3760 94493 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 15340 3716 15380 3760
rect 35683 3759 35741 3760
rect 44611 3759 44669 3760
rect 46051 3759 46109 3760
rect 58435 3759 58493 3760
rect 38083 3716 38141 3717
rect 47587 3716 47645 3717
rect 55363 3716 55421 3717
rect 8419 3676 8428 3716
rect 8468 3676 12020 3716
rect 12067 3676 12076 3716
rect 12116 3676 12460 3716
rect 12500 3676 15380 3716
rect 16771 3676 16780 3716
rect 16820 3676 21620 3716
rect 21667 3676 21676 3716
rect 21716 3676 27628 3716
rect 27668 3676 33388 3716
rect 33428 3676 38092 3716
rect 38132 3676 38141 3716
rect 38275 3676 38284 3716
rect 38324 3676 41740 3716
rect 41780 3676 44236 3716
rect 44276 3676 44285 3716
rect 47502 3676 47596 3716
rect 47636 3676 55372 3716
rect 55412 3676 55421 3716
rect 55555 3676 55564 3716
rect 55604 3676 58636 3716
rect 58676 3676 60652 3716
rect 60692 3676 60701 3716
rect 64003 3676 64012 3716
rect 64052 3676 70156 3716
rect 70196 3676 76012 3716
rect 76052 3676 76061 3716
rect 76771 3676 76780 3716
rect 76820 3676 82924 3716
rect 82964 3676 89164 3716
rect 89204 3676 89213 3716
rect 94252 3676 94636 3716
rect 94676 3676 94685 3716
rect 11980 3632 12020 3676
rect 21580 3632 21620 3676
rect 38083 3675 38141 3676
rect 47587 3675 47645 3676
rect 55363 3675 55421 3676
rect 32227 3632 32285 3633
rect 90691 3632 90749 3633
rect 94252 3632 94292 3676
rect 4387 3592 4396 3632
rect 4436 3592 10004 3632
rect 10147 3592 10156 3632
rect 10196 3592 10540 3632
rect 10580 3592 10924 3632
rect 10964 3592 11308 3632
rect 11348 3592 11692 3632
rect 11732 3592 11741 3632
rect 11980 3592 14476 3632
rect 14516 3592 14525 3632
rect 15235 3592 15244 3632
rect 15284 3592 21388 3632
rect 21428 3592 21437 3632
rect 21580 3592 23116 3632
rect 23156 3592 23165 3632
rect 32142 3592 32236 3632
rect 32276 3592 32285 3632
rect 32995 3592 33004 3632
rect 33044 3592 38380 3632
rect 38420 3592 38429 3632
rect 38563 3592 38572 3632
rect 38612 3592 40972 3632
rect 41012 3592 44620 3632
rect 44660 3592 44669 3632
rect 49123 3592 49132 3632
rect 49172 3592 57676 3632
rect 57716 3592 57725 3632
rect 57859 3592 57868 3632
rect 57908 3592 59116 3632
rect 59156 3592 67372 3632
rect 67412 3592 73324 3632
rect 73364 3592 73373 3632
rect 77644 3592 83788 3632
rect 83828 3592 89932 3632
rect 89972 3592 89981 3632
rect 90606 3592 90700 3632
rect 90740 3592 90749 3632
rect 92227 3592 92236 3632
rect 92276 3592 93100 3632
rect 93140 3592 93484 3632
rect 93524 3592 94252 3632
rect 94292 3592 94301 3632
rect 9571 3548 9629 3549
rect 9964 3548 10004 3592
rect 32227 3591 32285 3592
rect 41347 3548 41405 3549
rect 47875 3548 47933 3549
rect 69187 3548 69245 3549
rect 69763 3548 69821 3549
rect 71299 3548 71357 3549
rect 77644 3548 77684 3592
rect 90691 3591 90749 3592
rect 2092 3508 6320 3548
rect 6403 3508 6412 3548
rect 6452 3508 7276 3548
rect 7316 3508 7325 3548
rect 9486 3508 9580 3548
rect 9620 3508 9629 3548
rect 9955 3508 9964 3548
rect 10004 3508 13172 3548
rect 13219 3508 13228 3548
rect 13268 3508 13612 3548
rect 13652 3508 13996 3548
rect 14036 3508 14284 3548
rect 14324 3508 14668 3548
rect 14708 3508 15052 3548
rect 15092 3508 15436 3548
rect 15476 3508 15820 3548
rect 15860 3508 16204 3548
rect 16244 3508 16588 3548
rect 16628 3508 16972 3548
rect 17012 3508 17356 3548
rect 17396 3508 17780 3548
rect 17923 3508 17932 3548
rect 17972 3508 19372 3548
rect 19412 3508 19421 3548
rect 20707 3508 20716 3548
rect 20756 3508 26956 3548
rect 26996 3508 27005 3548
rect 28387 3508 28396 3548
rect 28436 3508 34156 3548
rect 34196 3508 40492 3548
rect 40532 3508 40541 3548
rect 41262 3508 41356 3548
rect 41396 3508 41405 3548
rect 43939 3508 43948 3548
rect 43988 3508 44428 3548
rect 44468 3508 44812 3548
rect 44852 3508 45196 3548
rect 45236 3508 45580 3548
rect 45620 3508 45964 3548
rect 46004 3508 46348 3548
rect 46388 3508 46640 3548
rect 47203 3508 47212 3548
rect 47252 3508 47884 3548
rect 47924 3508 48268 3548
rect 48308 3508 48317 3548
rect 48739 3508 48748 3548
rect 48788 3508 51148 3548
rect 51188 3508 52780 3548
rect 52820 3508 53260 3548
rect 53300 3508 53309 3548
rect 55420 3508 65452 3548
rect 65492 3508 65501 3548
rect 65635 3508 65644 3548
rect 65684 3508 66028 3548
rect 66068 3508 66316 3548
rect 66356 3508 66836 3548
rect 68611 3508 68620 3548
rect 68660 3508 69196 3548
rect 69236 3508 69245 3548
rect 69678 3508 69772 3548
rect 69812 3508 69821 3548
rect 71214 3508 71308 3548
rect 71348 3508 71357 3548
rect 71683 3508 71692 3548
rect 71732 3508 77644 3548
rect 77684 3508 77693 3548
rect 77923 3508 77932 3548
rect 77972 3508 84172 3548
rect 84212 3508 84221 3548
rect 87619 3508 87628 3548
rect 87668 3508 93332 3548
rect 94627 3508 94636 3548
rect 94676 3508 95020 3548
rect 95060 3508 95308 3548
rect 95348 3508 95692 3548
rect 95732 3508 96172 3548
rect 96212 3508 96556 3548
rect 96596 3508 96605 3548
rect 2092 3464 2132 3508
rect 5923 3464 5981 3465
rect 2083 3424 2092 3464
rect 2132 3424 2141 3464
rect 3715 3424 3724 3464
rect 3764 3424 4204 3464
rect 4244 3424 4588 3464
rect 4628 3424 4972 3464
rect 5012 3424 5021 3464
rect 5155 3424 5164 3464
rect 5204 3424 5213 3464
rect 5838 3424 5932 3464
rect 5972 3424 5981 3464
rect 6280 3464 6320 3508
rect 9571 3507 9629 3508
rect 6883 3464 6941 3465
rect 11107 3464 11165 3465
rect 11491 3464 11549 3465
rect 13027 3464 13085 3465
rect 6280 3424 6700 3464
rect 6740 3424 6749 3464
rect 6798 3424 6892 3464
rect 6932 3424 6941 3464
rect 7075 3424 7084 3464
rect 7124 3424 7468 3464
rect 7508 3424 7852 3464
rect 7892 3424 8236 3464
rect 8276 3424 8620 3464
rect 8660 3424 9004 3464
rect 9044 3424 9388 3464
rect 9428 3424 9772 3464
rect 9812 3424 10156 3464
rect 10196 3424 10205 3464
rect 11022 3424 11116 3464
rect 11156 3424 11165 3464
rect 11406 3424 11500 3464
rect 11540 3424 11549 3464
rect 11683 3424 11692 3464
rect 11732 3424 12076 3464
rect 12116 3424 12125 3464
rect 12942 3424 13036 3464
rect 13076 3424 13085 3464
rect 13132 3464 13172 3508
rect 17155 3464 17213 3465
rect 17539 3464 17597 3465
rect 17740 3464 17780 3508
rect 41347 3507 41405 3508
rect 18691 3464 18749 3465
rect 19939 3464 19997 3465
rect 23779 3464 23837 3465
rect 25315 3464 25373 3465
rect 29827 3464 29885 3465
rect 36835 3464 36893 3465
rect 46600 3464 46640 3508
rect 47875 3507 47933 3508
rect 50371 3464 50429 3465
rect 55420 3464 55460 3508
rect 65644 3464 65684 3508
rect 13132 3424 16012 3464
rect 16052 3424 16061 3464
rect 17070 3424 17164 3464
rect 17204 3424 17213 3464
rect 17454 3424 17548 3464
rect 17588 3424 17597 3464
rect 17731 3424 17740 3464
rect 17780 3424 18124 3464
rect 18164 3424 18508 3464
rect 18548 3424 18557 3464
rect 18691 3424 18700 3464
rect 18740 3424 18834 3464
rect 19854 3424 19948 3464
rect 19988 3424 19997 3464
rect 20140 3424 20149 3464
rect 20189 3424 20908 3464
rect 20948 3424 21292 3464
rect 21332 3424 21676 3464
rect 21716 3424 22060 3464
rect 22100 3424 22540 3464
rect 22580 3424 22924 3464
rect 22964 3424 23596 3464
rect 23636 3424 23645 3464
rect 23694 3424 23788 3464
rect 23828 3424 23837 3464
rect 25230 3424 25324 3464
rect 25364 3424 25373 3464
rect 25507 3424 25516 3464
rect 25556 3424 25900 3464
rect 25940 3424 26284 3464
rect 26324 3424 26764 3464
rect 26804 3424 27148 3464
rect 27188 3424 27820 3464
rect 27860 3424 28628 3464
rect 29742 3424 29836 3464
rect 29876 3424 29885 3464
rect 30211 3424 30220 3464
rect 30260 3424 30548 3464
rect 31459 3424 31468 3464
rect 31508 3424 31660 3464
rect 31700 3424 32044 3464
rect 32084 3424 32428 3464
rect 32468 3424 32812 3464
rect 32852 3424 33196 3464
rect 33236 3424 33580 3464
rect 33620 3424 33964 3464
rect 34004 3424 34348 3464
rect 34388 3424 34732 3464
rect 34772 3424 35116 3464
rect 35156 3424 35500 3464
rect 35540 3424 35884 3464
rect 35924 3424 36268 3464
rect 36308 3424 36652 3464
rect 36692 3424 36701 3464
rect 36835 3424 36844 3464
rect 36884 3424 36978 3464
rect 37507 3424 37516 3464
rect 37556 3424 37708 3464
rect 37748 3424 38476 3464
rect 38516 3424 38860 3464
rect 38900 3424 39244 3464
rect 39284 3424 39628 3464
rect 39668 3424 40012 3464
rect 40052 3424 40300 3464
rect 40340 3424 40780 3464
rect 40820 3424 41164 3464
rect 41204 3424 41644 3464
rect 41684 3424 41932 3464
rect 41972 3424 41981 3464
rect 42028 3424 45388 3464
rect 45428 3424 46444 3464
rect 46484 3424 46493 3464
rect 46600 3424 47020 3464
rect 47060 3424 47404 3464
rect 47444 3424 47788 3464
rect 47828 3424 47837 3464
rect 50083 3424 50092 3464
rect 50132 3424 50380 3464
rect 50420 3424 50668 3464
rect 50708 3424 50717 3464
rect 52003 3424 52012 3464
rect 52052 3424 55460 3464
rect 56131 3424 56140 3464
rect 56180 3424 56620 3464
rect 56660 3424 57100 3464
rect 57140 3424 57149 3464
rect 57955 3424 57964 3464
rect 58004 3424 58348 3464
rect 58388 3424 58397 3464
rect 58915 3424 58924 3464
rect 58964 3424 59308 3464
rect 59348 3424 59357 3464
rect 63139 3424 63148 3464
rect 63188 3424 63436 3464
rect 63476 3424 63820 3464
rect 63860 3424 64204 3464
rect 64244 3424 64588 3464
rect 64628 3424 65260 3464
rect 65300 3424 65684 3464
rect 65827 3464 65885 3465
rect 66211 3464 66269 3465
rect 66796 3464 66836 3508
rect 69187 3507 69245 3508
rect 69763 3507 69821 3508
rect 71299 3507 71357 3508
rect 72835 3464 72893 3465
rect 79171 3464 79229 3465
rect 80323 3464 80381 3465
rect 84547 3464 84605 3465
rect 92803 3464 92861 3465
rect 93292 3464 93332 3508
rect 65827 3424 65836 3464
rect 65876 3424 65970 3464
rect 66126 3424 66220 3464
rect 66260 3424 66269 3464
rect 66787 3424 66796 3464
rect 66836 3424 67180 3464
rect 67220 3424 67229 3464
rect 68803 3424 68812 3464
rect 68852 3424 69196 3464
rect 69236 3424 69580 3464
rect 69620 3424 69964 3464
rect 70004 3424 70348 3464
rect 70388 3424 70732 3464
rect 70772 3424 71116 3464
rect 71156 3424 71500 3464
rect 71540 3424 71884 3464
rect 71924 3424 72268 3464
rect 72308 3424 72652 3464
rect 72692 3424 72701 3464
rect 72750 3424 72844 3464
rect 72884 3424 72893 3464
rect 75139 3424 75148 3464
rect 75188 3424 75532 3464
rect 75572 3424 75820 3464
rect 75860 3424 76204 3464
rect 76244 3424 76588 3464
rect 76628 3424 76972 3464
rect 77012 3424 77452 3464
rect 77492 3424 78124 3464
rect 78164 3424 78508 3464
rect 78548 3424 78988 3464
rect 79028 3424 79037 3464
rect 79086 3424 79180 3464
rect 79220 3424 79229 3464
rect 80238 3424 80332 3464
rect 80372 3424 80381 3464
rect 81283 3424 81292 3464
rect 81332 3424 81676 3464
rect 81716 3424 82348 3464
rect 82388 3424 82732 3464
rect 82772 3424 83116 3464
rect 83156 3424 83596 3464
rect 83636 3424 83980 3464
rect 84020 3424 84364 3464
rect 84404 3424 84413 3464
rect 84462 3424 84556 3464
rect 84596 3424 84605 3464
rect 87043 3424 87052 3464
rect 87092 3424 87436 3464
rect 87476 3424 87820 3464
rect 87860 3424 88204 3464
rect 88244 3424 88588 3464
rect 88628 3424 88972 3464
rect 89012 3424 89356 3464
rect 89396 3424 89740 3464
rect 89780 3424 90124 3464
rect 90164 3424 90508 3464
rect 90548 3424 90892 3464
rect 90932 3424 91276 3464
rect 91316 3424 91660 3464
rect 91700 3424 92044 3464
rect 92084 3424 92428 3464
rect 92468 3424 92620 3464
rect 92660 3424 92669 3464
rect 92803 3424 92812 3464
rect 92852 3424 92946 3464
rect 93283 3424 93292 3464
rect 93332 3424 93341 3464
rect 94051 3424 94060 3464
rect 94100 3424 94109 3464
rect 94156 3424 94828 3464
rect 94868 3424 94877 3464
rect 5164 3380 5204 3424
rect 5923 3423 5981 3424
rect 6883 3423 6941 3424
rect 11107 3423 11165 3424
rect 11491 3423 11549 3424
rect 13027 3423 13085 3424
rect 16012 3380 16052 3424
rect 17155 3423 17213 3424
rect 17539 3423 17597 3424
rect 18691 3423 18749 3424
rect 19939 3423 19997 3424
rect 23779 3423 23837 3424
rect 25315 3423 25373 3424
rect 28588 3380 28628 3424
rect 29827 3423 29885 3424
rect 30508 3380 30548 3424
rect 36835 3423 36893 3424
rect 42028 3380 42068 3424
rect 50371 3423 50429 3424
rect 65827 3423 65885 3424
rect 66211 3423 66269 3424
rect 54307 3380 54365 3381
rect 64675 3380 64733 3381
rect 72451 3380 72509 3381
rect 5164 3340 10732 3380
rect 10772 3340 15956 3380
rect 16012 3340 22348 3380
rect 22388 3340 28396 3380
rect 28436 3340 28445 3380
rect 28579 3340 28588 3380
rect 28628 3340 28972 3380
rect 29012 3340 29356 3380
rect 29396 3340 29644 3380
rect 29684 3340 30028 3380
rect 30068 3340 30412 3380
rect 30452 3340 30461 3380
rect 30508 3340 36076 3380
rect 36116 3340 36125 3380
rect 38371 3340 38380 3380
rect 38420 3340 38429 3380
rect 39043 3340 39052 3380
rect 39092 3340 42068 3380
rect 42115 3340 42124 3380
rect 42164 3340 48076 3380
rect 48116 3340 48125 3380
rect 50275 3340 50284 3380
rect 50324 3340 50333 3380
rect 53923 3340 53932 3380
rect 53972 3340 54316 3380
rect 54356 3340 54365 3380
rect 56899 3340 56908 3380
rect 56948 3340 56957 3380
rect 58243 3340 58252 3380
rect 58292 3340 58301 3380
rect 58627 3340 58636 3380
rect 58676 3340 59116 3380
rect 59156 3340 59165 3380
rect 64675 3340 64684 3380
rect 64724 3340 64780 3380
rect 64820 3340 64829 3380
rect 65443 3340 65452 3380
rect 65492 3340 71692 3380
rect 71732 3340 71741 3380
rect 72366 3340 72460 3380
rect 72500 3340 72509 3380
rect 72652 3380 72692 3424
rect 72835 3423 72893 3424
rect 79171 3423 79229 3424
rect 80323 3423 80381 3424
rect 84547 3423 84605 3424
rect 92803 3423 92861 3424
rect 94060 3380 94100 3424
rect 72652 3340 73036 3380
rect 73076 3340 73085 3380
rect 76003 3340 76012 3380
rect 76052 3340 82156 3380
rect 82196 3340 88396 3380
rect 88436 3340 94100 3380
rect 15811 3296 15869 3297
rect 2659 3256 2668 3296
rect 2708 3256 8428 3296
rect 8468 3256 8477 3296
rect 10339 3256 10348 3296
rect 10388 3256 11692 3296
rect 11732 3256 11741 3296
rect 11788 3256 12268 3296
rect 12308 3256 12317 3296
rect 15726 3256 15820 3296
rect 15860 3256 15869 3296
rect 15916 3296 15956 3340
rect 30508 3296 30548 3340
rect 15916 3256 16780 3296
rect 16820 3256 16829 3296
rect 20140 3256 24172 3296
rect 24212 3256 30548 3296
rect 38380 3296 38420 3340
rect 50284 3296 50324 3340
rect 54307 3339 54365 3340
rect 56908 3296 56948 3340
rect 38380 3256 39436 3296
rect 39476 3256 39485 3296
rect 40483 3256 40492 3296
rect 40532 3256 46828 3296
rect 46868 3256 49268 3296
rect 50284 3256 50764 3296
rect 50804 3256 56620 3296
rect 56660 3256 56948 3296
rect 58252 3296 58292 3340
rect 64675 3339 64733 3340
rect 72451 3339 72509 3340
rect 66979 3296 67037 3297
rect 94156 3296 94196 3424
rect 94339 3340 94348 3380
rect 94388 3340 98188 3380
rect 98228 3340 98237 3380
rect 58252 3256 58540 3296
rect 58580 3256 58589 3296
rect 63331 3256 63340 3296
rect 63380 3256 63389 3296
rect 66894 3256 66988 3296
rect 67028 3256 67037 3296
rect 67363 3256 67372 3296
rect 67412 3256 70540 3296
rect 70580 3256 76396 3296
rect 76436 3256 76445 3296
rect 78979 3256 78988 3296
rect 79028 3256 79372 3296
rect 79412 3256 79756 3296
rect 79796 3256 80140 3296
rect 80180 3256 80189 3296
rect 81475 3256 81484 3296
rect 81524 3256 87628 3296
rect 87668 3256 87677 3296
rect 89155 3256 89164 3296
rect 89204 3256 94196 3296
rect 4195 3212 4253 3213
rect 10348 3212 10388 3256
rect 4195 3172 4204 3212
rect 4244 3172 4684 3212
rect 4724 3172 4733 3212
rect 4867 3172 4876 3212
rect 4916 3172 10388 3212
rect 4195 3171 4253 3172
rect 11788 3128 11828 3256
rect 15811 3255 15869 3256
rect 20140 3212 20180 3256
rect 31747 3212 31805 3213
rect 11875 3172 11884 3212
rect 11924 3172 17932 3212
rect 17972 3172 17981 3212
rect 18307 3172 18316 3212
rect 18356 3172 18836 3212
rect 19363 3172 19372 3212
rect 19412 3172 20180 3212
rect 23587 3172 23596 3212
rect 23636 3172 23980 3212
rect 24020 3172 24364 3212
rect 24404 3172 24652 3212
rect 24692 3172 24701 3212
rect 31662 3172 31756 3212
rect 31796 3172 31805 3212
rect 1603 3088 1612 3128
rect 1652 3088 6412 3128
rect 6452 3088 6461 3128
rect 6787 3088 6796 3128
rect 6836 3088 11828 3128
rect 11884 3044 11924 3172
rect 18316 3128 18356 3172
rect 12259 3088 12268 3128
rect 12308 3088 18356 3128
rect 18796 3044 18836 3172
rect 31747 3171 31805 3172
rect 34339 3212 34397 3213
rect 38083 3212 38141 3213
rect 49228 3212 49268 3256
rect 55075 3212 55133 3213
rect 34339 3172 34348 3212
rect 34388 3172 34444 3212
rect 34484 3172 34493 3212
rect 38083 3172 38092 3212
rect 38132 3172 39820 3212
rect 39860 3172 41836 3212
rect 41876 3172 41885 3212
rect 42019 3172 42028 3212
rect 42068 3172 42604 3212
rect 42644 3172 42653 3212
rect 43171 3172 43180 3212
rect 43220 3172 49132 3212
rect 49172 3172 49181 3212
rect 49228 3172 52012 3212
rect 52052 3172 52061 3212
rect 53347 3172 53356 3212
rect 53396 3172 54220 3212
rect 54260 3172 54269 3212
rect 54979 3172 54988 3212
rect 55028 3172 55084 3212
rect 55124 3172 55133 3212
rect 34339 3171 34397 3172
rect 38083 3171 38141 3172
rect 55075 3171 55133 3172
rect 41923 3128 41981 3129
rect 63340 3128 63380 3256
rect 66979 3255 67037 3256
rect 65347 3212 65405 3213
rect 65262 3172 65356 3212
rect 65396 3172 65405 3212
rect 66988 3212 67028 3255
rect 72931 3212 72989 3213
rect 83779 3212 83837 3213
rect 66988 3172 72940 3212
rect 72980 3172 72989 3212
rect 73699 3172 73708 3212
rect 73748 3172 79948 3212
rect 79988 3172 79997 3212
rect 80227 3172 80236 3212
rect 80276 3172 80620 3212
rect 80660 3172 80669 3212
rect 83683 3172 83692 3212
rect 83732 3172 83788 3212
rect 83828 3172 83837 3212
rect 89923 3172 89932 3212
rect 89972 3172 95500 3212
rect 95540 3172 95549 3212
rect 65347 3171 65405 3172
rect 72931 3171 72989 3172
rect 83779 3171 83837 3172
rect 18979 3088 18988 3128
rect 19028 3088 21100 3128
rect 21140 3088 21149 3128
rect 26083 3088 26092 3128
rect 26132 3088 31564 3128
rect 31604 3088 31613 3128
rect 39427 3088 39436 3128
rect 39476 3088 41932 3128
rect 41972 3088 41981 3128
rect 42115 3088 42124 3128
rect 42164 3088 42173 3128
rect 44611 3088 44620 3128
rect 44660 3088 69388 3128
rect 69428 3088 69437 3128
rect 72451 3088 72460 3128
rect 72500 3088 78220 3128
rect 78260 3088 78269 3128
rect 81091 3088 81100 3128
rect 81140 3088 87244 3128
rect 87284 3088 92908 3128
rect 92948 3088 92957 3128
rect 93004 3088 95980 3128
rect 96020 3088 96029 3128
rect 41923 3087 41981 3088
rect 35299 3044 35357 3045
rect 42124 3044 42164 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 4963 3004 4972 3044
rect 5012 3004 5740 3044
rect 5780 3004 5789 3044
rect 6307 3004 6316 3044
rect 6356 3004 11924 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 18796 3004 24556 3044
rect 24596 3004 24605 3044
rect 26947 3004 26956 3044
rect 26996 3004 32620 3044
rect 32660 3004 32669 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 35214 3004 35308 3044
rect 35348 3004 35357 3044
rect 36067 3004 36076 3044
rect 36116 3004 42164 3044
rect 42211 3044 42269 3045
rect 46147 3044 46205 3045
rect 93004 3044 93044 3088
rect 42211 3004 42220 3044
rect 42260 3004 45772 3044
rect 45812 3004 45821 3044
rect 46062 3004 46156 3044
rect 46196 3004 46205 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 50371 3004 50380 3044
rect 50420 3004 50572 3044
rect 50612 3004 50621 3044
rect 54499 3004 54508 3044
rect 54548 3004 55372 3044
rect 55412 3004 55421 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 64387 3004 64396 3044
rect 64436 3004 67372 3044
rect 67412 3004 67421 3044
rect 70915 3004 70924 3044
rect 70964 3004 76684 3044
rect 76724 3004 76733 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 90307 3004 90316 3044
rect 90356 3004 93044 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 35299 3003 35357 3004
rect 42211 3003 42269 3004
rect 46147 3003 46205 3004
rect 46156 2960 46196 3003
rect 6691 2920 6700 2960
rect 6740 2920 7660 2960
rect 7700 2920 13804 2960
rect 13844 2920 13853 2960
rect 16396 2920 22732 2960
rect 22772 2920 28780 2960
rect 28820 2920 34540 2960
rect 34580 2920 40972 2960
rect 41012 2920 41021 2960
rect 41827 2920 41836 2960
rect 41876 2920 46196 2960
rect 54979 2960 55037 2961
rect 65827 2960 65885 2961
rect 54979 2920 54988 2960
rect 55028 2920 55180 2960
rect 55220 2920 55229 2960
rect 57667 2920 57676 2960
rect 57716 2920 64204 2960
rect 64244 2920 64253 2960
rect 65827 2920 65836 2960
rect 65876 2920 72076 2960
rect 72116 2920 72125 2960
rect 76387 2920 76396 2960
rect 76436 2920 82540 2960
rect 82580 2920 88780 2960
rect 88820 2920 88829 2960
rect 92227 2920 92236 2960
rect 92276 2920 98092 2960
rect 98132 2920 98141 2960
rect 16396 2876 16436 2920
rect 54979 2919 55037 2920
rect 65827 2919 65885 2920
rect 20131 2876 20189 2877
rect 44035 2876 44093 2877
rect 44995 2876 45053 2877
rect 91459 2876 91517 2877
rect 11683 2836 11692 2876
rect 11732 2836 16396 2876
rect 16436 2836 16445 2876
rect 20035 2836 20044 2876
rect 20084 2836 20140 2876
rect 20180 2836 20189 2876
rect 24547 2836 24556 2876
rect 24596 2836 30700 2876
rect 30740 2836 36460 2876
rect 36500 2836 36509 2876
rect 37987 2836 37996 2876
rect 38036 2836 38284 2876
rect 38324 2836 38333 2876
rect 43950 2836 44044 2876
rect 44084 2836 45004 2876
rect 45044 2836 45053 2876
rect 48067 2836 48076 2876
rect 48116 2836 48844 2876
rect 48884 2836 57964 2876
rect 58004 2836 58013 2876
rect 60643 2836 60652 2876
rect 60692 2836 60940 2876
rect 60980 2836 60989 2876
rect 69379 2836 69388 2876
rect 69428 2836 75340 2876
rect 75380 2836 75389 2876
rect 84163 2836 84172 2876
rect 84212 2836 90316 2876
rect 90356 2836 90365 2876
rect 91374 2836 91468 2876
rect 91508 2836 91517 2876
rect 20131 2835 20189 2836
rect 44035 2835 44093 2836
rect 44995 2835 45053 2836
rect 91459 2835 91517 2836
rect 20035 2792 20093 2793
rect 54883 2792 54941 2793
rect 64675 2792 64733 2793
rect 74755 2792 74813 2793
rect 84739 2792 84797 2793
rect 84931 2792 84989 2793
rect 92236 2792 92276 2920
rect 92803 2876 92861 2877
rect 92803 2836 92812 2876
rect 92852 2836 94348 2876
rect 94388 2836 94397 2876
rect 92803 2835 92861 2836
rect 3139 2752 3148 2792
rect 3188 2752 8812 2792
rect 8852 2752 14860 2792
rect 14900 2752 18988 2792
rect 19028 2752 19037 2792
rect 19843 2752 19852 2792
rect 19892 2752 20044 2792
rect 20084 2752 20093 2792
rect 40963 2752 40972 2792
rect 41012 2752 47212 2792
rect 47252 2752 47261 2792
rect 47779 2752 47788 2792
rect 47828 2752 48268 2792
rect 48308 2752 48652 2792
rect 48692 2752 48940 2792
rect 48980 2752 49132 2792
rect 49172 2752 49181 2792
rect 54883 2752 54892 2792
rect 54932 2752 55276 2792
rect 55316 2752 55564 2792
rect 55604 2752 55613 2792
rect 55747 2752 55756 2792
rect 55796 2752 56044 2792
rect 56084 2752 58252 2792
rect 58292 2752 61420 2792
rect 61460 2752 61804 2792
rect 61844 2752 61853 2792
rect 62851 2752 62860 2792
rect 62900 2752 63340 2792
rect 63380 2752 63389 2792
rect 64675 2752 64684 2792
rect 64724 2752 70924 2792
rect 70964 2752 70973 2792
rect 74670 2752 74764 2792
rect 74804 2752 74813 2792
rect 20035 2751 20093 2752
rect 54883 2751 54941 2752
rect 64675 2751 64733 2752
rect 74755 2751 74813 2752
rect 78028 2752 79564 2792
rect 79604 2752 84748 2792
rect 84788 2752 84797 2792
rect 84846 2752 84940 2792
rect 84980 2752 84989 2792
rect 14275 2708 14333 2709
rect 48067 2708 48125 2709
rect 61315 2708 61373 2709
rect 72931 2708 72989 2709
rect 3532 2668 9196 2708
rect 9236 2668 9245 2708
rect 14190 2668 14284 2708
rect 14324 2668 14333 2708
rect 14467 2668 14476 2708
rect 14516 2668 20716 2708
rect 20756 2668 20765 2708
rect 23107 2668 23116 2708
rect 23156 2668 29164 2708
rect 29204 2668 34924 2708
rect 34964 2668 41356 2708
rect 41396 2668 41405 2708
rect 41635 2668 41644 2708
rect 41684 2668 42028 2708
rect 42068 2668 42796 2708
rect 42836 2668 42845 2708
rect 47982 2668 48076 2708
rect 48116 2668 48125 2708
rect 48355 2668 48364 2708
rect 48404 2668 48413 2708
rect 49132 2668 55220 2708
rect 61230 2668 61324 2708
rect 61364 2668 61373 2708
rect 2275 2624 2333 2625
rect 3532 2624 3572 2668
rect 14275 2667 14333 2668
rect 48067 2667 48125 2668
rect 3907 2624 3965 2625
rect 7171 2624 7229 2625
rect 8035 2624 8093 2625
rect 12739 2624 12797 2625
rect 20035 2624 20093 2625
rect 20419 2624 20477 2625
rect 21859 2624 21917 2625
rect 23395 2624 23453 2625
rect 26563 2624 26621 2625
rect 28099 2624 28157 2625
rect 29539 2624 29597 2625
rect 30883 2624 30941 2625
rect 31651 2624 31709 2625
rect 33763 2624 33821 2625
rect 38755 2624 38813 2625
rect 40195 2624 40253 2625
rect 41827 2624 41885 2625
rect 42211 2624 42269 2625
rect 42979 2624 43037 2625
rect 46531 2624 46589 2625
rect 2190 2584 2284 2624
rect 2324 2584 2333 2624
rect 3523 2584 3532 2624
rect 3572 2584 3581 2624
rect 3822 2584 3916 2624
rect 3956 2584 3965 2624
rect 5347 2584 5356 2624
rect 5396 2584 5740 2624
rect 5780 2584 6124 2624
rect 6164 2584 6604 2624
rect 6644 2584 6988 2624
rect 7028 2584 7037 2624
rect 7086 2584 7180 2624
rect 7220 2584 7229 2624
rect 7950 2584 8044 2624
rect 8084 2584 8093 2624
rect 12654 2584 12748 2624
rect 12788 2584 12797 2624
rect 19459 2584 19468 2624
rect 19508 2584 19660 2624
rect 19700 2584 19988 2624
rect 2275 2583 2333 2584
rect 3907 2583 3965 2584
rect 7171 2583 7229 2584
rect 8035 2583 8093 2584
rect 12739 2583 12797 2584
rect 6595 2540 6653 2541
rect 19948 2540 19988 2584
rect 20035 2584 20044 2624
rect 20084 2584 20236 2624
rect 20276 2584 20285 2624
rect 20334 2584 20428 2624
rect 20468 2584 20477 2624
rect 21774 2584 21868 2624
rect 21908 2584 21917 2624
rect 23310 2584 23404 2624
rect 23444 2584 23453 2624
rect 26478 2584 26572 2624
rect 26612 2584 26621 2624
rect 28014 2584 28108 2624
rect 28148 2584 28157 2624
rect 29454 2584 29548 2624
rect 29588 2584 29597 2624
rect 29731 2584 29740 2624
rect 29780 2584 30700 2624
rect 30740 2584 30749 2624
rect 30798 2584 30892 2624
rect 30932 2584 30941 2624
rect 31566 2584 31660 2624
rect 31700 2584 32780 2624
rect 33678 2584 33772 2624
rect 33812 2584 33821 2624
rect 37795 2584 37804 2624
rect 37844 2584 38572 2624
rect 38612 2584 38621 2624
rect 38755 2584 38764 2624
rect 38804 2584 38898 2624
rect 40110 2584 40204 2624
rect 40244 2584 40253 2624
rect 41742 2584 41836 2624
rect 41876 2584 41885 2624
rect 42126 2584 42220 2624
rect 42260 2584 42269 2624
rect 42894 2584 42988 2624
rect 43028 2584 43037 2624
rect 46446 2584 46540 2624
rect 46580 2584 46589 2624
rect 20035 2583 20093 2584
rect 20419 2583 20477 2584
rect 21859 2583 21917 2584
rect 23395 2583 23453 2584
rect 26563 2583 26621 2584
rect 28099 2583 28157 2584
rect 29539 2583 29597 2584
rect 30883 2583 30941 2584
rect 31651 2583 31709 2584
rect 2500 2500 2860 2540
rect 2900 2500 3244 2540
rect 3284 2500 3628 2540
rect 3668 2500 3677 2540
rect 6595 2500 6604 2540
rect 6644 2500 7084 2540
rect 7124 2500 7133 2540
rect 19948 2500 20180 2540
rect 2500 2456 2540 2500
rect 6595 2499 6653 2500
rect 19939 2456 19997 2457
rect 1795 2416 1804 2456
rect 1844 2416 2092 2456
rect 2132 2416 2476 2456
rect 2516 2416 2540 2456
rect 6403 2416 6412 2456
rect 6452 2416 13420 2456
rect 13460 2416 13469 2456
rect 13795 2416 13804 2456
rect 13844 2416 19948 2456
rect 19988 2416 19997 2456
rect 20140 2456 20180 2500
rect 20140 2416 25708 2456
rect 25748 2416 29000 2456
rect 13420 2288 13460 2416
rect 19939 2415 19997 2416
rect 20419 2372 20477 2373
rect 14275 2332 14284 2372
rect 14324 2332 20428 2372
rect 20468 2332 20477 2372
rect 20419 2331 20477 2332
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 5539 2248 5548 2288
rect 5588 2248 11116 2288
rect 11156 2248 11165 2288
rect 13420 2248 19372 2288
rect 19412 2248 19421 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 19939 2204 19997 2205
rect 28960 2204 29000 2416
rect 32740 2372 32780 2584
rect 33763 2583 33821 2584
rect 38188 2540 38228 2584
rect 38755 2583 38813 2584
rect 40195 2583 40253 2584
rect 41827 2583 41885 2584
rect 42211 2583 42269 2584
rect 42979 2583 43037 2584
rect 46531 2583 46589 2584
rect 46636 2584 48212 2624
rect 38179 2500 38188 2540
rect 38228 2500 38268 2540
rect 38764 2456 38804 2583
rect 41923 2540 41981 2541
rect 42307 2540 42365 2541
rect 46636 2540 46676 2584
rect 41731 2500 41740 2540
rect 41780 2500 41932 2540
rect 41972 2500 41981 2540
rect 42222 2500 42316 2540
rect 42356 2500 42365 2540
rect 41923 2499 41981 2500
rect 42307 2499 42365 2500
rect 46600 2500 46676 2540
rect 46600 2456 46640 2500
rect 34819 2416 34828 2456
rect 34868 2416 35308 2456
rect 35348 2416 35357 2456
rect 35404 2416 38804 2456
rect 42019 2416 42028 2456
rect 42068 2416 42412 2456
rect 42452 2416 42461 2456
rect 44227 2416 44236 2456
rect 44276 2416 46640 2456
rect 48172 2456 48212 2584
rect 48364 2541 48404 2668
rect 48451 2624 48509 2625
rect 48451 2584 48460 2624
rect 48500 2584 48594 2624
rect 48451 2583 48509 2584
rect 48355 2540 48413 2541
rect 48355 2500 48364 2540
rect 48404 2500 48413 2540
rect 49132 2540 49172 2668
rect 49315 2624 49373 2625
rect 49230 2584 49324 2624
rect 49364 2584 49373 2624
rect 49315 2583 49373 2584
rect 54883 2624 54941 2625
rect 54883 2576 54892 2624
rect 54932 2584 55019 2624
rect 54932 2576 54941 2584
rect 55180 2540 55220 2668
rect 61315 2667 61373 2668
rect 61420 2668 61996 2708
rect 62036 2668 62045 2708
rect 63052 2668 69004 2708
rect 69044 2668 69053 2708
rect 72846 2668 72940 2708
rect 72980 2668 72989 2708
rect 73123 2668 73132 2708
rect 73172 2668 73516 2708
rect 73556 2668 73900 2708
rect 73940 2668 74092 2708
rect 74132 2668 74141 2708
rect 74947 2668 74956 2708
rect 74996 2668 75820 2708
rect 75860 2668 75869 2708
rect 58627 2624 58685 2625
rect 61420 2624 61460 2668
rect 61699 2624 61757 2625
rect 63052 2624 63092 2668
rect 72931 2667 72989 2668
rect 63523 2624 63581 2625
rect 64003 2624 64061 2625
rect 75619 2624 75677 2625
rect 55363 2584 55372 2624
rect 55412 2584 55756 2624
rect 55796 2584 56236 2624
rect 56276 2584 56285 2624
rect 58542 2584 58636 2624
rect 58676 2584 58924 2624
rect 58964 2584 58973 2624
rect 60451 2584 60460 2624
rect 60500 2584 60940 2624
rect 60980 2584 61420 2624
rect 61460 2584 61469 2624
rect 61614 2584 61708 2624
rect 61748 2584 61757 2624
rect 62957 2584 63052 2624
rect 63092 2584 63101 2624
rect 63438 2584 63532 2624
rect 63572 2584 64012 2624
rect 64052 2584 64061 2624
rect 64195 2584 64204 2624
rect 64244 2584 67372 2624
rect 67412 2584 73708 2624
rect 73748 2584 73757 2624
rect 75534 2584 75628 2624
rect 75668 2584 75677 2624
rect 58627 2583 58685 2584
rect 61699 2583 61757 2584
rect 49132 2500 49268 2540
rect 55180 2500 55604 2540
rect 48355 2499 48413 2500
rect 49228 2456 49268 2500
rect 55459 2456 55517 2457
rect 48172 2416 49268 2456
rect 49612 2416 55468 2456
rect 55508 2416 55517 2456
rect 55564 2456 55604 2500
rect 59107 2456 59165 2457
rect 55564 2416 55892 2456
rect 59022 2416 59116 2456
rect 59156 2416 59165 2456
rect 60547 2416 60556 2456
rect 60596 2416 61324 2456
rect 61364 2416 61373 2456
rect 35299 2372 35357 2373
rect 32740 2332 35308 2372
rect 35348 2332 35357 2372
rect 35299 2331 35357 2332
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 32227 2204 32285 2205
rect 35404 2204 35444 2416
rect 35587 2372 35645 2373
rect 35587 2332 35596 2372
rect 35636 2332 37612 2372
rect 37652 2332 37661 2372
rect 35587 2331 35645 2332
rect 36451 2248 36460 2288
rect 36500 2248 43180 2288
rect 43220 2248 43229 2288
rect 49612 2204 49652 2416
rect 55459 2415 55517 2416
rect 55852 2372 55892 2416
rect 59107 2415 59165 2416
rect 63052 2372 63092 2584
rect 63523 2583 63581 2584
rect 64003 2583 64061 2584
rect 75619 2583 75677 2584
rect 76867 2624 76925 2625
rect 76867 2584 76876 2624
rect 76916 2584 77260 2624
rect 77300 2584 77309 2624
rect 76867 2583 76925 2584
rect 74275 2540 74333 2541
rect 77251 2540 77309 2541
rect 66787 2500 66796 2540
rect 66836 2500 66845 2540
rect 73284 2500 73324 2540
rect 73364 2500 73373 2540
rect 74190 2500 74284 2540
rect 74324 2500 74333 2540
rect 77155 2500 77164 2540
rect 77204 2500 77260 2540
rect 77300 2500 77309 2540
rect 64291 2456 64349 2457
rect 66595 2456 66653 2457
rect 64291 2416 64300 2456
rect 64340 2416 66604 2456
rect 66644 2416 66653 2456
rect 66796 2456 66836 2500
rect 73324 2456 73364 2500
rect 74275 2499 74333 2500
rect 77251 2499 77309 2500
rect 78028 2456 78068 2752
rect 84739 2751 84797 2752
rect 84931 2751 84989 2752
rect 85036 2752 86092 2792
rect 86132 2752 92276 2792
rect 92332 2752 97516 2792
rect 97556 2752 97565 2792
rect 85036 2708 85076 2752
rect 85315 2708 85373 2709
rect 88003 2708 88061 2709
rect 92332 2708 92372 2752
rect 93667 2708 93725 2709
rect 79939 2668 79948 2708
rect 79988 2668 85076 2708
rect 85230 2668 85324 2708
rect 85364 2668 85373 2708
rect 85315 2667 85373 2668
rect 85516 2668 85900 2708
rect 85940 2668 86284 2708
rect 86324 2668 86333 2708
rect 87918 2668 88012 2708
rect 88052 2668 88061 2708
rect 78595 2624 78653 2625
rect 81475 2624 81533 2625
rect 83395 2624 83453 2625
rect 85516 2624 85556 2668
rect 88003 2667 88061 2668
rect 89356 2668 91852 2708
rect 91892 2668 92372 2708
rect 93582 2668 93676 2708
rect 93716 2668 93725 2708
rect 96547 2668 96556 2708
rect 96596 2668 96940 2708
rect 96980 2668 97324 2708
rect 97364 2668 97708 2708
rect 97748 2668 97900 2708
rect 97940 2668 97949 2708
rect 86467 2624 86525 2625
rect 78595 2584 78604 2624
rect 78644 2584 78796 2624
rect 78836 2584 78845 2624
rect 81475 2584 81484 2624
rect 81524 2584 81868 2624
rect 81908 2584 81917 2624
rect 83310 2584 83404 2624
rect 83444 2584 83453 2624
rect 84355 2584 84364 2624
rect 84404 2584 84748 2624
rect 84788 2584 85132 2624
rect 85172 2584 85516 2624
rect 85556 2584 85565 2624
rect 85699 2584 85708 2624
rect 85748 2584 85788 2624
rect 86382 2584 86476 2624
rect 86516 2584 86525 2624
rect 78595 2583 78653 2584
rect 81475 2583 81533 2584
rect 83395 2583 83453 2584
rect 85219 2540 85277 2541
rect 85134 2500 85228 2540
rect 85268 2500 85277 2540
rect 85219 2499 85277 2500
rect 84547 2456 84605 2457
rect 66796 2416 67564 2456
rect 67604 2416 67613 2456
rect 73324 2416 78068 2456
rect 78211 2416 78220 2456
rect 78260 2416 84556 2456
rect 84596 2416 84605 2456
rect 64291 2415 64349 2416
rect 66595 2415 66653 2416
rect 84547 2415 84605 2416
rect 84739 2456 84797 2457
rect 85708 2456 85748 2584
rect 86467 2583 86525 2584
rect 89356 2456 89396 2668
rect 93667 2667 93725 2668
rect 89539 2624 89597 2625
rect 95107 2624 95165 2625
rect 96355 2624 96413 2625
rect 96739 2624 96797 2625
rect 97123 2624 97181 2625
rect 89454 2584 89548 2624
rect 89588 2584 89597 2624
rect 92707 2584 92716 2624
rect 92756 2584 93100 2624
rect 93140 2584 93772 2624
rect 93812 2584 93821 2624
rect 95022 2584 95116 2624
rect 95156 2584 95165 2624
rect 96270 2584 96364 2624
rect 96404 2584 96413 2624
rect 96654 2584 96748 2624
rect 96788 2584 96797 2624
rect 97038 2584 97132 2624
rect 97172 2584 97181 2624
rect 89539 2583 89597 2584
rect 95107 2583 95165 2584
rect 96355 2583 96413 2584
rect 96739 2583 96797 2584
rect 97123 2583 97181 2584
rect 91075 2540 91133 2541
rect 97987 2540 98045 2541
rect 90990 2500 91084 2540
rect 91124 2500 91133 2540
rect 97603 2500 97612 2540
rect 97652 2500 97996 2540
rect 98036 2500 98045 2540
rect 91075 2499 91133 2500
rect 97987 2499 98045 2500
rect 84739 2416 84748 2456
rect 84788 2416 89396 2456
rect 92995 2416 93004 2456
rect 93044 2416 93484 2456
rect 93524 2416 93533 2456
rect 84739 2415 84797 2416
rect 66604 2372 66644 2415
rect 93859 2372 93917 2373
rect 50380 2332 55460 2372
rect 55852 2332 63092 2372
rect 66595 2332 66604 2372
rect 66644 2332 66684 2372
rect 75331 2332 75340 2372
rect 75380 2332 81484 2372
rect 81524 2332 81533 2372
rect 91075 2332 91084 2372
rect 91124 2332 93868 2372
rect 93908 2332 93917 2372
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 19939 2164 19948 2204
rect 19988 2164 26092 2204
rect 26132 2164 26141 2204
rect 28960 2164 31180 2204
rect 31220 2164 31229 2204
rect 32227 2164 32236 2204
rect 32276 2164 35444 2204
rect 35683 2164 35692 2204
rect 35732 2164 38092 2204
rect 38132 2164 38141 2204
rect 45475 2164 45484 2204
rect 45524 2164 49652 2204
rect 19939 2163 19997 2164
rect 32227 2163 32285 2164
rect 50380 2120 50420 2332
rect 55420 2288 55460 2332
rect 93859 2331 93917 2332
rect 55555 2288 55613 2289
rect 51811 2248 51820 2288
rect 51860 2248 52300 2288
rect 52340 2248 52876 2288
rect 52916 2248 53356 2288
rect 53396 2248 54316 2288
rect 54356 2248 54700 2288
rect 54740 2248 55276 2288
rect 55316 2248 55325 2288
rect 55420 2248 55508 2288
rect 55468 2204 55508 2248
rect 55555 2248 55564 2288
rect 55604 2248 64108 2288
rect 64148 2248 64157 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 55555 2247 55613 2248
rect 55468 2164 64396 2204
rect 64436 2164 64445 2204
rect 68995 2164 69004 2204
rect 69044 2164 74668 2204
rect 74708 2164 81100 2204
rect 81140 2164 81149 2204
rect 6979 2080 6988 2120
rect 7028 2080 12172 2120
rect 12212 2080 12221 2120
rect 31555 2080 31564 2120
rect 31604 2080 32852 2120
rect 6403 1996 6412 2036
rect 6452 1996 6796 2036
rect 6836 1996 7276 2036
rect 7316 1996 7325 2036
rect 6883 1952 6941 1953
rect 19363 1952 19421 1953
rect 24835 1952 24893 1953
rect 32812 1952 32852 2080
rect 35788 2080 38380 2120
rect 38420 2080 38429 2120
rect 45763 2080 45772 2120
rect 45812 2080 50420 2120
rect 56995 2080 57004 2120
rect 57044 2080 57484 2120
rect 57524 2080 58060 2120
rect 58100 2080 58109 2120
rect 58732 2080 59020 2120
rect 59060 2080 59069 2120
rect 35788 1952 35828 2080
rect 58435 2036 58493 2037
rect 42883 1996 42892 2036
rect 42932 1996 43468 2036
rect 43508 1996 43517 2036
rect 51043 1996 51052 2036
rect 51092 1996 51436 2036
rect 51476 1996 51485 2036
rect 52108 1996 57388 2036
rect 57428 1996 57868 2036
rect 57908 1996 57917 2036
rect 58350 1996 58444 2036
rect 58484 1996 58493 2036
rect 52108 1953 52148 1996
rect 58435 1995 58493 1996
rect 50371 1952 50429 1953
rect 51427 1952 51485 1953
rect 52099 1952 52157 1953
rect 58732 1952 58772 2080
rect 69187 2036 69245 2037
rect 62572 1996 69196 2036
rect 69236 1996 69245 2036
rect 62572 1953 62612 1996
rect 69187 1995 69245 1996
rect 62563 1952 62621 1953
rect 1507 1912 1516 1952
rect 1556 1912 6892 1952
rect 6932 1912 6941 1952
rect 19278 1912 19372 1952
rect 19412 1912 19421 1952
rect 19555 1912 19564 1952
rect 19604 1912 20044 1952
rect 20084 1912 20093 1952
rect 24750 1912 24844 1952
rect 24884 1912 24893 1952
rect 31939 1912 31948 1952
rect 31988 1912 32716 1952
rect 32756 1912 32765 1952
rect 32812 1912 35828 1952
rect 37603 1912 37612 1952
rect 37652 1912 43852 1952
rect 43892 1912 46252 1952
rect 46292 1912 50380 1952
rect 50420 1912 50429 1952
rect 51235 1912 51244 1952
rect 51284 1912 51436 1952
rect 51476 1912 51724 1952
rect 51764 1912 51773 1952
rect 51907 1912 51916 1952
rect 51956 1912 52108 1952
rect 52148 1912 52157 1952
rect 52963 1912 52972 1952
rect 53012 1912 53164 1952
rect 53204 1912 58732 1952
rect 58772 1912 58781 1952
rect 58915 1912 58924 1952
rect 58964 1912 59980 1952
rect 60020 1912 60460 1952
rect 60500 1912 60509 1952
rect 62478 1912 62572 1952
rect 62612 1912 62621 1952
rect 6883 1911 6941 1912
rect 19363 1911 19421 1912
rect 24835 1911 24893 1912
rect 50371 1911 50429 1912
rect 51427 1911 51485 1912
rect 52099 1911 52157 1912
rect 62563 1911 62621 1912
rect 64579 1952 64637 1953
rect 67843 1952 67901 1953
rect 64579 1912 64588 1952
rect 64628 1912 65068 1952
rect 65108 1912 65117 1952
rect 67758 1912 67852 1952
rect 67892 1912 67901 1952
rect 74755 1912 74764 1952
rect 74804 1912 80812 1952
rect 80852 1912 86764 1952
rect 86804 1912 92524 1952
rect 92564 1912 92573 1952
rect 64579 1911 64637 1912
rect 67843 1911 67901 1912
rect 37315 1868 37373 1869
rect 79939 1868 79997 1869
rect 26083 1828 26092 1868
rect 26132 1828 32140 1868
rect 32180 1828 37324 1868
rect 37364 1828 37373 1868
rect 51427 1828 51436 1868
rect 51476 1828 57196 1868
rect 57236 1828 57245 1868
rect 61891 1828 61900 1868
rect 61940 1828 62380 1868
rect 62420 1828 62429 1868
rect 79854 1828 79948 1868
rect 79988 1828 79997 1868
rect 37315 1827 37373 1828
rect 79939 1827 79997 1828
rect 32611 1744 32620 1784
rect 32660 1744 39052 1784
rect 39092 1744 39101 1784
rect 55363 1744 55372 1784
rect 55412 1744 60652 1784
rect 60692 1744 60701 1784
rect 55459 1700 55517 1701
rect 55939 1700 55997 1701
rect 64003 1700 64061 1701
rect 24739 1660 24748 1700
rect 24788 1660 25132 1700
rect 25172 1660 25181 1700
rect 31171 1660 31180 1700
rect 31220 1660 35692 1700
rect 35732 1660 35741 1700
rect 54019 1660 54028 1700
rect 54068 1660 54508 1700
rect 54548 1660 54557 1700
rect 55459 1660 55468 1700
rect 55508 1660 55564 1700
rect 55604 1660 55613 1700
rect 55843 1660 55852 1700
rect 55892 1660 55948 1700
rect 55988 1660 55997 1700
rect 56227 1660 56236 1700
rect 56276 1660 57004 1700
rect 57044 1660 57053 1700
rect 58723 1660 58732 1700
rect 58772 1660 59020 1700
rect 59060 1660 59069 1700
rect 59299 1660 59308 1700
rect 59348 1660 60268 1700
rect 60308 1660 60317 1700
rect 63918 1660 64012 1700
rect 64052 1660 64061 1700
rect 92611 1660 92620 1700
rect 92660 1660 93100 1700
rect 93140 1660 93149 1700
rect 55459 1659 55517 1660
rect 55939 1659 55997 1660
rect 64003 1659 64061 1660
rect 42307 1616 42365 1617
rect 55075 1616 55133 1617
rect 71299 1616 71357 1617
rect 79843 1616 79901 1617
rect 13027 1576 13036 1616
rect 13076 1576 18892 1616
rect 18932 1576 18941 1616
rect 31459 1576 31468 1616
rect 31508 1576 37804 1616
rect 37844 1576 42316 1616
rect 42356 1576 42365 1616
rect 50275 1576 50284 1616
rect 50324 1576 50668 1616
rect 50708 1576 50717 1616
rect 53731 1576 53740 1616
rect 53780 1576 54124 1616
rect 54164 1576 55084 1616
rect 55124 1576 59500 1616
rect 59540 1576 59549 1616
rect 68707 1576 68716 1616
rect 68756 1576 69100 1616
rect 69140 1576 69149 1616
rect 71299 1576 71308 1616
rect 71348 1576 77452 1616
rect 77492 1576 77501 1616
rect 79758 1576 79852 1616
rect 79892 1576 79901 1616
rect 80035 1576 80044 1616
rect 80084 1576 86092 1616
rect 86132 1576 86141 1616
rect 42307 1575 42365 1576
rect 55075 1575 55133 1576
rect 71299 1575 71357 1576
rect 79843 1575 79901 1576
rect 20419 1532 20477 1533
rect 23875 1532 23933 1533
rect 55459 1532 55517 1533
rect 70723 1532 70781 1533
rect 79747 1532 79805 1533
rect 94819 1532 94877 1533
rect 97219 1532 97277 1533
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 20334 1492 20428 1532
rect 20468 1492 20477 1532
rect 23683 1492 23692 1532
rect 23732 1492 23884 1532
rect 23924 1492 23933 1532
rect 28963 1492 28972 1532
rect 29012 1492 33243 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 35971 1492 35980 1532
rect 36020 1492 36748 1532
rect 36788 1492 36797 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 55267 1492 55276 1532
rect 55316 1492 55468 1532
rect 55508 1492 55517 1532
rect 20419 1491 20477 1492
rect 23875 1491 23933 1492
rect 6403 1448 6461 1449
rect 11203 1448 11261 1449
rect 32995 1448 33053 1449
rect 6403 1408 6412 1448
rect 6452 1408 6796 1448
rect 6836 1408 6845 1448
rect 11203 1408 11212 1448
rect 11252 1408 15956 1448
rect 19459 1408 19468 1448
rect 19508 1408 25516 1448
rect 25556 1408 25565 1448
rect 32515 1408 32524 1448
rect 32564 1408 33004 1448
rect 33044 1408 33053 1448
rect 33203 1448 33243 1492
rect 55459 1491 55517 1492
rect 55564 1492 60172 1532
rect 60212 1492 60221 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 70638 1492 70732 1532
rect 70772 1492 70781 1532
rect 70915 1492 70924 1532
rect 70964 1492 77068 1532
rect 77108 1492 77117 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 79662 1492 79756 1532
rect 79796 1492 85708 1532
rect 85748 1492 85757 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 94627 1492 94636 1532
rect 94676 1492 94828 1532
rect 94868 1492 94877 1532
rect 97027 1492 97036 1532
rect 97076 1492 97228 1532
rect 97268 1492 97277 1532
rect 35107 1448 35165 1449
rect 33203 1408 34924 1448
rect 34964 1408 35116 1448
rect 35156 1408 35165 1448
rect 6403 1407 6461 1408
rect 11203 1407 11261 1408
rect 5827 1364 5885 1365
rect 14275 1364 14333 1365
rect 5827 1324 5836 1364
rect 5876 1324 6220 1364
rect 6260 1324 6269 1364
rect 14190 1324 14284 1364
rect 14324 1324 14333 1364
rect 5827 1323 5885 1324
rect 14275 1323 14333 1324
rect 14380 1324 14612 1364
rect 4771 1280 4829 1281
rect 6211 1280 6269 1281
rect 14380 1280 14420 1324
rect 1027 1240 1036 1280
rect 1076 1240 1420 1280
rect 1460 1240 1844 1280
rect 1804 1196 1844 1240
rect 3340 1240 3724 1280
rect 3764 1240 4108 1280
rect 4148 1240 4532 1280
rect 3340 1196 3380 1240
rect 4492 1196 4532 1240
rect 4771 1240 4780 1280
rect 4820 1240 5068 1280
rect 5108 1240 5117 1280
rect 6211 1240 6220 1280
rect 6260 1240 6700 1280
rect 6740 1240 6749 1280
rect 6988 1240 7412 1280
rect 9091 1240 9100 1280
rect 9140 1240 14420 1280
rect 14572 1280 14612 1324
rect 15916 1280 15956 1408
rect 32995 1407 33053 1408
rect 35107 1407 35165 1408
rect 35299 1448 35357 1449
rect 44323 1448 44381 1449
rect 55564 1448 55604 1492
rect 70723 1491 70781 1492
rect 79747 1491 79805 1492
rect 94819 1491 94877 1492
rect 97219 1491 97277 1492
rect 69379 1448 69437 1449
rect 35299 1408 35308 1448
rect 35348 1408 35442 1448
rect 36355 1408 36364 1448
rect 36404 1408 37132 1448
rect 37172 1408 37181 1448
rect 37228 1408 37820 1448
rect 44238 1408 44332 1448
rect 44372 1408 44381 1448
rect 54403 1408 54412 1448
rect 54452 1408 55084 1448
rect 55124 1408 55604 1448
rect 55660 1408 57772 1448
rect 57812 1408 58156 1448
rect 58196 1408 58205 1448
rect 63628 1408 69388 1448
rect 69428 1408 69437 1448
rect 35299 1407 35357 1408
rect 30691 1364 30749 1365
rect 37228 1364 37268 1408
rect 19084 1324 26092 1364
rect 26132 1324 26141 1364
rect 30606 1324 30700 1364
rect 30740 1324 30749 1364
rect 31843 1324 31852 1364
rect 31892 1324 37268 1364
rect 37780 1364 37820 1408
rect 44323 1407 44381 1408
rect 51427 1364 51485 1365
rect 55660 1364 55700 1408
rect 62851 1364 62909 1365
rect 37780 1324 38092 1364
rect 38132 1324 43372 1364
rect 43412 1324 43421 1364
rect 45859 1324 45868 1364
rect 45908 1324 49804 1364
rect 49844 1324 49853 1364
rect 50380 1324 51052 1364
rect 51092 1324 51436 1364
rect 51476 1324 51485 1364
rect 54211 1324 54220 1364
rect 54260 1324 55372 1364
rect 55412 1324 55421 1364
rect 55564 1324 55700 1364
rect 55747 1324 55756 1364
rect 55796 1324 56332 1364
rect 56372 1324 56381 1364
rect 62851 1324 62860 1364
rect 62900 1324 63052 1364
rect 63092 1324 63101 1364
rect 16771 1280 16829 1281
rect 14572 1240 15244 1280
rect 15284 1240 15293 1280
rect 15916 1240 16396 1280
rect 16436 1240 16445 1280
rect 16686 1240 16780 1280
rect 16820 1240 16829 1280
rect 4771 1239 4829 1240
rect 6211 1239 6269 1240
rect 6988 1196 7028 1240
rect 7171 1196 7229 1197
rect 7372 1196 7412 1240
rect 16771 1239 16829 1240
rect 17539 1280 17597 1281
rect 19084 1280 19124 1324
rect 30691 1323 30749 1324
rect 19267 1280 19325 1281
rect 26179 1280 26237 1281
rect 32611 1280 32669 1281
rect 35107 1280 35165 1281
rect 39619 1280 39677 1281
rect 49219 1280 49277 1281
rect 49507 1280 49565 1281
rect 17539 1240 17548 1280
rect 17588 1240 19084 1280
rect 19124 1240 19133 1280
rect 19267 1240 19276 1280
rect 19316 1240 19468 1280
rect 19508 1240 19517 1280
rect 19843 1240 19852 1280
rect 19892 1240 25268 1280
rect 25699 1240 25708 1280
rect 25748 1240 25900 1280
rect 25940 1240 26132 1280
rect 17539 1239 17597 1240
rect 19267 1239 19325 1240
rect 7555 1196 7613 1197
rect 8323 1196 8381 1197
rect 13315 1196 13373 1197
rect 14083 1196 14141 1197
rect 14851 1196 14909 1197
rect 18307 1196 18365 1197
rect 19939 1196 19997 1197
rect 835 1156 844 1196
rect 884 1156 1516 1196
rect 1556 1156 1565 1196
rect 1795 1156 1804 1196
rect 1844 1156 2572 1196
rect 2612 1156 2956 1196
rect 2996 1156 3340 1196
rect 3380 1156 3389 1196
rect 3532 1156 4436 1196
rect 4483 1156 4492 1196
rect 4532 1156 4876 1196
rect 4916 1156 5260 1196
rect 5300 1156 5644 1196
rect 5684 1156 6124 1196
rect 6164 1156 6412 1196
rect 6452 1156 6461 1196
rect 6979 1156 6988 1196
rect 7028 1156 7037 1196
rect 7086 1156 7180 1196
rect 7220 1156 7229 1196
rect 7363 1156 7372 1196
rect 7412 1156 7421 1196
rect 7555 1156 7564 1196
rect 7604 1156 7698 1196
rect 8238 1156 8332 1196
rect 8372 1156 8381 1196
rect 8515 1156 8524 1196
rect 8564 1156 8908 1196
rect 8948 1156 9292 1196
rect 9332 1156 9676 1196
rect 9716 1156 10060 1196
rect 10100 1156 10444 1196
rect 10484 1156 10828 1196
rect 10868 1156 11212 1196
rect 11252 1156 11596 1196
rect 11636 1156 11980 1196
rect 12020 1156 12364 1196
rect 12404 1156 12652 1196
rect 12692 1156 13036 1196
rect 13076 1156 13085 1196
rect 13230 1156 13324 1196
rect 13364 1156 13373 1196
rect 13998 1156 14092 1196
rect 14132 1156 14141 1196
rect 14766 1156 14860 1196
rect 14900 1156 14909 1196
rect 15043 1156 15052 1196
rect 15092 1156 15436 1196
rect 15476 1156 15820 1196
rect 15860 1156 16204 1196
rect 16244 1156 16588 1196
rect 16628 1156 16972 1196
rect 17012 1156 17356 1196
rect 17396 1156 17876 1196
rect 18222 1156 18316 1196
rect 18356 1156 18365 1196
rect 19267 1156 19276 1196
rect 19316 1156 19325 1196
rect 19854 1156 19948 1196
rect 19988 1156 19997 1196
rect 1219 1112 1277 1113
rect 1603 1112 1661 1113
rect 1987 1112 2045 1113
rect 2188 1112 2228 1156
rect 2755 1112 2813 1113
rect 3532 1112 3572 1156
rect 4291 1112 4349 1113
rect 1134 1072 1228 1112
rect 1268 1072 1277 1112
rect 1518 1072 1612 1112
rect 1652 1072 1661 1112
rect 1902 1072 1996 1112
rect 2036 1072 2045 1112
rect 2179 1072 2188 1112
rect 2228 1072 2237 1112
rect 2670 1072 2764 1112
rect 2804 1072 2813 1112
rect 3139 1072 3148 1112
rect 3188 1072 3197 1112
rect 3523 1072 3532 1112
rect 3572 1072 3581 1112
rect 3907 1072 3916 1112
rect 3956 1072 3965 1112
rect 4206 1072 4300 1112
rect 4340 1072 4349 1112
rect 1219 1071 1277 1072
rect 1603 1071 1661 1072
rect 1987 1071 2045 1072
rect 2755 1071 2813 1072
rect 2371 652 2380 692
rect 2420 652 2540 692
rect 2500 104 2540 652
rect 3148 440 3188 1072
rect 3916 860 3956 1072
rect 4291 1071 4349 1072
rect 4396 944 4436 1156
rect 7171 1155 7229 1156
rect 4675 1112 4733 1113
rect 6499 1112 6557 1113
rect 4590 1072 4684 1112
rect 4724 1072 4733 1112
rect 6414 1072 6508 1112
rect 6548 1072 6557 1112
rect 7372 1112 7412 1156
rect 7555 1155 7613 1156
rect 8323 1155 8381 1156
rect 8524 1112 8564 1156
rect 13315 1155 13373 1156
rect 14083 1155 14141 1156
rect 14851 1155 14909 1156
rect 9859 1112 9917 1113
rect 10243 1112 10301 1113
rect 10627 1112 10685 1113
rect 7372 1072 7756 1112
rect 7796 1072 8140 1112
rect 8180 1072 8564 1112
rect 9091 1072 9100 1112
rect 9140 1072 9149 1112
rect 9774 1072 9868 1112
rect 9908 1072 9917 1112
rect 10158 1072 10252 1112
rect 10292 1072 10301 1112
rect 10542 1072 10636 1112
rect 10676 1072 10685 1112
rect 4675 1071 4733 1072
rect 6499 1071 6557 1072
rect 9100 1028 9140 1072
rect 9859 1071 9917 1072
rect 10243 1071 10301 1072
rect 10627 1071 10685 1072
rect 11491 1112 11549 1113
rect 12259 1112 12317 1113
rect 12547 1112 12605 1113
rect 12931 1112 12989 1113
rect 15052 1112 15092 1156
rect 16003 1112 16061 1113
rect 17836 1112 17876 1156
rect 18307 1155 18365 1156
rect 19276 1112 19316 1156
rect 19939 1155 19997 1156
rect 20227 1196 20285 1197
rect 20995 1196 21053 1197
rect 22531 1196 22589 1197
rect 23299 1196 23357 1197
rect 24451 1196 24509 1197
rect 20227 1156 20236 1196
rect 20276 1156 20370 1196
rect 20910 1156 21004 1196
rect 21044 1156 21053 1196
rect 21187 1156 21196 1196
rect 21236 1156 21580 1196
rect 21620 1156 21964 1196
rect 22004 1156 22388 1196
rect 22446 1156 22540 1196
rect 22580 1156 22589 1196
rect 23214 1156 23308 1196
rect 23348 1156 23357 1196
rect 24366 1156 24460 1196
rect 24500 1156 24509 1196
rect 24643 1156 24652 1196
rect 24692 1156 25036 1196
rect 25076 1156 25085 1196
rect 20227 1155 20285 1156
rect 20995 1155 21053 1156
rect 21196 1112 21236 1156
rect 22147 1112 22205 1113
rect 22348 1112 22388 1156
rect 22531 1155 22589 1156
rect 23299 1155 23357 1156
rect 24451 1155 24509 1156
rect 23779 1112 23837 1113
rect 24652 1112 24692 1156
rect 24835 1112 24893 1113
rect 11491 1072 11500 1112
rect 11540 1072 11634 1112
rect 12163 1072 12172 1112
rect 12212 1072 12268 1112
rect 12308 1072 12317 1112
rect 12462 1072 12556 1112
rect 12596 1072 12605 1112
rect 12846 1072 12940 1112
rect 12980 1072 12989 1112
rect 13123 1072 13132 1112
rect 13172 1072 13516 1112
rect 13556 1072 13900 1112
rect 13940 1072 14284 1112
rect 14324 1072 14668 1112
rect 14708 1072 15092 1112
rect 15918 1072 16012 1112
rect 16052 1072 16061 1112
rect 11491 1071 11549 1072
rect 12259 1071 12317 1072
rect 12547 1071 12605 1072
rect 12931 1071 12989 1072
rect 16003 1071 16061 1072
rect 16684 1072 17164 1112
rect 17204 1072 17213 1112
rect 17635 1072 17644 1112
rect 17684 1072 17693 1112
rect 17827 1072 17836 1112
rect 17876 1072 18028 1112
rect 18068 1072 18508 1112
rect 18548 1072 18892 1112
rect 18932 1072 19180 1112
rect 19220 1072 19229 1112
rect 19276 1072 19660 1112
rect 19700 1072 20044 1112
rect 20084 1072 20428 1112
rect 20468 1072 20812 1112
rect 20852 1072 21236 1112
rect 22062 1072 22156 1112
rect 22196 1072 22205 1112
rect 22339 1072 22348 1112
rect 22388 1072 22732 1112
rect 22772 1072 23116 1112
rect 23156 1072 23500 1112
rect 23540 1072 23549 1112
rect 23694 1072 23788 1112
rect 23828 1072 23837 1112
rect 16387 1028 16445 1029
rect 6316 988 9140 1028
rect 9475 988 9484 1028
rect 9524 988 14324 1028
rect 6316 944 6356 988
rect 4396 904 6356 944
rect 6403 944 6461 945
rect 6883 944 6941 945
rect 14284 944 14324 988
rect 14476 988 15628 1028
rect 15668 988 16148 1028
rect 16302 988 16396 1028
rect 16436 988 16445 1028
rect 14476 944 14516 988
rect 16108 944 16148 988
rect 16387 987 16445 988
rect 16579 944 16637 945
rect 6403 904 6412 944
rect 6452 904 6546 944
rect 6798 904 6807 944
rect 6847 904 6892 944
rect 6932 904 6941 944
rect 7267 904 7276 944
rect 7316 904 7564 944
rect 7604 904 7613 944
rect 8035 904 8044 944
rect 8084 904 8332 944
rect 8372 904 8381 944
rect 8803 904 8812 944
rect 8852 904 9100 944
rect 9140 904 9149 944
rect 9571 904 9580 944
rect 9620 904 9868 944
rect 9908 904 9917 944
rect 10339 904 10348 944
rect 10388 904 10636 944
rect 10676 904 10685 944
rect 11107 904 11116 944
rect 11156 904 11404 944
rect 11444 904 11453 944
rect 12259 904 12268 944
rect 12308 904 12556 944
rect 12596 904 12605 944
rect 13027 904 13036 944
rect 13076 904 13324 944
rect 13364 904 13373 944
rect 13795 904 13804 944
rect 13844 904 14092 944
rect 14132 904 14141 944
rect 14284 904 14516 944
rect 14563 904 14572 944
rect 14612 904 14860 944
rect 14900 904 14909 944
rect 15715 904 15724 944
rect 15764 904 16012 944
rect 16052 904 16061 944
rect 16108 904 16588 944
rect 16628 904 16637 944
rect 6403 903 6461 904
rect 6883 903 6941 904
rect 16579 903 16637 904
rect 12067 860 12125 861
rect 14371 860 14429 861
rect 16684 860 16724 1072
rect 17539 944 17597 945
rect 16867 904 16876 944
rect 16916 904 17164 944
rect 17204 904 17213 944
rect 17454 904 17548 944
rect 17588 904 17597 944
rect 17539 903 17597 904
rect 3916 820 9484 860
rect 9524 820 9533 860
rect 11320 820 11692 860
rect 11732 820 11741 860
rect 12067 820 12076 860
rect 12116 820 14380 860
rect 14420 820 14429 860
rect 16675 820 16684 860
rect 16724 820 16733 860
rect 11320 776 11360 820
rect 12067 819 12125 820
rect 14371 819 14429 820
rect 13699 776 13757 777
rect 16771 776 16829 777
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 6211 736 6220 776
rect 6260 736 11360 776
rect 13614 736 13708 776
rect 13748 736 13757 776
rect 14563 736 14572 776
rect 14612 736 16780 776
rect 16820 736 16829 776
rect 17644 776 17684 1072
rect 22147 1071 22205 1072
rect 18691 1028 18749 1029
rect 17923 988 17932 1028
rect 17972 988 18452 1028
rect 18606 988 18700 1028
rect 18740 988 18749 1028
rect 17731 904 17740 944
rect 17780 904 17972 944
rect 18019 904 18028 944
rect 18068 904 18316 944
rect 18356 904 18365 944
rect 17932 860 17972 904
rect 18412 860 18452 988
rect 18691 987 18749 988
rect 19363 1028 19421 1029
rect 20611 1028 20669 1029
rect 22915 1028 22973 1029
rect 19363 988 19372 1028
rect 19412 988 19852 1028
rect 19892 988 19901 1028
rect 20526 988 20620 1028
rect 20660 988 20669 1028
rect 22830 988 22924 1028
rect 22964 988 22973 1028
rect 23500 1028 23540 1072
rect 23779 1071 23837 1072
rect 23884 1072 24268 1112
rect 24308 1072 24692 1112
rect 24750 1072 24844 1112
rect 24884 1072 24893 1112
rect 23884 1028 23924 1072
rect 24835 1071 24893 1072
rect 25228 1028 25268 1240
rect 25507 1112 25565 1113
rect 26092 1112 26132 1240
rect 26179 1240 26188 1280
rect 26228 1240 27436 1280
rect 27476 1240 31028 1280
rect 31651 1240 31660 1280
rect 31700 1240 32140 1280
rect 32180 1240 32189 1280
rect 32526 1240 32620 1280
rect 32660 1240 32669 1280
rect 33859 1240 33868 1280
rect 33908 1240 34444 1280
rect 34484 1240 34493 1280
rect 35107 1240 35116 1280
rect 35156 1240 39572 1280
rect 26179 1239 26237 1240
rect 26659 1196 26717 1197
rect 28195 1196 28253 1197
rect 26574 1156 26668 1196
rect 26708 1156 26717 1196
rect 28110 1156 28204 1196
rect 28244 1156 28253 1196
rect 26659 1155 26717 1156
rect 28195 1155 28253 1156
rect 28780 1156 29164 1196
rect 29204 1156 29548 1196
rect 29588 1156 29932 1196
rect 29972 1156 30316 1196
rect 30356 1156 30740 1196
rect 28780 1112 28820 1156
rect 29731 1112 29789 1113
rect 30115 1112 30173 1113
rect 30700 1112 30740 1156
rect 25422 1072 25516 1112
rect 25556 1072 25565 1112
rect 25987 1072 25996 1112
rect 26036 1072 26045 1112
rect 26092 1072 26476 1112
rect 26516 1072 26860 1112
rect 26900 1072 27244 1112
rect 27284 1072 27628 1112
rect 27668 1072 28012 1112
rect 28052 1072 28300 1112
rect 28340 1072 28780 1112
rect 28820 1072 28829 1112
rect 28963 1072 28972 1112
rect 29012 1072 29021 1112
rect 29646 1072 29740 1112
rect 29780 1072 29789 1112
rect 30030 1072 30124 1112
rect 30164 1072 30173 1112
rect 30691 1072 30700 1112
rect 30740 1072 30892 1112
rect 30932 1072 30941 1112
rect 25507 1071 25565 1072
rect 25891 1028 25949 1029
rect 23500 988 23884 1028
rect 23924 988 23933 1028
rect 25228 988 25900 1028
rect 25940 988 25949 1028
rect 19363 987 19421 988
rect 20611 987 20669 988
rect 22915 987 22973 988
rect 25891 987 25949 988
rect 25996 944 26036 1072
rect 26092 1028 26132 1072
rect 27619 1028 27677 1029
rect 28972 1028 29012 1072
rect 29731 1071 29789 1072
rect 30115 1071 30173 1072
rect 26083 988 26092 1028
rect 26132 988 26141 1028
rect 27619 988 27628 1028
rect 27668 988 29012 1028
rect 30988 1028 31028 1240
rect 32611 1239 32669 1240
rect 35107 1239 35165 1240
rect 31843 1196 31901 1197
rect 32227 1196 32285 1197
rect 31758 1156 31852 1196
rect 31892 1156 31901 1196
rect 32142 1156 32236 1196
rect 32276 1156 32285 1196
rect 31843 1155 31901 1156
rect 32227 1155 32285 1156
rect 34147 1196 34205 1197
rect 38467 1196 38525 1197
rect 38851 1196 38909 1197
rect 39235 1196 39293 1197
rect 34147 1156 34156 1196
rect 34196 1156 34290 1196
rect 34348 1156 34732 1196
rect 34772 1156 35116 1196
rect 35156 1156 35500 1196
rect 35540 1156 35884 1196
rect 35924 1156 36268 1196
rect 36308 1156 36692 1196
rect 38382 1156 38476 1196
rect 38516 1156 38525 1196
rect 38766 1156 38860 1196
rect 38900 1156 38909 1196
rect 39150 1156 39244 1196
rect 39284 1156 39293 1196
rect 39532 1196 39572 1240
rect 39619 1240 39628 1280
rect 39668 1240 42028 1280
rect 42068 1240 42077 1280
rect 42307 1240 42316 1280
rect 42356 1240 48556 1280
rect 48596 1240 49228 1280
rect 49268 1240 49277 1280
rect 49422 1240 49516 1280
rect 49556 1240 49565 1280
rect 39619 1239 39677 1240
rect 49219 1239 49277 1240
rect 49507 1239 49565 1240
rect 40003 1196 40061 1197
rect 40387 1196 40445 1197
rect 42691 1196 42749 1197
rect 44419 1196 44477 1197
rect 46243 1196 46301 1197
rect 47779 1196 47837 1197
rect 39532 1156 40012 1196
rect 40052 1156 40061 1196
rect 40302 1156 40396 1196
rect 40436 1156 40445 1196
rect 34147 1155 34205 1156
rect 31075 1112 31133 1113
rect 31459 1112 31517 1113
rect 34348 1112 34388 1156
rect 31075 1072 31084 1112
rect 31124 1072 31218 1112
rect 31374 1072 31468 1112
rect 31508 1072 31517 1112
rect 31651 1072 31660 1112
rect 31700 1072 32044 1112
rect 32084 1072 32428 1112
rect 32468 1072 32812 1112
rect 32852 1072 33196 1112
rect 33236 1072 33580 1112
rect 33620 1072 33964 1112
rect 34004 1072 34252 1112
rect 34292 1072 34388 1112
rect 34531 1112 34589 1113
rect 35011 1112 35069 1113
rect 34531 1072 34540 1112
rect 34580 1072 35020 1112
rect 35060 1072 35069 1112
rect 31075 1071 31133 1072
rect 31459 1071 31517 1072
rect 34531 1071 34589 1072
rect 35011 1071 35069 1072
rect 35395 1112 35453 1113
rect 36652 1112 36692 1156
rect 38467 1155 38525 1156
rect 38851 1155 38909 1156
rect 39235 1155 39293 1156
rect 40003 1155 40061 1156
rect 40387 1155 40445 1156
rect 40588 1156 40972 1196
rect 41012 1156 42124 1196
rect 42164 1156 42508 1196
rect 42548 1156 42557 1196
rect 42606 1156 42700 1196
rect 42740 1156 42749 1196
rect 43363 1156 43372 1196
rect 43412 1156 44343 1196
rect 44383 1156 44428 1196
rect 44468 1156 44477 1196
rect 45091 1156 45100 1196
rect 45140 1156 45964 1196
rect 46004 1156 46013 1196
rect 46158 1156 46252 1196
rect 46292 1156 46301 1196
rect 46627 1156 46636 1196
rect 46676 1156 47788 1196
rect 47828 1156 47837 1196
rect 37027 1112 37085 1113
rect 37315 1112 37373 1113
rect 40588 1112 40628 1156
rect 40771 1112 40829 1113
rect 41356 1112 41396 1156
rect 41539 1112 41597 1113
rect 41740 1112 41780 1156
rect 42403 1112 42461 1113
rect 35395 1072 35404 1112
rect 35444 1072 35538 1112
rect 35971 1072 35980 1112
rect 36020 1072 36364 1112
rect 36404 1072 36413 1112
rect 36643 1072 36652 1112
rect 36692 1072 36844 1112
rect 36884 1072 36893 1112
rect 37027 1072 37036 1112
rect 37076 1072 37170 1112
rect 37315 1072 37324 1112
rect 37364 1072 37458 1112
rect 37507 1072 37516 1112
rect 37556 1072 37900 1112
rect 37940 1072 38284 1112
rect 38324 1072 38668 1112
rect 38708 1072 39052 1112
rect 39092 1072 39436 1112
rect 39476 1072 39820 1112
rect 39860 1072 40204 1112
rect 40244 1072 40588 1112
rect 40628 1072 40637 1112
rect 40686 1072 40780 1112
rect 40820 1072 40829 1112
rect 41155 1072 41164 1112
rect 41204 1072 41213 1112
rect 41347 1072 41356 1112
rect 41396 1072 41405 1112
rect 41454 1072 41548 1112
rect 41588 1072 41597 1112
rect 41731 1072 41740 1112
rect 41780 1072 41789 1112
rect 42019 1072 42028 1112
rect 42068 1072 42164 1112
rect 42307 1072 42316 1112
rect 42356 1072 42412 1112
rect 42452 1072 42461 1112
rect 42508 1112 42548 1156
rect 42691 1155 42749 1156
rect 44419 1155 44477 1156
rect 46243 1155 46301 1156
rect 47779 1155 47837 1156
rect 48067 1196 48125 1197
rect 49699 1196 49757 1197
rect 50380 1196 50420 1324
rect 51427 1323 51485 1324
rect 55564 1280 55604 1324
rect 62851 1323 62909 1324
rect 63628 1280 63668 1408
rect 69379 1407 69437 1408
rect 73027 1448 73085 1449
rect 81475 1448 81533 1449
rect 88387 1448 88445 1449
rect 94915 1448 94973 1449
rect 73027 1408 73036 1448
rect 73076 1408 73748 1448
rect 73987 1408 73996 1448
rect 74036 1408 74956 1448
rect 74996 1408 75005 1448
rect 75532 1408 81484 1448
rect 81524 1408 81533 1448
rect 83875 1408 83884 1448
rect 83924 1408 88220 1448
rect 88302 1408 88396 1448
rect 88436 1408 94348 1448
rect 94388 1408 94397 1448
rect 94830 1408 94924 1448
rect 94964 1408 94973 1448
rect 73027 1407 73085 1408
rect 64195 1364 64253 1365
rect 64675 1364 64733 1365
rect 65251 1364 65309 1365
rect 66883 1364 66941 1365
rect 71491 1364 71549 1365
rect 72259 1364 72317 1365
rect 64110 1324 64204 1364
rect 64244 1324 64253 1364
rect 64590 1324 64684 1364
rect 64724 1324 64733 1364
rect 64195 1323 64253 1324
rect 64675 1323 64733 1324
rect 64780 1324 65260 1364
rect 65300 1324 65309 1364
rect 66798 1324 66892 1364
rect 66932 1324 66941 1364
rect 64780 1280 64820 1324
rect 65251 1323 65309 1324
rect 66883 1323 66941 1324
rect 70156 1324 70772 1364
rect 70156 1280 70196 1324
rect 70732 1280 70772 1324
rect 71491 1324 71500 1364
rect 71540 1324 71788 1364
rect 71828 1324 71837 1364
rect 72174 1324 72268 1364
rect 72308 1324 72317 1364
rect 71491 1323 71549 1324
rect 72259 1323 72317 1324
rect 72835 1280 72893 1281
rect 50563 1240 50572 1280
rect 50612 1240 50956 1280
rect 50996 1240 51005 1280
rect 52195 1240 52204 1280
rect 52244 1240 52588 1280
rect 52628 1240 55604 1280
rect 55651 1240 55660 1280
rect 55700 1240 56140 1280
rect 56180 1240 56189 1280
rect 56428 1240 56716 1280
rect 56756 1240 56765 1280
rect 59299 1240 59308 1280
rect 59348 1240 59884 1280
rect 59924 1240 59933 1280
rect 60643 1240 60652 1280
rect 60692 1240 60940 1280
rect 60980 1240 60989 1280
rect 63052 1240 63668 1280
rect 63715 1240 63724 1280
rect 63764 1240 64820 1280
rect 64867 1240 64876 1280
rect 64916 1240 66508 1280
rect 66548 1240 69236 1280
rect 50956 1196 50996 1240
rect 56428 1196 56468 1240
rect 62755 1196 62813 1197
rect 63052 1196 63092 1240
rect 63523 1196 63581 1197
rect 67267 1196 67325 1197
rect 68035 1196 68093 1197
rect 48067 1156 48076 1196
rect 48116 1156 48167 1196
rect 48207 1156 48216 1196
rect 48259 1156 48268 1196
rect 48308 1156 48317 1196
rect 48739 1156 48748 1196
rect 48788 1156 49132 1196
rect 49172 1156 49324 1196
rect 49364 1156 49373 1196
rect 49614 1156 49708 1196
rect 49748 1156 49757 1196
rect 50371 1156 50380 1196
rect 50420 1156 50429 1196
rect 50956 1156 56428 1196
rect 56468 1156 56477 1196
rect 62755 1156 62764 1196
rect 62804 1156 63052 1196
rect 63092 1156 63101 1196
rect 63438 1156 63532 1196
rect 63572 1156 63581 1196
rect 64003 1156 64012 1196
rect 64052 1156 64396 1196
rect 64436 1156 64780 1196
rect 64820 1156 65164 1196
rect 65204 1156 65548 1196
rect 65588 1156 65932 1196
rect 65972 1156 66316 1196
rect 66356 1156 66700 1196
rect 66740 1156 67084 1196
rect 67124 1156 67133 1196
rect 67267 1156 67276 1196
rect 67316 1156 67410 1196
rect 67950 1156 68044 1196
rect 68084 1156 68093 1196
rect 69196 1196 69236 1240
rect 69580 1240 70196 1280
rect 70243 1240 70252 1280
rect 70292 1240 70636 1280
rect 70676 1240 70685 1280
rect 70732 1240 72844 1280
rect 72884 1240 72893 1280
rect 69580 1196 69620 1240
rect 72835 1239 72893 1240
rect 69763 1196 69821 1197
rect 70147 1196 70205 1197
rect 70435 1196 70493 1197
rect 72067 1196 72125 1197
rect 72451 1196 72509 1197
rect 72931 1196 72989 1197
rect 73603 1196 73661 1197
rect 69196 1156 69620 1196
rect 69678 1156 69772 1196
rect 69812 1156 69821 1196
rect 70062 1156 70156 1196
rect 70196 1156 70205 1196
rect 70426 1156 70444 1196
rect 70484 1156 70521 1196
rect 70561 1156 70570 1196
rect 71982 1156 72076 1196
rect 72116 1156 72125 1196
rect 72366 1156 72460 1196
rect 72500 1156 72940 1196
rect 72980 1156 72989 1196
rect 73518 1156 73612 1196
rect 73652 1156 73661 1196
rect 73708 1196 73748 1408
rect 74851 1324 74860 1364
rect 74900 1324 75052 1364
rect 75092 1324 75101 1364
rect 75532 1281 75572 1408
rect 81475 1407 81533 1408
rect 80515 1364 80573 1365
rect 82819 1364 82877 1365
rect 85315 1364 85373 1365
rect 79852 1324 80044 1364
rect 80084 1324 80093 1364
rect 80430 1324 80524 1364
rect 80564 1324 80573 1364
rect 82734 1324 82828 1364
rect 82868 1324 82877 1364
rect 85230 1324 85324 1364
rect 85364 1324 85373 1364
rect 75523 1280 75581 1281
rect 79171 1280 79229 1281
rect 75438 1240 75532 1280
rect 75572 1240 75581 1280
rect 79086 1240 79180 1280
rect 79220 1240 79229 1280
rect 79363 1240 79372 1280
rect 79412 1240 79564 1280
rect 79604 1240 79613 1280
rect 75523 1239 75581 1240
rect 79171 1239 79229 1240
rect 79852 1196 79892 1324
rect 80515 1323 80573 1324
rect 82819 1323 82877 1324
rect 85315 1323 85373 1324
rect 81091 1280 81149 1281
rect 85699 1280 85757 1281
rect 87619 1280 87677 1281
rect 80419 1240 80428 1280
rect 80468 1240 80908 1280
rect 80948 1240 80957 1280
rect 81091 1240 81100 1280
rect 81140 1240 81234 1280
rect 85614 1240 85708 1280
rect 85748 1240 85757 1280
rect 87534 1240 87628 1280
rect 87668 1240 87677 1280
rect 88180 1280 88220 1408
rect 88387 1407 88445 1408
rect 94915 1407 94973 1408
rect 88771 1364 88829 1365
rect 88686 1324 88780 1364
rect 88820 1324 88829 1364
rect 89347 1324 89356 1364
rect 89396 1324 89740 1364
rect 89780 1324 90124 1364
rect 90164 1324 90508 1364
rect 90548 1324 90892 1364
rect 90932 1324 91276 1364
rect 91316 1324 91660 1364
rect 91700 1324 92044 1364
rect 92084 1324 92428 1364
rect 92468 1324 92477 1364
rect 97987 1324 97996 1364
rect 98036 1324 98045 1364
rect 88771 1323 88829 1324
rect 89923 1280 89981 1281
rect 90307 1280 90365 1281
rect 88180 1240 89932 1280
rect 89972 1240 89981 1280
rect 90222 1240 90316 1280
rect 90356 1240 90365 1280
rect 73708 1156 73996 1196
rect 74036 1156 79892 1196
rect 80908 1196 80948 1240
rect 81091 1239 81149 1240
rect 85699 1239 85757 1240
rect 87619 1239 87677 1240
rect 89923 1239 89981 1240
rect 90307 1239 90365 1240
rect 92611 1280 92669 1281
rect 93187 1280 93245 1281
rect 94531 1280 94589 1281
rect 97996 1280 98036 1324
rect 92611 1240 92620 1280
rect 92660 1240 92754 1280
rect 93102 1240 93196 1280
rect 93236 1240 93245 1280
rect 94243 1240 94252 1280
rect 94292 1240 94540 1280
rect 94580 1240 94589 1280
rect 95587 1240 95596 1280
rect 95636 1240 96172 1280
rect 96212 1240 96221 1280
rect 97996 1240 98860 1280
rect 98900 1240 98909 1280
rect 92611 1239 92669 1240
rect 93187 1239 93245 1240
rect 94531 1239 94589 1240
rect 86947 1196 87005 1197
rect 88003 1196 88061 1197
rect 89155 1196 89213 1197
rect 89539 1196 89597 1197
rect 80908 1156 81292 1196
rect 81332 1156 81676 1196
rect 81716 1156 82060 1196
rect 82100 1156 82444 1196
rect 82484 1156 82828 1196
rect 82868 1156 83212 1196
rect 83252 1156 83596 1196
rect 83636 1156 83980 1196
rect 84020 1156 84364 1196
rect 84404 1156 84748 1196
rect 84788 1156 85132 1196
rect 85172 1156 85516 1196
rect 85556 1156 85900 1196
rect 85940 1156 86284 1196
rect 86324 1156 86668 1196
rect 86708 1156 86717 1196
rect 86947 1156 86956 1196
rect 86996 1156 87047 1196
rect 87087 1156 87096 1196
rect 88003 1156 88012 1196
rect 88052 1156 88146 1196
rect 89070 1156 89164 1196
rect 89204 1156 89213 1196
rect 89454 1156 89548 1196
rect 89588 1156 95540 1196
rect 48067 1155 48125 1156
rect 43267 1112 43325 1113
rect 43555 1112 43613 1113
rect 47011 1112 47069 1113
rect 42508 1072 42892 1112
rect 42932 1072 43084 1112
rect 43124 1072 43133 1112
rect 43182 1072 43276 1112
rect 43316 1072 43325 1112
rect 43470 1072 43564 1112
rect 43604 1072 43613 1112
rect 43747 1072 43756 1112
rect 43796 1072 44140 1112
rect 44180 1072 44428 1112
rect 44468 1072 44908 1112
rect 44948 1072 45292 1112
rect 45332 1072 45676 1112
rect 45716 1072 46060 1112
rect 46100 1072 46444 1112
rect 46484 1072 46828 1112
rect 46868 1072 46877 1112
rect 46926 1072 47020 1112
rect 47060 1072 47069 1112
rect 35395 1071 35453 1072
rect 37027 1071 37085 1072
rect 37315 1071 37373 1072
rect 40771 1071 40829 1072
rect 34051 1028 34109 1029
rect 30988 988 33388 1028
rect 33428 988 34060 1028
rect 34100 988 34109 1028
rect 27619 987 27677 988
rect 34051 987 34109 988
rect 34243 1028 34301 1029
rect 39619 1028 39677 1029
rect 34243 988 34252 1028
rect 34292 988 39628 1028
rect 39668 988 39677 1028
rect 34243 987 34301 988
rect 39619 987 39677 988
rect 30499 944 30557 945
rect 31747 944 31805 945
rect 18787 904 18796 944
rect 18836 904 19084 944
rect 19124 904 19133 944
rect 19555 904 19564 944
rect 19604 904 19613 944
rect 19939 904 19948 944
rect 19988 904 20236 944
rect 20276 904 20285 944
rect 20707 904 20716 944
rect 20756 904 21004 944
rect 21044 904 21053 944
rect 22243 904 22252 944
rect 22292 904 22540 944
rect 22580 904 22589 944
rect 23011 904 23020 944
rect 23060 904 23308 944
rect 23348 904 23357 944
rect 23779 904 23788 944
rect 23828 904 24071 944
rect 24111 904 24120 944
rect 24163 904 24172 944
rect 24212 904 24460 944
rect 24500 904 24509 944
rect 24931 904 24940 944
rect 24980 904 25228 944
rect 25268 904 25277 944
rect 25699 904 25708 944
rect 25748 904 26036 944
rect 26371 904 26380 944
rect 26420 904 26668 944
rect 26708 904 26717 944
rect 27139 904 27148 944
rect 27188 904 27436 944
rect 27476 904 27485 944
rect 27907 904 27916 944
rect 27956 904 28204 944
rect 28244 904 28253 944
rect 28675 904 28684 944
rect 28724 904 28972 944
rect 29012 904 29021 944
rect 29827 904 29836 944
rect 29876 904 30124 944
rect 30164 904 30173 944
rect 30414 904 30508 944
rect 30548 904 30557 944
rect 30979 904 30988 944
rect 31028 904 31372 944
rect 31412 904 31421 944
rect 31747 904 31756 944
rect 31796 904 32236 944
rect 32276 904 32285 944
rect 32707 904 32716 944
rect 32756 904 33292 944
rect 33332 904 33341 944
rect 34627 904 34636 944
rect 34676 904 35212 944
rect 35252 904 35261 944
rect 35395 904 35404 944
rect 35444 904 35980 944
rect 36020 904 36029 944
rect 36163 904 36172 944
rect 36212 904 36884 944
rect 37411 904 37420 944
rect 37460 904 37900 944
rect 37940 904 37949 944
rect 38179 904 38188 944
rect 38228 904 38668 944
rect 38708 904 38717 944
rect 38947 904 38956 944
rect 38996 904 39436 944
rect 39476 904 39485 944
rect 39715 904 39724 944
rect 39764 904 40204 944
rect 40244 904 40253 944
rect 40483 904 40492 944
rect 40532 904 40972 944
rect 41012 904 41021 944
rect 19564 860 19604 904
rect 30499 903 30557 904
rect 31747 903 31805 904
rect 20035 860 20093 861
rect 26179 860 26237 861
rect 35107 860 35165 861
rect 36067 860 36125 861
rect 36451 860 36509 861
rect 36844 860 36884 904
rect 41164 860 41204 1072
rect 41539 1071 41597 1072
rect 42019 1028 42077 1029
rect 41934 988 41943 1028
rect 41983 988 42028 1028
rect 42068 988 42077 1028
rect 42124 1028 42164 1072
rect 42403 1071 42461 1072
rect 43267 1071 43325 1072
rect 43555 1071 43613 1072
rect 46627 1028 46685 1029
rect 46828 1028 46868 1072
rect 47011 1071 47069 1072
rect 47683 1112 47741 1113
rect 48268 1112 48308 1156
rect 49699 1155 49757 1156
rect 62755 1155 62813 1156
rect 63523 1155 63581 1156
rect 48931 1112 48989 1113
rect 47683 1072 47692 1112
rect 47732 1072 47788 1112
rect 47828 1072 48308 1112
rect 48846 1072 48940 1112
rect 48980 1072 48989 1112
rect 47683 1071 47741 1072
rect 48931 1071 48989 1072
rect 49123 1112 49181 1113
rect 51427 1112 51485 1113
rect 55939 1112 55997 1113
rect 62659 1112 62717 1113
rect 49123 1072 49132 1112
rect 49172 1072 51148 1112
rect 51188 1072 51197 1112
rect 51342 1072 51436 1112
rect 51476 1072 52204 1112
rect 52244 1072 52684 1112
rect 52724 1072 53548 1112
rect 53588 1072 54124 1112
rect 54164 1072 54508 1112
rect 54548 1072 55084 1112
rect 55124 1072 55564 1112
rect 55604 1072 55613 1112
rect 55854 1072 55948 1112
rect 55988 1072 55997 1112
rect 56611 1072 56620 1112
rect 56660 1072 57100 1112
rect 57140 1072 57772 1112
rect 57812 1072 58348 1112
rect 58388 1072 59116 1112
rect 59156 1072 59596 1112
rect 59636 1072 60172 1112
rect 60212 1072 60652 1112
rect 60692 1072 61132 1112
rect 61172 1072 61181 1112
rect 62574 1072 62668 1112
rect 62708 1072 62717 1112
rect 49123 1071 49181 1072
rect 51427 1071 51485 1072
rect 55939 1071 55997 1072
rect 62659 1071 62717 1072
rect 62947 1112 63005 1113
rect 64012 1112 64052 1156
rect 62947 1072 62956 1112
rect 62996 1072 63244 1112
rect 63284 1072 63628 1112
rect 63668 1072 64052 1112
rect 64291 1112 64349 1113
rect 64579 1112 64637 1113
rect 65443 1112 65501 1113
rect 65731 1112 65789 1113
rect 66787 1112 66845 1113
rect 64291 1072 64300 1112
rect 64340 1072 64434 1112
rect 64494 1072 64588 1112
rect 64628 1072 64637 1112
rect 65358 1072 65452 1112
rect 65492 1072 65501 1112
rect 65646 1072 65740 1112
rect 65780 1072 65789 1112
rect 66115 1072 66124 1112
rect 66164 1072 66796 1112
rect 66836 1072 66845 1112
rect 67084 1112 67124 1156
rect 67267 1155 67325 1156
rect 68035 1155 68093 1156
rect 69763 1155 69821 1156
rect 70147 1155 70205 1156
rect 70435 1155 70493 1156
rect 72067 1155 72125 1156
rect 72451 1155 72509 1156
rect 72931 1155 72989 1156
rect 73603 1155 73661 1156
rect 86947 1155 87005 1156
rect 88003 1155 88061 1156
rect 89155 1155 89213 1156
rect 89539 1155 89597 1156
rect 68611 1112 68669 1113
rect 68803 1112 68861 1113
rect 74755 1112 74813 1113
rect 75907 1112 75965 1113
rect 76291 1112 76349 1113
rect 81859 1112 81917 1113
rect 82243 1112 82301 1113
rect 82627 1112 82685 1113
rect 83011 1112 83069 1113
rect 84163 1112 84221 1113
rect 84547 1112 84605 1113
rect 85603 1112 85661 1113
rect 86467 1112 86525 1113
rect 86851 1112 86909 1113
rect 91075 1112 91133 1113
rect 91459 1112 91517 1113
rect 91843 1112 91901 1113
rect 92995 1112 93053 1113
rect 93571 1112 93629 1113
rect 93955 1112 94013 1113
rect 94723 1112 94781 1113
rect 95500 1112 95540 1156
rect 95788 1156 96076 1196
rect 96116 1156 96460 1196
rect 96500 1156 96844 1196
rect 96884 1156 97228 1196
rect 97268 1156 97612 1196
rect 97652 1156 97996 1196
rect 98036 1156 98380 1196
rect 98420 1156 98764 1196
rect 98804 1156 98956 1196
rect 98996 1156 99005 1196
rect 67084 1072 67468 1112
rect 67508 1072 67852 1112
rect 67892 1072 68236 1112
rect 68276 1072 68428 1112
rect 68468 1072 68477 1112
rect 68611 1072 68620 1112
rect 68660 1072 68754 1112
rect 68803 1072 68812 1112
rect 68852 1072 68946 1112
rect 68995 1072 69004 1112
rect 69044 1072 69196 1112
rect 69236 1072 69676 1112
rect 69716 1072 69964 1112
rect 70004 1072 70348 1112
rect 70388 1072 70636 1112
rect 70676 1072 71116 1112
rect 71156 1072 71500 1112
rect 71540 1072 71884 1112
rect 71924 1072 72268 1112
rect 72308 1072 72652 1112
rect 72692 1072 73036 1112
rect 73076 1072 73420 1112
rect 73460 1072 73804 1112
rect 73844 1072 74188 1112
rect 74228 1072 74572 1112
rect 74612 1072 74621 1112
rect 74670 1072 74764 1112
rect 74804 1072 74813 1112
rect 74947 1072 74956 1112
rect 74996 1072 75340 1112
rect 75380 1072 75724 1112
rect 75764 1072 75773 1112
rect 75907 1072 75916 1112
rect 75956 1072 76050 1112
rect 76099 1072 76108 1112
rect 76148 1072 76157 1112
rect 76206 1072 76300 1112
rect 76340 1072 76349 1112
rect 62947 1071 63005 1072
rect 64291 1071 64349 1072
rect 64579 1071 64637 1072
rect 65443 1071 65501 1072
rect 65731 1071 65789 1072
rect 66787 1071 66845 1072
rect 68611 1071 68669 1072
rect 68803 1071 68861 1072
rect 74755 1071 74813 1072
rect 71299 1028 71357 1029
rect 42124 988 45868 1028
rect 45908 988 45917 1028
rect 46627 988 46636 1028
rect 46676 988 46770 1028
rect 46828 988 47212 1028
rect 47252 988 47596 1028
rect 47636 988 47980 1028
rect 48020 988 48364 1028
rect 48404 988 48748 1028
rect 48788 988 48797 1028
rect 49795 988 49804 1028
rect 49844 988 64972 1028
rect 65012 988 71308 1028
rect 71348 988 71357 1028
rect 75724 1028 75764 1072
rect 75907 1071 75965 1072
rect 76108 1028 76148 1072
rect 76291 1071 76349 1072
rect 77260 1072 77644 1112
rect 77684 1072 78028 1112
rect 78068 1072 78412 1112
rect 78452 1072 78796 1112
rect 78836 1072 79564 1112
rect 79604 1072 79948 1112
rect 79988 1072 80332 1112
rect 80372 1072 80381 1112
rect 81774 1072 81868 1112
rect 81908 1072 81917 1112
rect 82158 1072 82252 1112
rect 82292 1072 82301 1112
rect 82542 1072 82636 1112
rect 82676 1072 82685 1112
rect 82926 1072 83020 1112
rect 83060 1072 83069 1112
rect 83299 1072 83308 1112
rect 83348 1072 83357 1112
rect 84078 1072 84172 1112
rect 84212 1072 84221 1112
rect 84462 1072 84556 1112
rect 84596 1072 84605 1112
rect 84931 1072 84940 1112
rect 84980 1072 85612 1112
rect 85652 1072 85661 1112
rect 86382 1072 86476 1112
rect 86516 1072 86525 1112
rect 86766 1072 86860 1112
rect 86900 1072 86909 1112
rect 87235 1072 87244 1112
rect 87284 1072 87436 1112
rect 87476 1072 87820 1112
rect 87860 1072 88204 1112
rect 88244 1072 88588 1112
rect 88628 1072 88972 1112
rect 89012 1072 89356 1112
rect 89396 1072 89405 1112
rect 90990 1072 91084 1112
rect 91124 1072 91133 1112
rect 91374 1072 91468 1112
rect 91508 1072 91517 1112
rect 91758 1072 91852 1112
rect 91892 1072 91901 1112
rect 92419 1072 92428 1112
rect 92468 1072 92812 1112
rect 92852 1072 92861 1112
rect 92995 1072 93004 1112
rect 93044 1072 93138 1112
rect 93283 1072 93292 1112
rect 93332 1072 93341 1112
rect 93386 1072 93395 1112
rect 93435 1072 93444 1112
rect 93486 1072 93580 1112
rect 93620 1072 93629 1112
rect 93870 1072 93964 1112
rect 94004 1072 94013 1112
rect 94147 1072 94156 1112
rect 94196 1072 94205 1112
rect 94638 1072 94732 1112
rect 94772 1072 94781 1112
rect 77260 1028 77300 1072
rect 81859 1071 81917 1072
rect 82243 1071 82301 1072
rect 82627 1071 82685 1072
rect 83011 1071 83069 1072
rect 78595 1028 78653 1029
rect 83308 1028 83348 1072
rect 84163 1071 84221 1072
rect 84547 1071 84605 1072
rect 85603 1071 85661 1072
rect 86467 1071 86525 1072
rect 86851 1071 86909 1072
rect 91075 1071 91133 1072
rect 91459 1071 91517 1072
rect 91843 1071 91901 1072
rect 92995 1071 93053 1072
rect 89539 1028 89597 1029
rect 75724 988 76492 1028
rect 76532 988 76876 1028
rect 76916 988 77260 1028
rect 77300 988 77309 1028
rect 77443 988 77452 1028
rect 77492 988 78356 1028
rect 42019 987 42077 988
rect 46627 987 46685 988
rect 71299 987 71357 988
rect 45475 944 45533 945
rect 62947 944 63005 945
rect 64003 944 64061 945
rect 65347 944 65405 945
rect 66883 944 66941 945
rect 70915 944 70973 945
rect 72259 944 72317 945
rect 78211 944 78269 945
rect 41251 904 41260 944
rect 41300 904 41740 944
rect 41780 904 41789 944
rect 42019 904 42028 944
rect 42068 904 42508 944
rect 42548 904 42557 944
rect 42787 904 42796 944
rect 42836 904 43276 944
rect 43316 904 43325 944
rect 45390 904 45484 944
rect 45524 904 45533 944
rect 45955 904 45964 944
rect 46004 904 46252 944
rect 46292 904 46301 944
rect 46723 904 46732 944
rect 46772 904 47020 944
rect 47060 904 47069 944
rect 47491 904 47500 944
rect 47540 904 47788 944
rect 47828 904 47837 944
rect 48259 904 48268 944
rect 48308 904 48556 944
rect 48596 904 48605 944
rect 50467 904 50476 944
rect 50516 904 50956 944
rect 50996 904 51005 944
rect 52099 904 52108 944
rect 52148 904 52588 944
rect 52628 904 52637 944
rect 53443 904 53452 944
rect 53492 904 53932 944
rect 53972 904 53981 944
rect 59299 904 59308 944
rect 59348 904 59500 944
rect 59540 904 59549 944
rect 60547 904 60556 944
rect 60596 904 61036 944
rect 61076 904 61085 944
rect 62467 904 62476 944
rect 62516 904 62764 944
rect 62804 904 62813 944
rect 62856 904 62865 944
rect 62905 904 62956 944
rect 62996 904 63005 944
rect 63235 904 63244 944
rect 63284 904 63532 944
rect 63572 904 63581 944
rect 63811 904 63820 944
rect 63860 904 64012 944
rect 64052 904 64061 944
rect 64176 904 64204 944
rect 64244 904 64300 944
rect 64340 904 64349 944
rect 64588 904 64876 944
rect 64916 904 64925 944
rect 65059 904 65068 944
rect 65108 904 65117 944
rect 65262 904 65356 944
rect 65396 904 65405 944
rect 65539 904 65548 944
rect 65588 904 65836 944
rect 65876 904 65885 944
rect 66691 904 66700 944
rect 66740 904 66892 944
rect 66932 904 66941 944
rect 67075 904 67084 944
rect 67124 904 67372 944
rect 67412 904 67421 944
rect 68227 904 68236 944
rect 68276 904 68524 944
rect 68564 904 68573 944
rect 69379 904 69388 944
rect 69428 904 69676 944
rect 69716 904 69725 944
rect 70147 904 70156 944
rect 70196 904 70444 944
rect 70484 904 70493 944
rect 70915 904 70924 944
rect 70964 904 71212 944
rect 71252 904 71261 944
rect 71683 904 71692 944
rect 71732 904 71884 944
rect 71924 904 71933 944
rect 72067 904 72076 944
rect 72116 904 72268 944
rect 72308 904 72317 944
rect 72835 904 72844 944
rect 72884 904 73132 944
rect 73172 904 73181 944
rect 73603 904 73612 944
rect 73652 904 73900 944
rect 73940 904 73949 944
rect 74371 904 74380 944
rect 74420 904 74429 944
rect 74755 904 74764 944
rect 74804 904 75052 944
rect 75092 904 75101 944
rect 75523 904 75532 944
rect 75572 904 75820 944
rect 75860 904 75869 944
rect 76291 904 76300 944
rect 76340 904 76588 944
rect 76628 904 76637 944
rect 77059 904 77068 944
rect 77108 904 77356 944
rect 77396 904 77405 944
rect 78126 904 78220 944
rect 78260 904 78269 944
rect 78316 944 78356 988
rect 78595 988 78604 1028
rect 78644 988 78738 1028
rect 78796 988 89548 1028
rect 89588 988 89597 1028
rect 78595 987 78653 988
rect 78796 944 78836 988
rect 89539 987 89597 988
rect 90691 1028 90749 1029
rect 92035 1028 92093 1029
rect 90691 988 90700 1028
rect 90740 988 92044 1028
rect 92084 988 92093 1028
rect 90691 987 90749 988
rect 92035 987 92093 988
rect 82243 944 82301 945
rect 88387 944 88445 945
rect 78316 904 78836 944
rect 78979 904 78988 944
rect 79028 904 79276 944
rect 79316 904 79325 944
rect 79747 904 79756 944
rect 79796 904 80044 944
rect 80084 904 80093 944
rect 80227 904 80236 944
rect 80276 904 80524 944
rect 80564 904 80573 944
rect 82243 904 82252 944
rect 82292 904 88396 944
rect 88436 904 88445 944
rect 45475 903 45533 904
rect 62947 903 63005 904
rect 64003 903 64061 904
rect 54979 860 55037 861
rect 64588 860 64628 904
rect 65068 860 65108 904
rect 65347 903 65405 904
rect 66883 903 66941 904
rect 70915 903 70973 904
rect 72259 903 72317 904
rect 74380 861 74420 904
rect 78211 903 78269 904
rect 82243 903 82301 904
rect 88387 903 88445 904
rect 17923 820 17932 860
rect 17972 820 17981 860
rect 18412 820 18700 860
rect 18740 820 18749 860
rect 19564 820 20044 860
rect 20084 820 20093 860
rect 20035 819 20093 820
rect 20140 820 21388 860
rect 21428 820 26188 860
rect 26228 820 26237 860
rect 27811 820 27820 860
rect 27860 820 33772 860
rect 33812 820 35116 860
rect 35156 820 35165 860
rect 35683 820 35692 860
rect 35732 820 36076 860
rect 36116 820 36125 860
rect 36366 820 36460 860
rect 36500 820 36509 860
rect 36835 820 36844 860
rect 36884 820 36893 860
rect 37780 820 47404 860
rect 47444 820 54988 860
rect 55028 820 64628 860
rect 64684 820 65108 860
rect 65251 860 65309 861
rect 70147 860 70205 861
rect 71491 860 71549 861
rect 74371 860 74429 861
rect 74851 860 74909 861
rect 75139 860 75197 861
rect 76675 860 76733 861
rect 65251 820 65260 860
rect 65300 820 70156 860
rect 70196 820 70205 860
rect 71406 820 71500 860
rect 71540 820 71549 860
rect 74286 820 74380 860
rect 74420 820 74860 860
rect 74900 820 74909 860
rect 75054 820 75148 860
rect 75188 820 75197 860
rect 76590 820 76684 860
rect 76724 820 76733 860
rect 78220 860 78260 903
rect 84163 860 84221 861
rect 78220 820 84172 860
rect 84212 820 84221 860
rect 17644 736 17740 776
rect 17780 736 17789 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 13699 735 13757 736
rect 16771 735 16829 736
rect 11203 692 11261 693
rect 14275 692 14333 693
rect 20140 692 20180 820
rect 26179 819 26237 820
rect 35107 819 35165 820
rect 36067 819 36125 820
rect 36451 819 36509 820
rect 20227 776 20285 777
rect 32227 776 32285 777
rect 35203 776 35261 777
rect 37780 776 37820 820
rect 54979 819 55037 820
rect 20227 736 20236 776
rect 20276 736 26284 776
rect 26324 736 32236 776
rect 32276 736 33620 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 35203 736 35212 776
rect 35252 736 37820 776
rect 40003 776 40061 777
rect 44323 776 44381 777
rect 45091 776 45149 777
rect 52483 776 52541 777
rect 64684 776 64724 820
rect 65251 819 65309 820
rect 70147 819 70205 820
rect 71491 819 71549 820
rect 74371 819 74429 820
rect 74851 819 74909 820
rect 75139 819 75197 820
rect 76675 819 76733 820
rect 84163 819 84221 820
rect 85219 860 85277 861
rect 89923 860 89981 861
rect 93292 860 93332 1072
rect 93388 1028 93428 1072
rect 93571 1071 93629 1072
rect 93955 1071 94013 1072
rect 94156 1028 94196 1072
rect 94723 1071 94781 1072
rect 94924 1072 95348 1112
rect 95491 1072 95500 1112
rect 95540 1072 95549 1112
rect 94924 1028 94964 1072
rect 95308 1028 95348 1072
rect 95788 1028 95828 1156
rect 96259 1112 96317 1113
rect 96643 1112 96701 1113
rect 99139 1112 99197 1113
rect 95875 1072 95884 1112
rect 95924 1072 96020 1112
rect 96174 1072 96268 1112
rect 96308 1072 96317 1112
rect 96558 1072 96652 1112
rect 96692 1072 96701 1112
rect 97027 1072 97036 1112
rect 97076 1072 97085 1112
rect 98659 1072 98668 1112
rect 98708 1072 98717 1112
rect 99054 1072 99148 1112
rect 99188 1072 99197 1112
rect 93388 988 93772 1028
rect 93812 988 94540 1028
rect 94580 988 94924 1028
rect 94964 988 94973 1028
rect 95020 988 95111 1028
rect 95151 988 95160 1028
rect 95299 988 95308 1028
rect 95348 988 95828 1028
rect 93859 904 93868 944
rect 93908 904 94156 944
rect 94196 904 94205 944
rect 94723 904 94732 944
rect 94772 904 94828 944
rect 94868 904 94877 944
rect 94531 860 94589 861
rect 95020 860 95060 988
rect 95203 904 95212 944
rect 95252 904 95261 944
rect 95395 904 95404 944
rect 95444 904 95692 944
rect 95732 904 95741 944
rect 85219 820 85228 860
rect 85268 820 85324 860
rect 85364 820 85373 860
rect 85603 820 85612 860
rect 85652 820 85661 860
rect 89923 820 89932 860
rect 89972 820 92468 860
rect 93292 820 93772 860
rect 93812 820 93821 860
rect 94446 820 94540 860
rect 94580 820 94589 860
rect 85219 819 85277 820
rect 40003 736 40012 776
rect 40052 736 44332 776
rect 44372 736 44381 776
rect 45006 736 45100 776
rect 45140 736 45149 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 50275 736 50284 776
rect 50324 736 50860 776
rect 50900 736 50909 776
rect 52398 736 52492 776
rect 52532 736 52541 776
rect 55555 736 55564 776
rect 55604 736 56044 776
rect 56084 736 56093 776
rect 56323 736 56332 776
rect 56372 736 57100 776
rect 57140 736 57149 776
rect 62572 736 63724 776
rect 63764 736 63773 776
rect 64675 736 64684 776
rect 64724 736 64733 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 20227 735 20285 736
rect 32227 735 32285 736
rect 5347 652 5356 692
rect 5396 652 11020 692
rect 11060 652 11069 692
rect 11203 652 11212 692
rect 11252 652 14132 692
rect 11203 651 11261 652
rect 14092 609 14132 652
rect 14275 652 14284 692
rect 14324 652 14476 692
rect 14516 652 14525 692
rect 15235 652 15244 692
rect 15284 652 20180 692
rect 14275 651 14333 652
rect 4195 608 4253 609
rect 10627 608 10685 609
rect 14083 608 14141 609
rect 20236 608 20276 735
rect 33580 692 33620 736
rect 35203 735 35261 736
rect 40003 735 40061 736
rect 44323 735 44381 736
rect 45091 735 45149 736
rect 52483 735 52541 736
rect 38467 692 38525 693
rect 43843 692 43901 693
rect 62572 692 62612 736
rect 25987 652 25996 692
rect 26036 652 26380 692
rect 26420 652 26429 692
rect 26755 652 26764 692
rect 26804 652 27148 692
rect 27188 652 27197 692
rect 27523 652 27532 692
rect 27572 652 27916 692
rect 27956 652 27965 692
rect 28291 652 28300 692
rect 28340 652 28684 692
rect 28724 652 28733 692
rect 29443 652 29452 692
rect 29492 652 29836 692
rect 29876 652 29885 692
rect 30211 652 30220 692
rect 30260 652 30604 692
rect 30644 652 30653 692
rect 31267 652 31276 692
rect 31316 652 31948 692
rect 31988 652 31997 692
rect 32899 652 32908 692
rect 32948 652 33484 692
rect 33524 652 33533 692
rect 33580 652 38476 692
rect 38516 652 43852 692
rect 43892 652 43901 692
rect 44131 652 44140 692
rect 44180 652 44428 692
rect 44468 652 44477 692
rect 44803 652 44812 692
rect 44852 652 45196 692
rect 45236 652 45245 692
rect 45571 652 45580 692
rect 45620 652 45964 692
rect 46004 652 46013 692
rect 46339 652 46348 692
rect 46388 652 46732 692
rect 46772 652 46781 692
rect 47107 652 47116 692
rect 47156 652 47500 692
rect 47540 652 47549 692
rect 47875 652 47884 692
rect 47924 652 48268 692
rect 48308 652 48317 692
rect 48643 652 48652 692
rect 48692 652 49036 692
rect 49076 652 49085 692
rect 49132 652 62612 692
rect 62659 692 62717 693
rect 66691 692 66749 693
rect 70156 692 70196 819
rect 72931 776 72989 777
rect 73603 776 73661 777
rect 79747 776 79805 777
rect 82819 776 82877 777
rect 83779 776 83837 777
rect 71875 736 71884 776
rect 71924 736 72172 776
rect 72212 736 72221 776
rect 72931 736 72940 776
rect 72980 736 73612 776
rect 73652 736 79756 776
rect 79796 736 79805 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 82734 736 82828 776
rect 82868 736 82877 776
rect 83694 736 83788 776
rect 83828 736 83837 776
rect 85612 776 85652 820
rect 89923 819 89981 820
rect 85612 736 85708 776
rect 85748 736 85757 776
rect 72931 735 72989 736
rect 73603 735 73661 736
rect 79747 735 79805 736
rect 82819 735 82877 736
rect 83779 735 83837 736
rect 70531 692 70589 693
rect 73027 692 73085 693
rect 85315 692 85373 693
rect 62659 652 62668 692
rect 62708 652 66700 692
rect 66740 652 66749 692
rect 67459 652 67468 692
rect 67508 652 67852 692
rect 67892 652 67901 692
rect 68611 652 68620 692
rect 68660 652 68908 692
rect 68948 652 68957 692
rect 70156 652 70540 692
rect 70580 652 70589 692
rect 38467 651 38525 652
rect 43843 651 43901 652
rect 4195 568 4204 608
rect 4244 568 4300 608
rect 4340 568 4349 608
rect 5059 568 5068 608
rect 5108 568 10636 608
rect 10676 568 10685 608
rect 4195 567 4253 568
rect 10627 567 10685 568
rect 10732 568 14036 608
rect 5827 524 5885 525
rect 6211 524 6269 525
rect 5742 484 5836 524
rect 5876 484 5885 524
rect 6126 484 6220 524
rect 6260 484 6269 524
rect 7651 484 7660 524
rect 7700 484 7948 524
rect 7988 484 7997 524
rect 8419 484 8428 524
rect 8468 484 8716 524
rect 8756 484 8765 524
rect 9187 484 9196 524
rect 9236 484 9484 524
rect 9524 484 9533 524
rect 9955 484 9964 524
rect 10004 484 10252 524
rect 10292 484 10301 524
rect 5827 483 5885 484
rect 6211 483 6269 484
rect 10732 440 10772 568
rect 13996 524 14036 568
rect 14083 568 14092 608
rect 14132 568 20276 608
rect 20995 608 21053 609
rect 28579 608 28637 609
rect 30691 608 30749 609
rect 32995 608 33053 609
rect 35395 608 35453 609
rect 41923 608 41981 609
rect 43939 608 43997 609
rect 20995 568 21004 608
rect 21044 568 27052 608
rect 27092 568 27101 608
rect 28494 568 28588 608
rect 28628 568 28637 608
rect 28771 568 28780 608
rect 28820 568 29356 608
rect 29396 568 29405 608
rect 30691 568 30700 608
rect 30740 568 30988 608
rect 31028 568 31037 608
rect 32995 568 33004 608
rect 33044 568 33100 608
rect 33140 568 33149 608
rect 34147 568 34156 608
rect 34196 568 34636 608
rect 34676 568 34685 608
rect 35260 568 35404 608
rect 35444 568 41588 608
rect 41838 568 41932 608
rect 41972 568 41981 608
rect 43854 568 43948 608
rect 43988 568 43997 608
rect 45283 568 45292 608
rect 45332 568 45484 608
rect 45524 568 45533 608
rect 14083 567 14141 568
rect 20995 567 21053 568
rect 28579 567 28637 568
rect 30691 567 30749 568
rect 32995 567 33053 568
rect 14851 524 14909 525
rect 11875 484 11884 524
rect 11924 484 12172 524
rect 12212 484 12221 524
rect 12643 484 12652 524
rect 12692 484 12940 524
rect 12980 484 12989 524
rect 13411 484 13420 524
rect 13460 484 13708 524
rect 13748 484 13757 524
rect 13996 484 14860 524
rect 14900 484 14909 524
rect 14851 483 14909 484
rect 15043 524 15101 525
rect 16483 524 16541 525
rect 19939 524 19997 525
rect 15043 484 15052 524
rect 15092 484 16492 524
rect 16532 484 16541 524
rect 17251 484 17260 524
rect 17300 484 17548 524
rect 17588 484 17597 524
rect 18403 484 18412 524
rect 18452 484 18700 524
rect 18740 484 18749 524
rect 19171 484 19180 524
rect 19220 484 19468 524
rect 19508 484 19517 524
rect 19854 484 19948 524
rect 19988 484 19997 524
rect 15043 483 15101 484
rect 16483 483 16541 484
rect 19939 483 19997 484
rect 20419 524 20477 525
rect 23875 524 23933 525
rect 26179 524 26237 525
rect 27619 524 27677 525
rect 27811 524 27869 525
rect 35260 524 35300 568
rect 35395 567 35453 568
rect 41548 525 41588 568
rect 41923 567 41981 568
rect 43939 567 43997 568
rect 41539 524 41597 525
rect 49132 524 49172 652
rect 62659 651 62717 652
rect 66691 651 66749 652
rect 70531 651 70589 652
rect 71308 652 73036 692
rect 73076 652 73085 692
rect 73219 652 73228 692
rect 73268 652 79372 692
rect 79412 652 85324 692
rect 85364 652 85373 692
rect 49219 608 49277 609
rect 49987 608 50045 609
rect 71308 608 71348 652
rect 73027 651 73085 652
rect 85315 651 85373 652
rect 85603 692 85661 693
rect 91075 692 91133 693
rect 92428 692 92468 820
rect 94531 819 94589 820
rect 94636 820 95060 860
rect 95212 860 95252 904
rect 95491 860 95549 861
rect 95788 860 95828 988
rect 95212 820 95500 860
rect 95540 820 95549 860
rect 95779 820 95788 860
rect 95828 820 95837 860
rect 94636 776 94676 820
rect 95491 819 95549 820
rect 94819 776 94877 777
rect 94627 736 94636 776
rect 94676 736 94685 776
rect 94819 736 94828 776
rect 94868 736 94962 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
rect 94819 735 94877 736
rect 95980 692 96020 1072
rect 96259 1071 96317 1072
rect 96643 1071 96701 1072
rect 85603 652 85612 692
rect 85652 652 90988 692
rect 91028 652 91084 692
rect 91124 652 91152 692
rect 92428 652 96020 692
rect 85603 651 85661 652
rect 91075 651 91133 652
rect 79843 608 79901 609
rect 83011 608 83069 609
rect 89155 608 89213 609
rect 94915 608 94973 609
rect 49219 568 49228 608
rect 49268 568 49940 608
rect 49219 567 49277 568
rect 49900 524 49940 568
rect 49987 568 49996 608
rect 50036 568 66796 608
rect 66836 568 66845 608
rect 67747 568 67756 608
rect 67796 568 71348 608
rect 71779 568 71788 608
rect 71828 568 77836 608
rect 77876 568 79400 608
rect 49987 567 50045 568
rect 62851 524 62909 525
rect 64675 524 64733 525
rect 70915 524 70973 525
rect 77251 524 77309 525
rect 79171 524 79229 525
rect 20419 484 20428 524
rect 20468 484 20620 524
rect 20660 484 20669 524
rect 21091 484 21100 524
rect 21140 484 21388 524
rect 21428 484 21437 524
rect 22627 484 22636 524
rect 22676 484 22924 524
rect 22964 484 22973 524
rect 23790 484 23884 524
rect 23924 484 23933 524
rect 25603 484 25612 524
rect 25652 484 25996 524
rect 26036 484 26045 524
rect 26179 484 26188 524
rect 26228 484 27628 524
rect 27668 484 27677 524
rect 27726 484 27820 524
rect 27860 484 27869 524
rect 29059 484 29068 524
rect 29108 484 29452 524
rect 29492 484 29501 524
rect 32323 484 32332 524
rect 32372 484 32908 524
rect 32948 484 32957 524
rect 33187 484 33196 524
rect 33236 484 33676 524
rect 33716 484 33725 524
rect 33859 484 33868 524
rect 33908 484 34444 524
rect 34484 484 34493 524
rect 34723 484 34732 524
rect 34772 484 35300 524
rect 35779 484 35788 524
rect 35828 484 36364 524
rect 36404 484 36413 524
rect 36547 484 36556 524
rect 36596 484 37132 524
rect 37172 484 37181 524
rect 37795 484 37804 524
rect 37844 484 38284 524
rect 38324 484 38333 524
rect 38563 484 38572 524
rect 38612 484 39052 524
rect 39092 484 39101 524
rect 40099 484 40108 524
rect 40148 484 40588 524
rect 40628 484 40637 524
rect 40867 484 40876 524
rect 40916 484 41356 524
rect 41396 484 41405 524
rect 41539 484 41548 524
rect 41588 484 43028 524
rect 43651 484 43660 524
rect 43700 484 44044 524
rect 44084 484 44093 524
rect 44236 484 44716 524
rect 44756 484 49172 524
rect 49411 484 49420 524
rect 49460 484 49804 524
rect 49844 484 49853 524
rect 49900 484 53548 524
rect 53588 484 53597 524
rect 53827 484 53836 524
rect 53876 484 54892 524
rect 54932 484 54941 524
rect 55843 484 55852 524
rect 55892 484 56332 524
rect 56372 484 56381 524
rect 62766 484 62860 524
rect 62900 484 62909 524
rect 63619 484 63628 524
rect 63668 484 63916 524
rect 63956 484 63965 524
rect 64579 484 64588 524
rect 64628 484 64684 524
rect 64724 484 64733 524
rect 65923 484 65932 524
rect 65972 484 66220 524
rect 66260 484 66269 524
rect 67843 484 67852 524
rect 67892 484 68140 524
rect 68180 484 68189 524
rect 68995 484 69004 524
rect 69044 484 69292 524
rect 69332 484 69341 524
rect 69763 484 69772 524
rect 69812 484 70060 524
rect 70100 484 70109 524
rect 70830 484 70924 524
rect 70964 484 70973 524
rect 71299 484 71308 524
rect 71348 484 71596 524
rect 71636 484 71645 524
rect 72451 484 72460 524
rect 72500 484 72748 524
rect 72788 484 72797 524
rect 73315 484 73324 524
rect 73364 484 73516 524
rect 73556 484 73565 524
rect 74371 484 74380 524
rect 74420 484 74668 524
rect 74708 484 74717 524
rect 75139 484 75148 524
rect 75188 484 75436 524
rect 75476 484 75485 524
rect 75907 484 75916 524
rect 75956 484 76204 524
rect 76244 484 76253 524
rect 76675 484 76684 524
rect 76724 484 76972 524
rect 77012 484 77021 524
rect 77166 484 77260 524
rect 77300 484 77309 524
rect 77443 484 77452 524
rect 77492 484 77740 524
rect 77780 484 77789 524
rect 78595 484 78604 524
rect 78644 484 78892 524
rect 78932 484 78941 524
rect 79086 484 79180 524
rect 79220 484 79229 524
rect 79360 524 79400 568
rect 79843 568 79852 608
rect 79892 568 79948 608
rect 79988 568 79997 608
rect 83011 568 83020 608
rect 83060 568 89164 608
rect 89204 568 94636 608
rect 94676 568 94685 608
rect 94915 568 94924 608
rect 94964 568 95308 608
rect 95348 568 95357 608
rect 79843 567 79901 568
rect 83011 567 83069 568
rect 89155 567 89213 568
rect 94915 567 94973 568
rect 97036 524 97076 1072
rect 97987 944 98045 945
rect 97902 904 97996 944
rect 98036 904 98045 944
rect 97987 903 98045 904
rect 98668 860 98708 1072
rect 99139 1071 99197 1072
rect 98179 820 98188 860
rect 98228 820 98708 860
rect 97219 776 97277 777
rect 97219 736 97228 776
rect 97268 736 97362 776
rect 97219 735 97277 736
rect 79360 484 83884 524
rect 83924 484 83933 524
rect 90979 484 90988 524
rect 91028 484 97076 524
rect 20419 483 20477 484
rect 23875 483 23933 484
rect 26179 483 26237 484
rect 27619 483 27677 484
rect 27811 483 27869 484
rect 41539 483 41597 484
rect 35011 440 35069 441
rect 35299 440 35357 441
rect 42988 440 43028 484
rect 43843 440 43901 441
rect 44236 440 44276 484
rect 62851 483 62909 484
rect 64675 483 64733 484
rect 70915 483 70973 484
rect 77251 483 77309 484
rect 79171 483 79229 484
rect 46243 440 46301 441
rect 85315 440 85373 441
rect 91459 440 91517 441
rect 3148 400 8620 440
rect 8660 400 10772 440
rect 11011 400 11020 440
rect 11060 400 11360 440
rect 11779 400 11788 440
rect 11828 400 18796 440
rect 18836 400 23980 440
rect 24020 400 30164 440
rect 32035 400 32044 440
rect 32084 400 32524 440
rect 32564 400 32573 440
rect 33571 400 33580 440
rect 33620 400 34060 440
rect 34100 400 34109 440
rect 34243 400 34252 440
rect 34292 400 34828 440
rect 34868 400 34877 440
rect 35011 400 35020 440
rect 35060 400 35154 440
rect 35299 400 35308 440
rect 35348 400 35404 440
rect 35444 400 35453 440
rect 36931 400 36940 440
rect 36980 400 37516 440
rect 37556 400 37565 440
rect 39331 400 39340 440
rect 39380 400 39820 440
rect 39860 400 39869 440
rect 41635 400 41644 440
rect 41684 400 42124 440
rect 42164 400 42173 440
rect 42403 400 42412 440
rect 42452 400 42892 440
rect 42932 400 42941 440
rect 42988 400 43796 440
rect 4771 356 4829 357
rect 10627 356 10685 357
rect 11320 356 11360 400
rect 30124 357 30164 400
rect 35011 399 35069 400
rect 35299 399 35357 400
rect 14851 356 14909 357
rect 20995 356 21053 357
rect 23779 356 23837 357
rect 29731 356 29789 357
rect 4675 316 4684 356
rect 4724 316 4780 356
rect 4820 316 4829 356
rect 6499 316 6508 356
rect 6548 316 6796 356
rect 6836 316 6845 356
rect 7564 316 10580 356
rect 4771 315 4829 316
rect 7564 272 7604 316
rect 5923 232 5932 272
rect 5972 232 7604 272
rect 7756 232 7852 272
rect 7892 232 7901 272
rect 6595 188 6653 189
rect 6510 148 6604 188
rect 6644 148 6653 188
rect 6595 147 6653 148
rect 7756 104 7796 232
rect 10540 188 10580 316
rect 10627 316 10636 356
rect 10676 316 11156 356
rect 11320 316 14804 356
rect 10627 315 10685 316
rect 11116 272 11156 316
rect 10723 232 10732 272
rect 10772 232 11020 272
rect 11060 232 11069 272
rect 11116 232 14572 272
rect 14612 232 14621 272
rect 14764 188 14804 316
rect 14851 316 14860 356
rect 14900 316 21004 356
rect 21044 316 21053 356
rect 21475 316 21484 356
rect 21524 316 21772 356
rect 21812 316 21821 356
rect 23779 316 23788 356
rect 23828 316 29740 356
rect 29780 316 29789 356
rect 14851 315 14909 316
rect 20995 315 21053 316
rect 23779 315 23837 316
rect 29731 315 29789 316
rect 30115 356 30173 357
rect 42403 356 42461 357
rect 43756 356 43796 400
rect 43843 400 43852 440
rect 43892 400 44276 440
rect 44323 400 44332 440
rect 44372 400 46252 440
rect 46292 400 65108 440
rect 65155 400 65164 440
rect 65204 400 65452 440
rect 65492 400 65501 440
rect 66307 400 66316 440
rect 66356 400 66604 440
rect 66644 400 66653 440
rect 66787 400 66796 440
rect 66836 400 73132 440
rect 73172 400 73181 440
rect 77827 400 77836 440
rect 77876 400 78124 440
rect 78164 400 78173 440
rect 78307 400 78316 440
rect 78356 400 78508 440
rect 78548 400 78557 440
rect 79084 400 81920 440
rect 43843 399 43901 400
rect 46243 399 46301 400
rect 47683 356 47741 357
rect 49987 356 50045 357
rect 65068 356 65108 400
rect 65443 356 65501 357
rect 72835 356 72893 357
rect 79084 356 79124 400
rect 81880 356 81920 400
rect 85315 400 85324 440
rect 85364 400 91468 440
rect 91508 400 97324 440
rect 97364 400 97373 440
rect 85315 399 85373 400
rect 91459 399 91517 400
rect 92611 356 92669 357
rect 30115 316 30124 356
rect 30164 316 36076 356
rect 36116 316 42412 356
rect 42452 316 42461 356
rect 43171 316 43180 356
rect 43220 316 43660 356
rect 43700 316 43709 356
rect 43756 316 47692 356
rect 47732 316 49996 356
rect 50036 316 50045 356
rect 54403 316 54412 356
rect 54452 316 55468 356
rect 55508 316 55517 356
rect 65068 316 65452 356
rect 65492 316 71788 356
rect 71828 316 71837 356
rect 72835 316 72844 356
rect 72884 316 79084 356
rect 79124 316 79133 356
rect 79363 316 79372 356
rect 79412 316 79660 356
rect 79700 316 79709 356
rect 80323 316 80332 356
rect 80372 316 80620 356
rect 80660 316 80669 356
rect 81880 316 85612 356
rect 85652 316 85661 356
rect 86179 316 86188 356
rect 86228 316 90740 356
rect 30115 315 30173 316
rect 42403 315 42461 316
rect 47683 315 47741 316
rect 49987 315 50045 316
rect 65443 315 65501 316
rect 72835 315 72893 316
rect 39235 272 39293 273
rect 45475 272 45533 273
rect 64579 272 64637 273
rect 76291 272 76349 273
rect 82243 272 82301 273
rect 14947 232 14956 272
rect 14996 232 15148 272
rect 15188 232 15197 272
rect 15331 232 15340 272
rect 15380 232 15628 272
rect 15668 232 15677 272
rect 16099 232 16108 272
rect 16148 232 16396 272
rect 16436 232 16445 272
rect 16492 232 16684 272
rect 16724 232 21812 272
rect 21859 232 21868 272
rect 21908 232 22156 272
rect 22196 232 22205 272
rect 23395 232 23404 272
rect 23444 232 23692 272
rect 23732 232 23741 272
rect 27043 232 27052 272
rect 27092 232 33004 272
rect 33044 232 39244 272
rect 39284 232 44120 272
rect 44515 232 44524 272
rect 44564 232 44812 272
rect 44852 232 44861 272
rect 44908 232 45484 272
rect 45524 232 64588 272
rect 64628 232 70828 272
rect 70868 232 70877 272
rect 73987 232 73996 272
rect 74036 232 74284 272
rect 74324 232 74333 272
rect 76291 232 76300 272
rect 76340 232 82252 272
rect 82292 232 82301 272
rect 90700 272 90740 316
rect 92611 316 92620 356
rect 92660 316 98476 356
rect 98516 316 98525 356
rect 92611 315 92669 316
rect 90700 232 92140 272
rect 92180 232 98092 272
rect 98132 232 98141 272
rect 16492 188 16532 232
rect 10540 148 11360 188
rect 11491 148 11500 188
rect 11540 148 11788 188
rect 11828 148 11837 188
rect 14764 148 16532 188
rect 16579 188 16637 189
rect 21772 188 21812 232
rect 39235 231 39293 232
rect 23299 188 23357 189
rect 44080 188 44120 232
rect 44908 188 44948 232
rect 45475 231 45533 232
rect 64579 231 64637 232
rect 76291 231 76349 232
rect 82243 231 82301 232
rect 70723 188 70781 189
rect 83011 188 83069 189
rect 16579 148 16588 188
rect 16628 148 21676 188
rect 21716 148 21725 188
rect 21772 148 23308 188
rect 23348 148 28780 188
rect 28820 148 28829 188
rect 29347 148 29356 188
rect 29396 148 34732 188
rect 34772 148 34781 188
rect 35107 148 35116 188
rect 35156 148 35596 188
rect 35636 148 35645 188
rect 44080 148 44948 188
rect 49123 148 49132 188
rect 49172 148 49420 188
rect 49460 148 49469 188
rect 53539 148 53548 188
rect 53588 148 60268 188
rect 60308 148 67756 188
rect 67796 148 67805 188
rect 70531 148 70540 188
rect 70580 148 70732 188
rect 70772 148 70781 188
rect 77155 148 77164 188
rect 77204 148 83020 188
rect 83060 148 83069 188
rect 11203 104 11261 105
rect 2500 64 11212 104
rect 11252 64 11261 104
rect 11320 104 11360 148
rect 16579 147 16637 148
rect 11491 104 11549 105
rect 15043 104 15101 105
rect 11320 64 11500 104
rect 11540 64 15052 104
rect 15092 64 15101 104
rect 11203 63 11261 64
rect 11491 63 11549 64
rect 15043 63 15101 64
rect 16771 104 16829 105
rect 19651 104 19709 105
rect 16771 64 16780 104
rect 16820 64 19660 104
rect 19700 64 19709 104
rect 16771 63 16829 64
rect 19651 63 19709 64
rect 19843 104 19901 105
rect 20131 104 20189 105
rect 19843 64 19852 104
rect 19892 64 19986 104
rect 20035 64 20044 104
rect 20084 64 20140 104
rect 20180 64 20189 104
rect 21676 104 21716 148
rect 23299 147 23357 148
rect 70723 147 70781 148
rect 83011 147 83069 148
rect 85699 188 85757 189
rect 91843 188 91901 189
rect 85699 148 85708 188
rect 85748 148 91852 188
rect 91892 148 97708 188
rect 97748 148 97757 188
rect 85699 147 85757 148
rect 91843 147 91901 148
rect 27811 104 27869 105
rect 64195 104 64253 105
rect 21676 64 27820 104
rect 27860 64 27869 104
rect 64110 64 64204 104
rect 64244 64 64253 104
rect 19843 63 19901 64
rect 20131 63 20189 64
rect 27811 63 27869 64
rect 64195 63 64253 64
rect 67267 104 67325 105
rect 72931 104 72989 105
rect 95491 104 95549 105
rect 67267 64 67276 104
rect 67316 64 72940 104
rect 72980 64 72989 104
rect 95107 64 95116 104
rect 95156 64 95500 104
rect 95540 64 95549 104
rect 67267 63 67325 64
rect 72931 63 72989 64
rect 95491 63 95549 64
<< via3 >>
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 42220 5188 42260 5228
rect 46060 5104 46100 5144
rect 55372 5104 55412 5144
rect 50380 4936 50420 4976
rect 48364 4768 48404 4808
rect 48940 4768 48980 4808
rect 62380 4684 62420 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 38668 4348 38708 4388
rect 52108 4348 52148 4388
rect 52492 4348 52532 4388
rect 66796 4348 66836 4388
rect 28012 4264 28052 4304
rect 38956 4180 38996 4220
rect 68524 4180 68564 4220
rect 46060 4096 46100 4136
rect 58636 4096 58676 4136
rect 66508 4096 66548 4136
rect 26092 4012 26132 4052
rect 48940 4012 48980 4052
rect 39244 3928 39284 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 35692 3760 35732 3800
rect 44620 3760 44660 3800
rect 46060 3760 46100 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 58444 3760 58484 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 38092 3676 38132 3716
rect 47596 3676 47636 3716
rect 55372 3676 55412 3716
rect 32236 3592 32276 3632
rect 90700 3592 90740 3632
rect 9580 3508 9620 3548
rect 41356 3508 41396 3548
rect 47884 3508 47924 3548
rect 69196 3508 69236 3548
rect 69772 3508 69812 3548
rect 71308 3508 71348 3548
rect 5932 3424 5972 3464
rect 6892 3424 6932 3464
rect 11116 3424 11156 3464
rect 11500 3424 11540 3464
rect 13036 3424 13076 3464
rect 17164 3424 17204 3464
rect 17548 3424 17588 3464
rect 18700 3424 18740 3464
rect 19948 3424 19988 3464
rect 23788 3424 23828 3464
rect 25324 3424 25364 3464
rect 29836 3424 29876 3464
rect 36844 3424 36884 3464
rect 50380 3424 50420 3464
rect 65836 3424 65876 3464
rect 66220 3424 66260 3464
rect 72844 3424 72884 3464
rect 79180 3424 79220 3464
rect 80332 3424 80372 3464
rect 84556 3424 84596 3464
rect 92812 3424 92852 3464
rect 54316 3340 54356 3380
rect 64684 3340 64724 3380
rect 72460 3340 72500 3380
rect 15820 3256 15860 3296
rect 66988 3256 67028 3296
rect 4204 3172 4244 3212
rect 31756 3172 31796 3212
rect 34348 3172 34388 3212
rect 38092 3172 38132 3212
rect 55084 3172 55124 3212
rect 65356 3172 65396 3212
rect 72940 3172 72980 3212
rect 83788 3172 83828 3212
rect 41932 3088 41972 3128
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 35308 3004 35348 3044
rect 42220 3004 42260 3044
rect 46156 3004 46196 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 54988 2920 55028 2960
rect 65836 2920 65876 2960
rect 20140 2836 20180 2876
rect 44044 2836 44084 2876
rect 45004 2836 45044 2876
rect 91468 2836 91508 2876
rect 92812 2836 92852 2876
rect 20044 2752 20084 2792
rect 54892 2752 54932 2792
rect 64684 2752 64724 2792
rect 74764 2752 74804 2792
rect 84748 2752 84788 2792
rect 84940 2752 84980 2792
rect 14284 2668 14324 2708
rect 48076 2668 48116 2708
rect 61324 2668 61364 2708
rect 2284 2584 2324 2624
rect 3916 2584 3956 2624
rect 7180 2584 7220 2624
rect 8044 2584 8084 2624
rect 12748 2584 12788 2624
rect 20044 2584 20084 2624
rect 20428 2584 20468 2624
rect 21868 2584 21908 2624
rect 23404 2584 23444 2624
rect 26572 2584 26612 2624
rect 28108 2584 28148 2624
rect 29548 2584 29588 2624
rect 30892 2584 30932 2624
rect 31660 2584 31700 2624
rect 33772 2584 33812 2624
rect 38764 2584 38804 2624
rect 40204 2584 40244 2624
rect 41836 2584 41876 2624
rect 42220 2584 42260 2624
rect 42988 2584 43028 2624
rect 46540 2584 46580 2624
rect 6604 2500 6644 2540
rect 19948 2416 19988 2456
rect 20428 2332 20468 2372
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 41932 2500 41972 2540
rect 42316 2500 42356 2540
rect 48460 2584 48500 2624
rect 48364 2500 48404 2540
rect 49324 2584 49364 2624
rect 54892 2616 54932 2624
rect 54892 2584 54932 2616
rect 72940 2668 72980 2708
rect 58636 2584 58676 2624
rect 61708 2584 61748 2624
rect 63532 2584 63572 2624
rect 64012 2584 64052 2624
rect 75628 2584 75668 2624
rect 55468 2416 55508 2456
rect 59116 2416 59156 2456
rect 35308 2332 35348 2372
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 35596 2332 35636 2372
rect 76876 2584 76916 2624
rect 74284 2500 74324 2540
rect 77260 2500 77300 2540
rect 64300 2416 64340 2456
rect 66604 2416 66644 2456
rect 85324 2668 85364 2708
rect 88012 2668 88052 2708
rect 93676 2668 93716 2708
rect 78604 2584 78644 2624
rect 81484 2584 81524 2624
rect 83404 2584 83444 2624
rect 86476 2584 86516 2624
rect 85228 2500 85268 2540
rect 84556 2416 84596 2456
rect 89548 2584 89588 2624
rect 95116 2584 95156 2624
rect 96364 2584 96404 2624
rect 96748 2584 96788 2624
rect 97132 2584 97172 2624
rect 91084 2500 91124 2540
rect 97996 2500 98036 2540
rect 84748 2416 84788 2456
rect 93868 2332 93908 2372
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 19948 2164 19988 2204
rect 32236 2164 32276 2204
rect 55564 2248 55604 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 58444 1996 58484 2036
rect 69196 1996 69236 2036
rect 6892 1912 6932 1952
rect 19372 1912 19412 1952
rect 24844 1912 24884 1952
rect 50380 1912 50420 1952
rect 51436 1912 51476 1952
rect 52108 1912 52148 1952
rect 62572 1912 62612 1952
rect 64588 1912 64628 1952
rect 67852 1912 67892 1952
rect 37324 1828 37364 1868
rect 79948 1828 79988 1868
rect 55468 1660 55508 1700
rect 55948 1660 55988 1700
rect 64012 1660 64052 1700
rect 42316 1576 42356 1616
rect 55084 1576 55124 1616
rect 71308 1576 71348 1616
rect 79852 1576 79892 1616
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 20428 1492 20468 1532
rect 23884 1492 23924 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 55468 1492 55508 1532
rect 6412 1408 6452 1448
rect 11212 1408 11252 1448
rect 33004 1408 33044 1448
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 70732 1492 70772 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 79756 1492 79796 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 94828 1492 94868 1532
rect 97228 1492 97268 1532
rect 35116 1408 35156 1448
rect 5836 1324 5876 1364
rect 14284 1324 14324 1364
rect 4780 1240 4820 1280
rect 6220 1240 6260 1280
rect 35308 1408 35348 1448
rect 44332 1408 44372 1448
rect 69388 1408 69428 1448
rect 30700 1324 30740 1364
rect 51436 1324 51476 1364
rect 62860 1324 62900 1364
rect 16780 1240 16820 1280
rect 17548 1240 17588 1280
rect 19276 1240 19316 1280
rect 7180 1156 7220 1196
rect 7564 1156 7604 1196
rect 8332 1156 8372 1196
rect 13324 1156 13364 1196
rect 14092 1156 14132 1196
rect 14860 1156 14900 1196
rect 18316 1156 18356 1196
rect 19948 1156 19988 1196
rect 1228 1072 1268 1112
rect 1612 1072 1652 1112
rect 1996 1072 2036 1112
rect 2764 1072 2804 1112
rect 4300 1072 4340 1112
rect 4684 1072 4724 1112
rect 6508 1072 6548 1112
rect 9868 1072 9908 1112
rect 10252 1072 10292 1112
rect 10636 1072 10676 1112
rect 20236 1156 20276 1196
rect 21004 1156 21044 1196
rect 22540 1156 22580 1196
rect 23308 1156 23348 1196
rect 24460 1156 24500 1196
rect 11500 1072 11540 1112
rect 12268 1072 12308 1112
rect 12556 1072 12596 1112
rect 12940 1072 12980 1112
rect 16012 1072 16052 1112
rect 22156 1072 22196 1112
rect 23788 1072 23828 1112
rect 16396 988 16436 1028
rect 6412 904 6452 944
rect 6892 904 6932 944
rect 16588 904 16628 944
rect 17548 904 17588 944
rect 12076 820 12116 860
rect 14380 820 14420 860
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 13708 736 13748 776
rect 16780 736 16820 776
rect 18700 988 18740 1028
rect 19372 988 19412 1028
rect 20620 988 20660 1028
rect 22924 988 22964 1028
rect 24844 1072 24884 1112
rect 26188 1240 26228 1280
rect 32620 1240 32660 1280
rect 35116 1240 35156 1280
rect 26668 1156 26708 1196
rect 28204 1156 28244 1196
rect 25516 1072 25556 1112
rect 29740 1072 29780 1112
rect 30124 1072 30164 1112
rect 25900 988 25940 1028
rect 27628 988 27668 1028
rect 31852 1156 31892 1196
rect 32236 1156 32276 1196
rect 34156 1156 34196 1196
rect 38476 1156 38516 1196
rect 38860 1156 38900 1196
rect 39244 1156 39284 1196
rect 39628 1240 39668 1280
rect 49228 1240 49268 1280
rect 49516 1240 49556 1280
rect 40012 1156 40052 1196
rect 40396 1156 40436 1196
rect 31084 1072 31124 1112
rect 31468 1072 31508 1112
rect 34540 1072 34580 1112
rect 35020 1072 35060 1112
rect 42700 1156 42740 1196
rect 44428 1156 44468 1196
rect 46252 1156 46292 1196
rect 47788 1156 47828 1196
rect 35404 1072 35444 1112
rect 37036 1072 37076 1112
rect 37324 1072 37364 1112
rect 40780 1072 40820 1112
rect 41548 1072 41588 1112
rect 42412 1072 42452 1112
rect 73036 1408 73076 1448
rect 81484 1408 81524 1448
rect 88396 1408 88436 1448
rect 94924 1408 94964 1448
rect 64204 1324 64244 1364
rect 64684 1324 64724 1364
rect 65260 1324 65300 1364
rect 66892 1324 66932 1364
rect 71500 1324 71540 1364
rect 72268 1324 72308 1364
rect 48076 1156 48116 1196
rect 49708 1156 49748 1196
rect 62764 1156 62804 1196
rect 63532 1156 63572 1196
rect 67276 1156 67316 1196
rect 68044 1156 68084 1196
rect 72844 1240 72884 1280
rect 69772 1156 69812 1196
rect 70156 1156 70196 1196
rect 70444 1156 70484 1196
rect 72076 1156 72116 1196
rect 72460 1156 72500 1196
rect 72940 1156 72980 1196
rect 73612 1156 73652 1196
rect 80524 1324 80564 1364
rect 82828 1324 82868 1364
rect 85324 1324 85364 1364
rect 75532 1240 75572 1280
rect 79180 1240 79220 1280
rect 81100 1240 81140 1280
rect 85708 1240 85748 1280
rect 87628 1240 87668 1280
rect 88780 1324 88820 1364
rect 89932 1240 89972 1280
rect 90316 1240 90356 1280
rect 92620 1240 92660 1280
rect 93196 1240 93236 1280
rect 94540 1240 94580 1280
rect 86956 1156 86996 1196
rect 88012 1156 88052 1196
rect 89164 1156 89204 1196
rect 89548 1156 89588 1196
rect 43276 1072 43316 1112
rect 43564 1072 43604 1112
rect 47020 1072 47060 1112
rect 34060 988 34100 1028
rect 34252 988 34292 1028
rect 39628 988 39668 1028
rect 30508 904 30548 944
rect 31756 904 31796 944
rect 42028 988 42068 1028
rect 47692 1072 47732 1112
rect 48940 1072 48980 1112
rect 49132 1072 49172 1112
rect 51436 1072 51476 1112
rect 55948 1072 55988 1112
rect 62668 1072 62708 1112
rect 62956 1072 62996 1112
rect 64300 1072 64340 1112
rect 64588 1072 64628 1112
rect 65452 1072 65492 1112
rect 65740 1072 65780 1112
rect 66796 1072 66836 1112
rect 68620 1072 68660 1112
rect 68812 1072 68852 1112
rect 74764 1072 74804 1112
rect 75916 1072 75956 1112
rect 76300 1072 76340 1112
rect 46636 988 46676 1028
rect 71308 988 71348 1028
rect 81868 1072 81908 1112
rect 82252 1072 82292 1112
rect 82636 1072 82676 1112
rect 83020 1072 83060 1112
rect 84172 1072 84212 1112
rect 84556 1072 84596 1112
rect 85612 1072 85652 1112
rect 86476 1072 86516 1112
rect 86860 1072 86900 1112
rect 91084 1072 91124 1112
rect 91468 1072 91508 1112
rect 91852 1072 91892 1112
rect 93004 1072 93044 1112
rect 93580 1072 93620 1112
rect 93964 1072 94004 1112
rect 94732 1072 94772 1112
rect 45484 904 45524 944
rect 62956 904 62996 944
rect 64012 904 64052 944
rect 65356 904 65396 944
rect 66892 904 66932 944
rect 70924 904 70964 944
rect 72268 904 72308 944
rect 78220 904 78260 944
rect 78604 988 78644 1028
rect 89548 988 89588 1028
rect 90700 988 90740 1028
rect 92044 988 92084 1028
rect 82252 904 82292 944
rect 88396 904 88436 944
rect 20044 820 20084 860
rect 26188 820 26228 860
rect 35116 820 35156 860
rect 36076 820 36116 860
rect 36460 820 36500 860
rect 54988 820 55028 860
rect 65260 820 65300 860
rect 70156 820 70196 860
rect 71500 820 71540 860
rect 74380 820 74420 860
rect 74860 820 74900 860
rect 75148 820 75188 860
rect 76684 820 76724 860
rect 84172 820 84212 860
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 20236 736 20276 776
rect 32236 736 32276 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 35212 736 35252 776
rect 96268 1072 96308 1112
rect 96652 1072 96692 1112
rect 99148 1072 99188 1112
rect 85228 820 85268 860
rect 89932 820 89972 860
rect 94540 820 94580 860
rect 40012 736 40052 776
rect 44332 736 44372 776
rect 45100 736 45140 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 52492 736 52532 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 11212 652 11252 692
rect 14284 652 14324 692
rect 38476 652 38516 692
rect 43852 652 43892 692
rect 72940 736 72980 776
rect 73612 736 73652 776
rect 79756 736 79796 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 82828 736 82868 776
rect 83788 736 83828 776
rect 62668 652 62708 692
rect 66700 652 66740 692
rect 70540 652 70580 692
rect 4204 568 4244 608
rect 10636 568 10676 608
rect 5836 484 5876 524
rect 6220 484 6260 524
rect 14092 568 14132 608
rect 21004 568 21044 608
rect 28588 568 28628 608
rect 30700 568 30740 608
rect 33004 568 33044 608
rect 35404 568 35444 608
rect 41932 568 41972 608
rect 43948 568 43988 608
rect 14860 484 14900 524
rect 15052 484 15092 524
rect 16492 484 16532 524
rect 19948 484 19988 524
rect 73036 652 73076 692
rect 85324 652 85364 692
rect 95500 820 95540 860
rect 94828 736 94868 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
rect 85612 652 85652 692
rect 91084 652 91124 692
rect 49228 568 49268 608
rect 49996 568 50036 608
rect 20428 484 20468 524
rect 23884 484 23924 524
rect 26188 484 26228 524
rect 27628 484 27668 524
rect 27820 484 27860 524
rect 41548 484 41588 524
rect 62860 484 62900 524
rect 64684 484 64724 524
rect 70924 484 70964 524
rect 77260 484 77300 524
rect 79180 484 79220 524
rect 79852 568 79892 608
rect 83020 568 83060 608
rect 89164 568 89204 608
rect 94924 568 94964 608
rect 97996 904 98036 944
rect 97228 736 97268 776
rect 35020 400 35060 440
rect 35308 400 35348 440
rect 4780 316 4820 356
rect 6604 148 6644 188
rect 10636 316 10676 356
rect 14860 316 14900 356
rect 21004 316 21044 356
rect 23788 316 23828 356
rect 29740 316 29780 356
rect 43852 400 43892 440
rect 46252 400 46292 440
rect 85324 400 85364 440
rect 91468 400 91508 440
rect 30124 316 30164 356
rect 42412 316 42452 356
rect 47692 316 47732 356
rect 49996 316 50036 356
rect 65452 316 65492 356
rect 72844 316 72884 356
rect 39244 232 39284 272
rect 45484 232 45524 272
rect 64588 232 64628 272
rect 76300 232 76340 272
rect 82252 232 82292 272
rect 92620 316 92660 356
rect 16588 148 16628 188
rect 23308 148 23348 188
rect 70732 148 70772 188
rect 83020 148 83060 188
rect 11212 64 11252 104
rect 11500 64 11540 104
rect 15052 64 15092 104
rect 16780 64 16820 104
rect 19660 64 19700 104
rect 19852 64 19892 104
rect 20140 64 20180 104
rect 85708 148 85748 188
rect 91852 148 91892 188
rect 27820 64 27860 104
rect 64204 64 64244 104
rect 67276 64 67316 104
rect 72940 64 72980 104
rect 95500 64 95540 104
<< metal4 >>
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 42220 5228 42260 5237
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 38668 4388 38708 4397
rect 28012 4304 28052 4313
rect 26091 4136 26133 4145
rect 26091 4096 26092 4136
rect 26132 4096 26133 4136
rect 26091 4087 26133 4096
rect 26092 4052 26132 4087
rect 28012 4061 28052 4264
rect 26092 4001 26132 4012
rect 28011 4052 28053 4061
rect 28011 4012 28012 4052
rect 28052 4012 28053 4052
rect 28011 4003 28053 4012
rect 38668 3977 38708 4348
rect 38955 4220 38997 4229
rect 38955 4180 38956 4220
rect 38996 4180 38997 4220
rect 38955 4171 38997 4180
rect 38956 4086 38996 4171
rect 38667 3968 38709 3977
rect 38667 3928 38668 3968
rect 38708 3928 38709 3968
rect 38667 3919 38709 3928
rect 39244 3968 39284 3977
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 35692 3800 35732 3809
rect 11115 3716 11157 3725
rect 11115 3676 11116 3716
rect 11156 3676 11157 3716
rect 11115 3667 11157 3676
rect 17163 3716 17205 3725
rect 17163 3676 17164 3716
rect 17204 3676 17205 3716
rect 17163 3667 17205 3676
rect 9579 3548 9621 3557
rect 9579 3508 9580 3548
rect 9620 3508 9621 3548
rect 9579 3499 9621 3508
rect 5931 3464 5973 3473
rect 5931 3424 5932 3464
rect 5972 3424 5973 3464
rect 5931 3415 5973 3424
rect 6892 3464 6932 3473
rect 5932 3330 5972 3415
rect 6892 3221 6932 3424
rect 4204 3212 4244 3221
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 2283 2624 2325 2633
rect 2283 2584 2284 2624
rect 2324 2584 2325 2624
rect 2283 2575 2325 2584
rect 3915 2624 3957 2633
rect 3915 2584 3916 2624
rect 3956 2584 3957 2624
rect 3915 2575 3957 2584
rect 2284 2490 2324 2575
rect 3916 2490 3956 2575
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 1228 1112 1268 1121
rect 1228 953 1268 1072
rect 1612 1112 1652 1121
rect 1227 944 1269 953
rect 1227 904 1228 944
rect 1268 904 1269 944
rect 1227 895 1269 904
rect 1612 617 1652 1072
rect 1995 1112 2037 1121
rect 1995 1072 1996 1112
rect 2036 1072 2037 1112
rect 1995 1063 2037 1072
rect 2763 1112 2805 1121
rect 2763 1072 2764 1112
rect 2804 1072 2805 1112
rect 2763 1063 2805 1072
rect 1996 978 2036 1063
rect 2764 978 2804 1063
rect 1611 608 1653 617
rect 1611 568 1612 608
rect 1652 568 1653 608
rect 1611 559 1653 568
rect 4204 608 4244 3172
rect 6891 3212 6933 3221
rect 6891 3172 6892 3212
rect 6932 3172 6933 3212
rect 6891 3163 6933 3172
rect 6604 2540 6644 2549
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 6412 1448 6452 1457
rect 5836 1364 5876 1373
rect 4780 1280 4820 1289
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 4684 1112 4724 1121
rect 4300 978 4340 1063
rect 4684 953 4724 1072
rect 4683 944 4725 953
rect 4683 904 4684 944
rect 4724 904 4725 944
rect 4683 895 4725 904
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 4204 559 4244 568
rect 4780 356 4820 1240
rect 5836 524 5876 1324
rect 5836 475 5876 484
rect 6220 1280 6260 1289
rect 6220 524 6260 1240
rect 6412 944 6452 1408
rect 6412 895 6452 904
rect 6508 1112 6548 1121
rect 6508 869 6548 1072
rect 6507 860 6549 869
rect 6507 820 6508 860
rect 6548 820 6549 860
rect 6507 811 6549 820
rect 6220 475 6260 484
rect 4780 307 4820 316
rect 6604 188 6644 2500
rect 6892 1952 6932 3163
rect 8043 2708 8085 2717
rect 8043 2668 8044 2708
rect 8084 2668 8085 2708
rect 8043 2659 8085 2668
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 8044 2624 8084 2659
rect 7180 2490 7220 2575
rect 8044 2573 8084 2584
rect 9580 2549 9620 3499
rect 11116 3464 11156 3667
rect 15819 3548 15861 3557
rect 15819 3508 15820 3548
rect 15860 3508 15861 3548
rect 15819 3499 15861 3508
rect 11116 3415 11156 3424
rect 11500 3464 11540 3475
rect 11500 3389 11540 3424
rect 13036 3464 13076 3473
rect 11499 3380 11541 3389
rect 11499 3340 11500 3380
rect 11540 3340 11541 3380
rect 11499 3331 11541 3340
rect 13036 3221 13076 3424
rect 15820 3296 15860 3499
rect 13035 3212 13077 3221
rect 13035 3172 13036 3212
rect 13076 3172 13077 3212
rect 13035 3163 13077 3172
rect 12748 2633 12788 2718
rect 15820 2717 15860 3256
rect 17164 3464 17204 3667
rect 32236 3632 32276 3641
rect 19371 3548 19413 3557
rect 19371 3508 19372 3548
rect 19412 3508 19413 3548
rect 19371 3499 19413 3508
rect 25323 3548 25365 3557
rect 25323 3508 25324 3548
rect 25364 3508 25365 3548
rect 25323 3499 25365 3508
rect 31659 3548 31701 3557
rect 31659 3508 31660 3548
rect 31700 3508 31701 3548
rect 31659 3499 31701 3508
rect 17164 2885 17204 3424
rect 17548 3464 17588 3475
rect 17548 3389 17588 3424
rect 18700 3464 18740 3473
rect 17547 3380 17589 3389
rect 17547 3340 17548 3380
rect 17588 3340 17589 3380
rect 17547 3331 17589 3340
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 18700 2969 18740 3424
rect 19372 3221 19412 3499
rect 19948 3464 19988 3473
rect 19371 3212 19413 3221
rect 19371 3172 19372 3212
rect 19412 3172 19413 3212
rect 19371 3163 19413 3172
rect 18699 2960 18741 2969
rect 18699 2920 18700 2960
rect 18740 2920 18741 2960
rect 18699 2911 18741 2920
rect 17163 2876 17205 2885
rect 17163 2836 17164 2876
rect 17204 2836 17205 2876
rect 17163 2827 17205 2836
rect 14283 2708 14325 2717
rect 14283 2668 14284 2708
rect 14324 2668 14325 2708
rect 14283 2659 14325 2668
rect 15819 2708 15861 2717
rect 15819 2668 15820 2708
rect 15860 2668 15861 2708
rect 15819 2659 15861 2668
rect 12747 2624 12789 2633
rect 12747 2584 12748 2624
rect 12788 2584 12789 2624
rect 12747 2575 12789 2584
rect 14284 2574 14324 2659
rect 18700 2633 18740 2911
rect 18699 2624 18741 2633
rect 18699 2584 18700 2624
rect 18740 2584 18741 2624
rect 18699 2575 18741 2584
rect 9579 2540 9621 2549
rect 9579 2500 9580 2540
rect 9620 2500 9621 2540
rect 9579 2491 9621 2500
rect 6892 1903 6932 1912
rect 19372 1952 19412 3163
rect 19948 2456 19988 3424
rect 23788 3464 23828 3475
rect 23788 3389 23828 3424
rect 25324 3464 25364 3499
rect 25324 3413 25364 3424
rect 29836 3464 29876 3475
rect 29836 3389 29876 3424
rect 23787 3380 23829 3389
rect 23787 3340 23788 3380
rect 23828 3340 23829 3380
rect 23787 3331 23829 3340
rect 29835 3380 29877 3389
rect 29835 3340 29836 3380
rect 29876 3340 29877 3380
rect 29835 3331 29877 3340
rect 24843 2960 24885 2969
rect 24843 2920 24844 2960
rect 24884 2920 24885 2960
rect 24843 2911 24885 2920
rect 20140 2876 20180 2885
rect 20044 2792 20084 2801
rect 20044 2624 20084 2752
rect 20044 2575 20084 2584
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 19948 2204 19988 2416
rect 19948 2155 19988 2164
rect 19372 1903 19412 1912
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 11212 1448 11252 1457
rect 7563 1364 7605 1373
rect 7563 1324 7564 1364
rect 7604 1324 7605 1364
rect 7563 1315 7605 1324
rect 6891 1280 6933 1289
rect 6891 1240 6892 1280
rect 6932 1240 6933 1280
rect 6891 1231 6933 1240
rect 6892 1037 6932 1231
rect 7180 1196 7220 1205
rect 6891 1028 6933 1037
rect 6891 988 6892 1028
rect 6932 988 6933 1028
rect 6891 979 6933 988
rect 6892 944 6932 979
rect 6892 894 6932 904
rect 7180 617 7220 1156
rect 7564 1196 7604 1315
rect 10059 1280 10101 1289
rect 10059 1240 10060 1280
rect 10100 1240 10101 1280
rect 10059 1231 10101 1240
rect 7564 785 7604 1156
rect 8331 1196 8373 1205
rect 8331 1156 8332 1196
rect 8372 1156 8373 1196
rect 8331 1147 8373 1156
rect 8332 1037 8372 1147
rect 10060 1121 10100 1231
rect 9867 1112 9909 1121
rect 9867 1072 9868 1112
rect 9908 1072 9909 1112
rect 9867 1063 9909 1072
rect 10059 1112 10101 1121
rect 10059 1072 10060 1112
rect 10100 1072 10101 1112
rect 10059 1063 10101 1072
rect 10252 1112 10292 1121
rect 8331 1028 8373 1037
rect 8331 988 8332 1028
rect 8372 988 8373 1028
rect 8331 979 8373 988
rect 9868 978 9908 1063
rect 10252 953 10292 1072
rect 10636 1112 10676 1121
rect 10251 944 10293 953
rect 10251 904 10252 944
rect 10292 904 10293 944
rect 10251 895 10293 904
rect 7563 776 7605 785
rect 7563 736 7564 776
rect 7604 736 7605 776
rect 7563 727 7605 736
rect 7179 608 7221 617
rect 7179 568 7180 608
rect 7220 568 7221 608
rect 7179 559 7221 568
rect 10636 608 10676 1072
rect 11212 953 11252 1408
rect 14284 1364 14324 1373
rect 11403 1280 11445 1289
rect 11403 1240 11404 1280
rect 11444 1240 11445 1280
rect 11403 1231 11445 1240
rect 12555 1280 12597 1289
rect 12555 1240 12556 1280
rect 12596 1240 12597 1280
rect 12555 1231 12597 1240
rect 11404 953 11444 1231
rect 11500 1112 11540 1121
rect 11211 944 11253 953
rect 11211 904 11212 944
rect 11252 904 11253 944
rect 11211 895 11253 904
rect 11403 944 11445 953
rect 11403 904 11404 944
rect 11444 904 11445 944
rect 11403 895 11445 904
rect 10636 356 10676 568
rect 10636 307 10676 316
rect 11212 692 11252 701
rect 6604 139 6644 148
rect 11212 104 11252 652
rect 11212 55 11252 64
rect 11500 104 11540 1072
rect 12268 1112 12308 1123
rect 12268 1037 12308 1072
rect 12556 1112 12596 1231
rect 13324 1196 13364 1205
rect 12556 1063 12596 1072
rect 12939 1112 12981 1121
rect 12939 1072 12940 1112
rect 12980 1072 12981 1112
rect 12939 1063 12981 1072
rect 12075 1028 12117 1037
rect 12075 988 12076 1028
rect 12116 988 12117 1028
rect 12075 979 12117 988
rect 12267 1028 12309 1037
rect 12267 988 12268 1028
rect 12308 988 12309 1028
rect 12267 979 12309 988
rect 12076 860 12116 979
rect 12940 978 12980 1063
rect 12076 811 12116 820
rect 13324 449 13364 1156
rect 14092 1196 14132 1205
rect 13707 776 13749 785
rect 13707 736 13708 776
rect 13748 736 13749 776
rect 13707 727 13749 736
rect 13708 642 13748 727
rect 14092 608 14132 1156
rect 14284 692 14324 1324
rect 16780 1280 16820 1289
rect 14860 1196 14900 1205
rect 14284 643 14324 652
rect 14380 860 14420 869
rect 14092 559 14132 568
rect 13323 440 13365 449
rect 13323 400 13324 440
rect 13364 400 13365 440
rect 13323 391 13365 400
rect 14380 281 14420 820
rect 14860 524 14900 1156
rect 16011 1196 16053 1205
rect 16011 1156 16012 1196
rect 16052 1156 16053 1196
rect 16011 1147 16053 1156
rect 16012 1112 16052 1147
rect 16012 1061 16052 1072
rect 16396 1028 16436 1037
rect 16396 617 16436 988
rect 16491 944 16533 953
rect 16491 904 16492 944
rect 16532 904 16533 944
rect 16491 895 16533 904
rect 16588 944 16628 953
rect 16395 608 16437 617
rect 16395 568 16396 608
rect 16436 568 16437 608
rect 16395 559 16437 568
rect 14860 356 14900 484
rect 14860 307 14900 316
rect 15052 524 15092 533
rect 14379 272 14421 281
rect 14379 232 14380 272
rect 14420 232 14421 272
rect 14379 223 14421 232
rect 11500 55 11540 64
rect 15052 104 15092 484
rect 16492 524 16532 895
rect 16492 475 16532 484
rect 16588 188 16628 904
rect 16588 139 16628 148
rect 16780 776 16820 1240
rect 17548 1280 17588 1289
rect 17548 1121 17588 1240
rect 18699 1280 18741 1289
rect 18699 1240 18700 1280
rect 18740 1240 18741 1280
rect 18699 1231 18741 1240
rect 19276 1280 19316 1289
rect 18316 1196 18356 1207
rect 18316 1121 18356 1156
rect 17547 1112 17589 1121
rect 17547 1072 17548 1112
rect 17588 1072 17589 1112
rect 17547 1063 17589 1072
rect 18315 1112 18357 1121
rect 18315 1072 18316 1112
rect 18356 1072 18357 1112
rect 18315 1063 18357 1072
rect 18700 1028 18740 1231
rect 18700 979 18740 988
rect 17547 944 17589 953
rect 17547 904 17548 944
rect 17588 904 17589 944
rect 17547 895 17589 904
rect 17548 810 17588 895
rect 15052 55 15092 64
rect 16780 104 16820 736
rect 19276 449 19316 1240
rect 19948 1196 19988 1205
rect 19372 1028 19412 1037
rect 19372 785 19412 988
rect 19371 776 19413 785
rect 19371 736 19372 776
rect 19412 736 19413 776
rect 19371 727 19413 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 19948 524 19988 1156
rect 19948 475 19988 484
rect 20044 860 20084 869
rect 19275 440 19317 449
rect 19275 400 19276 440
rect 19316 400 19317 440
rect 19275 391 19317 400
rect 20044 356 20084 820
rect 19852 316 20084 356
rect 19660 113 19700 198
rect 16780 55 16820 64
rect 19659 104 19701 113
rect 19659 64 19660 104
rect 19700 64 19701 104
rect 19659 55 19701 64
rect 19852 104 19892 316
rect 19852 55 19892 64
rect 20140 104 20180 2836
rect 23403 2876 23445 2885
rect 23403 2836 23404 2876
rect 23444 2836 23445 2876
rect 23403 2827 23445 2836
rect 20427 2792 20469 2801
rect 20427 2752 20428 2792
rect 20468 2752 20469 2792
rect 20427 2743 20469 2752
rect 20428 2624 20468 2743
rect 21868 2633 21908 2718
rect 20428 2372 20468 2584
rect 21867 2624 21909 2633
rect 21867 2584 21868 2624
rect 21908 2584 21909 2624
rect 21867 2575 21909 2584
rect 23404 2624 23444 2827
rect 24844 2717 24884 2911
rect 26571 2792 26613 2801
rect 26571 2752 26572 2792
rect 26612 2752 26613 2792
rect 26571 2743 26613 2752
rect 24843 2708 24885 2717
rect 24843 2668 24844 2708
rect 24884 2668 24885 2708
rect 24843 2659 24885 2668
rect 23404 2549 23444 2584
rect 23403 2540 23445 2549
rect 23403 2500 23404 2540
rect 23444 2500 23445 2540
rect 23403 2491 23445 2500
rect 20428 2323 20468 2332
rect 24844 1952 24884 2659
rect 26572 2624 26612 2743
rect 28108 2633 28148 2718
rect 30891 2708 30933 2717
rect 30891 2668 30892 2708
rect 30932 2668 30933 2708
rect 30891 2659 30933 2668
rect 26572 2575 26612 2584
rect 28107 2624 28149 2633
rect 28107 2584 28108 2624
rect 28148 2584 28149 2624
rect 28107 2575 28149 2584
rect 29548 2624 29588 2635
rect 29548 2465 29588 2584
rect 30892 2624 30932 2659
rect 30892 2573 30932 2584
rect 31660 2624 31700 3499
rect 31660 2575 31700 2584
rect 31756 3212 31796 3221
rect 29547 2456 29589 2465
rect 29547 2416 29548 2456
rect 29588 2416 29589 2456
rect 29547 2407 29589 2416
rect 24844 1903 24884 1912
rect 20428 1532 20468 1541
rect 20236 1196 20276 1205
rect 20236 776 20276 1156
rect 20236 727 20276 736
rect 20428 524 20468 1492
rect 23884 1532 23924 1541
rect 21004 1196 21044 1205
rect 20620 1028 20660 1037
rect 20620 869 20660 988
rect 20619 860 20661 869
rect 20619 820 20620 860
rect 20660 820 20661 860
rect 20619 811 20661 820
rect 20428 475 20468 484
rect 20620 281 20660 811
rect 21004 608 21044 1156
rect 22155 1196 22197 1205
rect 22155 1156 22156 1196
rect 22196 1156 22197 1196
rect 22155 1147 22197 1156
rect 22540 1196 22580 1205
rect 22156 1112 22196 1147
rect 22156 1061 22196 1072
rect 22540 617 22580 1156
rect 23308 1196 23348 1205
rect 22924 1028 22964 1037
rect 21004 356 21044 568
rect 22539 608 22581 617
rect 22539 568 22540 608
rect 22580 568 22581 608
rect 22539 559 22581 568
rect 22924 533 22964 988
rect 22923 524 22965 533
rect 22923 484 22924 524
rect 22964 484 22965 524
rect 22923 475 22965 484
rect 21004 307 21044 316
rect 20619 272 20661 281
rect 20619 232 20620 272
rect 20660 232 20661 272
rect 20619 223 20661 232
rect 22924 113 22964 475
rect 23308 188 23348 1156
rect 23788 1112 23828 1121
rect 23788 953 23828 1072
rect 23787 944 23829 953
rect 23787 904 23788 944
rect 23828 904 23829 944
rect 23787 895 23829 904
rect 23788 356 23828 895
rect 23884 524 23924 1492
rect 30700 1364 30740 1373
rect 24843 1280 24885 1289
rect 24843 1240 24844 1280
rect 24884 1240 24885 1280
rect 24843 1231 24885 1240
rect 26188 1280 26228 1289
rect 24460 1196 24500 1205
rect 24460 1121 24500 1156
rect 24459 1112 24501 1121
rect 24459 1072 24460 1112
rect 24500 1072 24501 1112
rect 24459 1063 24501 1072
rect 24844 1112 24884 1231
rect 24844 1063 24884 1072
rect 25515 1112 25557 1121
rect 25515 1072 25516 1112
rect 25556 1072 25557 1112
rect 25515 1063 25557 1072
rect 24460 953 24500 1063
rect 25516 978 25556 1063
rect 25899 1028 25941 1037
rect 25899 988 25900 1028
rect 25940 988 25941 1028
rect 25899 979 25941 988
rect 24459 944 24501 953
rect 24459 904 24460 944
rect 24500 904 24501 944
rect 24459 895 24501 904
rect 25900 894 25940 979
rect 26188 860 26228 1240
rect 26668 1196 26708 1205
rect 26668 869 26708 1156
rect 28203 1196 28245 1205
rect 28203 1156 28204 1196
rect 28244 1156 28245 1196
rect 28203 1147 28245 1156
rect 28204 1062 28244 1147
rect 29740 1112 29780 1121
rect 27628 1028 27668 1037
rect 26188 811 26228 820
rect 26667 860 26709 869
rect 26667 820 26668 860
rect 26708 820 26709 860
rect 26667 811 26709 820
rect 23884 475 23924 484
rect 26187 524 26229 533
rect 26187 484 26188 524
rect 26228 484 26229 524
rect 26187 475 26229 484
rect 27628 524 27668 988
rect 28587 608 28629 617
rect 28587 568 28588 608
rect 28628 568 28629 608
rect 28587 559 28629 568
rect 27628 475 27668 484
rect 27820 524 27860 533
rect 26188 390 26228 475
rect 23788 307 23828 316
rect 23308 139 23348 148
rect 20140 55 20180 64
rect 22923 104 22965 113
rect 22923 64 22924 104
rect 22964 64 22965 104
rect 22923 55 22965 64
rect 27820 104 27860 484
rect 28588 474 28628 559
rect 29740 533 29780 1072
rect 30124 1112 30164 1121
rect 29739 524 29781 533
rect 29739 484 29740 524
rect 29780 484 29781 524
rect 29739 475 29781 484
rect 29740 356 29780 475
rect 29740 307 29780 316
rect 30124 356 30164 1072
rect 30507 944 30549 953
rect 30507 904 30508 944
rect 30548 904 30549 944
rect 30507 895 30549 904
rect 30508 810 30548 895
rect 30700 608 30740 1324
rect 31083 1280 31125 1289
rect 31083 1240 31084 1280
rect 31124 1240 31125 1280
rect 31083 1231 31125 1240
rect 31084 1112 31124 1231
rect 31084 1063 31124 1072
rect 31467 1112 31509 1121
rect 31467 1072 31468 1112
rect 31508 1072 31509 1112
rect 31467 1063 31509 1072
rect 31468 978 31508 1063
rect 31756 944 31796 3172
rect 32236 2801 32276 3592
rect 35692 3473 35732 3760
rect 38092 3716 38132 3725
rect 35691 3464 35733 3473
rect 35691 3424 35692 3464
rect 35732 3424 35733 3464
rect 35691 3415 35733 3424
rect 36844 3464 36884 3473
rect 34348 3212 34388 3221
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 32235 2792 32277 2801
rect 32235 2752 32236 2792
rect 32276 2752 32277 2792
rect 32235 2743 32277 2752
rect 32236 2204 32276 2743
rect 33771 2624 33813 2633
rect 33771 2584 33772 2624
rect 33812 2584 33813 2624
rect 33771 2575 33813 2584
rect 33772 2490 33812 2575
rect 32236 2155 32276 2164
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 33004 1448 33044 1457
rect 32620 1280 32660 1289
rect 31852 1196 31892 1205
rect 31852 1037 31892 1156
rect 32236 1196 32276 1205
rect 31851 1028 31893 1037
rect 31851 988 31852 1028
rect 31892 988 31893 1028
rect 31851 979 31893 988
rect 31756 895 31796 904
rect 32236 776 32276 1156
rect 32620 869 32660 1240
rect 32619 860 32661 869
rect 32619 820 32620 860
rect 32660 820 32661 860
rect 32619 811 32661 820
rect 32236 727 32276 736
rect 32620 617 32660 811
rect 30700 559 30740 568
rect 32619 608 32661 617
rect 32619 568 32620 608
rect 32660 568 32661 608
rect 32619 559 32661 568
rect 33004 608 33044 1408
rect 34155 1196 34197 1205
rect 34155 1156 34156 1196
rect 34196 1156 34197 1196
rect 34155 1147 34197 1156
rect 34156 1062 34196 1147
rect 34060 1028 34100 1037
rect 34060 944 34100 988
rect 34252 1028 34292 1037
rect 34252 944 34292 988
rect 34060 904 34292 944
rect 33004 559 33044 568
rect 34348 449 34388 3172
rect 35308 3044 35348 3055
rect 35308 2969 35348 3004
rect 35307 2960 35349 2969
rect 35307 2920 35308 2960
rect 35348 2920 35349 2960
rect 35307 2911 35349 2920
rect 35308 2549 35348 2911
rect 35307 2540 35349 2549
rect 35307 2500 35308 2540
rect 35348 2500 35349 2540
rect 35307 2491 35349 2500
rect 35692 2465 35732 3415
rect 36844 2717 36884 3424
rect 38092 3212 38132 3676
rect 38092 3163 38132 3172
rect 38763 2876 38805 2885
rect 38763 2836 38764 2876
rect 38804 2836 38805 2876
rect 38763 2827 38805 2836
rect 36843 2708 36885 2717
rect 36843 2668 36844 2708
rect 36884 2668 36885 2708
rect 36843 2659 36885 2668
rect 38764 2624 38804 2827
rect 38764 2575 38804 2584
rect 35691 2456 35733 2465
rect 35691 2416 35692 2456
rect 35732 2416 35733 2456
rect 35691 2407 35733 2416
rect 35308 2372 35348 2381
rect 35596 2372 35636 2381
rect 35348 2332 35596 2372
rect 35308 2323 35348 2332
rect 35596 2323 35636 2332
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 37324 1868 37364 1877
rect 35116 1448 35156 1457
rect 35308 1448 35348 1457
rect 35156 1408 35252 1448
rect 35116 1399 35156 1408
rect 35116 1280 35156 1289
rect 34540 1112 34580 1121
rect 34444 1072 34540 1112
rect 34444 701 34484 1072
rect 34540 1063 34580 1072
rect 35020 1112 35060 1121
rect 35020 785 35060 1072
rect 35116 860 35156 1240
rect 35116 811 35156 820
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 35019 776 35061 785
rect 35019 736 35020 776
rect 35060 736 35061 776
rect 35019 727 35061 736
rect 35212 776 35252 1408
rect 35212 727 35252 736
rect 34443 692 34485 701
rect 34443 652 34444 692
rect 34484 652 34485 692
rect 34443 643 34485 652
rect 34347 440 34389 449
rect 34347 400 34348 440
rect 34388 400 34389 440
rect 34347 391 34389 400
rect 35019 440 35061 449
rect 35019 400 35020 440
rect 35060 400 35061 440
rect 35019 391 35061 400
rect 35308 440 35348 1408
rect 37035 1280 37077 1289
rect 37035 1240 37036 1280
rect 37076 1240 37077 1280
rect 37035 1231 37077 1240
rect 35404 1112 35444 1121
rect 35404 608 35444 1072
rect 37036 1112 37076 1231
rect 37036 1063 37076 1072
rect 37324 1112 37364 1828
rect 37324 953 37364 1072
rect 38476 1196 38516 1205
rect 36459 944 36501 953
rect 36459 904 36460 944
rect 36500 904 36501 944
rect 36459 895 36501 904
rect 37323 944 37365 953
rect 37323 904 37324 944
rect 37364 904 37365 944
rect 37323 895 37365 904
rect 36076 860 36116 871
rect 36076 785 36116 820
rect 36460 860 36500 895
rect 36460 809 36500 820
rect 36075 776 36117 785
rect 36075 736 36076 776
rect 36116 736 36117 776
rect 36075 727 36117 736
rect 35404 559 35444 568
rect 36076 533 36116 727
rect 38476 692 38516 1156
rect 38476 643 38516 652
rect 38860 1196 38900 1205
rect 38860 617 38900 1156
rect 39244 1196 39284 3928
rect 41355 3548 41397 3557
rect 41355 3508 41356 3548
rect 41396 3508 41397 3548
rect 41355 3499 41397 3508
rect 41356 3414 41396 3499
rect 41932 3128 41972 3137
rect 42220 3128 42260 5188
rect 46060 5144 46100 5153
rect 46060 4136 46100 5104
rect 55372 5144 55412 5153
rect 50380 4976 50420 4985
rect 46060 4087 46100 4096
rect 48364 4808 48404 4817
rect 41972 3088 42260 3128
rect 41932 3079 41972 3088
rect 40203 3044 40245 3053
rect 40203 3004 40204 3044
rect 40244 3004 40245 3044
rect 40203 2995 40245 3004
rect 42220 3044 42260 3088
rect 44620 3800 44660 3809
rect 44620 3053 44660 3760
rect 46060 3800 46100 3809
rect 42220 2995 42260 3004
rect 44619 3044 44661 3053
rect 44619 3004 44620 3044
rect 44660 3004 44661 3044
rect 44619 2995 44661 3004
rect 40204 2633 40244 2995
rect 40587 2960 40629 2969
rect 40587 2920 40588 2960
rect 40628 2920 40629 2960
rect 40587 2911 40629 2920
rect 40203 2624 40245 2633
rect 40203 2584 40204 2624
rect 40244 2584 40245 2624
rect 40203 2575 40245 2584
rect 40588 2465 40628 2911
rect 44043 2876 44085 2885
rect 44043 2836 44044 2876
rect 44084 2836 44085 2876
rect 44043 2827 44085 2836
rect 45004 2876 45044 2885
rect 41643 2792 41685 2801
rect 41643 2752 41644 2792
rect 41684 2752 41685 2792
rect 41643 2743 41685 2752
rect 42219 2792 42261 2801
rect 42219 2752 42220 2792
rect 42260 2752 42261 2792
rect 42219 2743 42261 2752
rect 41644 2633 41684 2743
rect 41836 2633 41876 2718
rect 42220 2633 42260 2743
rect 44044 2742 44084 2827
rect 42987 2708 43029 2717
rect 42987 2668 42988 2708
rect 43028 2668 43029 2708
rect 42987 2659 43029 2668
rect 41643 2624 41685 2633
rect 41643 2584 41644 2624
rect 41684 2584 41685 2624
rect 41643 2575 41685 2584
rect 41835 2624 41877 2633
rect 41835 2584 41836 2624
rect 41876 2584 41877 2624
rect 41835 2575 41877 2584
rect 42219 2624 42261 2633
rect 42219 2584 42220 2624
rect 42260 2584 42261 2624
rect 42219 2575 42261 2584
rect 42988 2624 43028 2659
rect 42988 2573 43028 2584
rect 41932 2540 41972 2549
rect 40587 2456 40629 2465
rect 40587 2416 40588 2456
rect 40628 2416 40629 2456
rect 40587 2407 40629 2416
rect 38859 608 38901 617
rect 38859 568 38860 608
rect 38900 568 38901 608
rect 38859 559 38901 568
rect 36075 524 36117 533
rect 36075 484 36076 524
rect 36116 484 36117 524
rect 36075 475 36117 484
rect 35308 391 35348 400
rect 30124 307 30164 316
rect 35020 306 35060 391
rect 39244 272 39284 1156
rect 39628 1280 39668 1289
rect 39628 1028 39668 1240
rect 40300 1205 40340 1224
rect 39628 979 39668 988
rect 40012 1196 40052 1205
rect 40012 776 40052 1156
rect 40299 1196 40341 1205
rect 40396 1196 40436 1205
rect 40299 1156 40300 1196
rect 40340 1156 40396 1196
rect 40299 1147 40341 1156
rect 40012 727 40052 736
rect 40396 701 40436 1156
rect 40779 1112 40821 1121
rect 40779 1072 40780 1112
rect 40820 1072 40821 1112
rect 40779 1063 40821 1072
rect 41548 1112 41588 1121
rect 40780 978 40820 1063
rect 40395 692 40437 701
rect 40395 652 40396 692
rect 40436 652 40437 692
rect 40395 643 40437 652
rect 41548 524 41588 1072
rect 41932 608 41972 2500
rect 42316 2540 42356 2549
rect 42316 1616 42356 2500
rect 45004 1877 45044 2836
rect 45003 1868 45045 1877
rect 45003 1828 45004 1868
rect 45044 1828 45045 1868
rect 45003 1819 45045 1828
rect 46060 1709 46100 3760
rect 47596 3716 47636 3725
rect 47596 3557 47636 3676
rect 47595 3548 47637 3557
rect 47595 3508 47596 3548
rect 47636 3508 47637 3548
rect 47595 3499 47637 3508
rect 47884 3548 47924 3557
rect 46156 3044 46196 3053
rect 46156 2129 46196 3004
rect 46539 3044 46581 3053
rect 46539 3004 46540 3044
rect 46580 3004 46581 3044
rect 46539 2995 46581 3004
rect 46540 2801 46580 2995
rect 46635 2876 46677 2885
rect 46635 2836 46636 2876
rect 46676 2836 46677 2876
rect 46635 2827 46677 2836
rect 46539 2792 46581 2801
rect 46539 2752 46540 2792
rect 46580 2752 46581 2792
rect 46539 2743 46581 2752
rect 46540 2624 46580 2743
rect 46540 2575 46580 2584
rect 46636 2549 46676 2827
rect 46635 2540 46677 2549
rect 46635 2500 46636 2540
rect 46676 2500 46677 2540
rect 46635 2491 46677 2500
rect 46155 2120 46197 2129
rect 46155 2080 46156 2120
rect 46196 2080 46197 2120
rect 46155 2071 46197 2080
rect 47884 2045 47924 3508
rect 48364 2885 48404 4768
rect 48940 4808 48980 4817
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 48940 4052 48980 4768
rect 48940 4003 48980 4012
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 50380 3464 50420 4936
rect 50380 3415 50420 3424
rect 52108 4388 52148 4397
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 48075 2876 48117 2885
rect 48075 2836 48076 2876
rect 48116 2836 48117 2876
rect 48075 2827 48117 2836
rect 48363 2876 48405 2885
rect 48363 2836 48364 2876
rect 48404 2836 48405 2876
rect 48363 2827 48405 2836
rect 48076 2708 48116 2827
rect 48076 2659 48116 2668
rect 48460 2633 48500 2718
rect 49323 2708 49365 2717
rect 49323 2668 49324 2708
rect 49364 2668 49365 2708
rect 49323 2659 49365 2668
rect 48459 2624 48501 2633
rect 48459 2584 48460 2624
rect 48500 2584 48501 2624
rect 48459 2575 48501 2584
rect 49324 2624 49364 2659
rect 49324 2573 49364 2584
rect 48364 2540 48404 2549
rect 47883 2036 47925 2045
rect 47883 1996 47884 2036
rect 47924 1996 47925 2036
rect 47883 1987 47925 1996
rect 45387 1700 45429 1709
rect 45387 1660 45388 1700
rect 45428 1660 45429 1700
rect 45387 1651 45429 1660
rect 46059 1700 46101 1709
rect 46059 1660 46060 1700
rect 46100 1660 46101 1700
rect 46059 1651 46101 1660
rect 42028 1028 42068 1037
rect 42028 785 42068 988
rect 42027 776 42069 785
rect 42027 736 42028 776
rect 42068 736 42069 776
rect 42027 727 42069 736
rect 42316 617 42356 1576
rect 44332 1448 44372 1457
rect 43275 1280 43317 1289
rect 43275 1240 43276 1280
rect 43316 1240 43317 1280
rect 43275 1231 43317 1240
rect 42700 1196 42740 1205
rect 42412 1112 42452 1121
rect 41932 559 41972 568
rect 42315 608 42357 617
rect 42315 568 42316 608
rect 42356 568 42357 608
rect 42315 559 42357 568
rect 41548 475 41588 484
rect 42412 356 42452 1072
rect 42700 1037 42740 1156
rect 43276 1112 43316 1231
rect 43276 1063 43316 1072
rect 43564 1112 43604 1121
rect 42699 1028 42741 1037
rect 42699 988 42700 1028
rect 42740 988 42741 1028
rect 42699 979 42741 988
rect 42700 869 42740 979
rect 43564 953 43604 1072
rect 43563 944 43605 953
rect 43563 904 43564 944
rect 43604 904 43605 944
rect 43563 895 43605 904
rect 42699 860 42741 869
rect 42699 820 42700 860
rect 42740 820 42741 860
rect 42699 811 42741 820
rect 44332 776 44372 1408
rect 44332 727 44372 736
rect 44428 1196 44468 1205
rect 43852 692 43892 701
rect 43852 440 43892 652
rect 43947 608 43989 617
rect 43947 568 43948 608
rect 43988 568 43989 608
rect 43947 559 43989 568
rect 43948 474 43988 559
rect 43852 391 43892 400
rect 44428 365 44468 1156
rect 45388 953 45428 1651
rect 48364 1373 48404 2500
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 50379 1952 50421 1961
rect 50379 1912 50380 1952
rect 50420 1912 50421 1952
rect 50379 1903 50421 1912
rect 51436 1952 51476 1961
rect 50380 1818 50420 1903
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 47979 1364 48021 1373
rect 47884 1324 47980 1364
rect 48020 1324 48021 1364
rect 47884 1280 47924 1324
rect 47979 1315 48021 1324
rect 48363 1364 48405 1373
rect 48363 1324 48364 1364
rect 48404 1324 48405 1364
rect 48363 1315 48405 1324
rect 51436 1364 51476 1912
rect 52108 1952 52148 4348
rect 52108 1903 52148 1912
rect 52492 4388 52532 4397
rect 47788 1240 47924 1280
rect 49228 1280 49268 1289
rect 46252 1196 46292 1205
rect 45387 944 45429 953
rect 45387 904 45388 944
rect 45428 904 45429 944
rect 45387 895 45429 904
rect 45484 944 45524 953
rect 45100 776 45140 785
rect 45100 533 45140 736
rect 45099 524 45141 533
rect 45099 484 45100 524
rect 45140 484 45141 524
rect 45099 475 45141 484
rect 42412 307 42452 316
rect 44427 356 44469 365
rect 44427 316 44428 356
rect 44468 316 44469 356
rect 44427 307 44469 316
rect 39244 223 39284 232
rect 45484 272 45524 904
rect 46252 440 46292 1156
rect 47788 1196 47828 1240
rect 47788 1147 47828 1156
rect 48075 1196 48117 1205
rect 48075 1156 48076 1196
rect 48116 1156 48117 1196
rect 48075 1147 48117 1156
rect 47019 1112 47061 1121
rect 47019 1072 47020 1112
rect 47060 1072 47061 1112
rect 47019 1063 47061 1072
rect 47692 1112 47732 1121
rect 46636 1028 46676 1037
rect 46636 701 46676 988
rect 47020 978 47060 1063
rect 46635 692 46677 701
rect 46635 652 46636 692
rect 46676 652 46677 692
rect 46635 643 46677 652
rect 46252 391 46292 400
rect 47692 356 47732 1072
rect 48076 785 48116 1147
rect 48940 1112 48980 1123
rect 48940 1037 48980 1072
rect 49131 1112 49173 1121
rect 49131 1072 49132 1112
rect 49172 1072 49173 1112
rect 49131 1063 49173 1072
rect 48939 1028 48981 1037
rect 48939 988 48940 1028
rect 48980 988 48981 1028
rect 48939 979 48981 988
rect 49132 978 49172 1063
rect 48075 776 48117 785
rect 48075 736 48076 776
rect 48116 736 48117 776
rect 48075 727 48117 736
rect 49228 608 49268 1240
rect 49515 1280 49557 1289
rect 49515 1240 49516 1280
rect 49556 1240 49557 1280
rect 49515 1231 49557 1240
rect 49516 953 49556 1231
rect 49707 1196 49749 1205
rect 49707 1156 49708 1196
rect 49748 1156 49749 1196
rect 49707 1147 49749 1156
rect 49708 1062 49748 1147
rect 51436 1112 51476 1324
rect 51436 1063 51476 1072
rect 50187 1028 50229 1037
rect 50187 988 50188 1028
rect 50228 988 50229 1028
rect 50187 979 50229 988
rect 49515 944 49557 953
rect 49515 904 49516 944
rect 49556 904 49557 944
rect 49515 895 49557 904
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 49228 559 49268 568
rect 49996 608 50036 617
rect 47692 307 47732 316
rect 49996 356 50036 568
rect 50188 533 50228 979
rect 52492 776 52532 4348
rect 55372 3716 55412 5104
rect 62380 4724 62420 4733
rect 58636 4136 58676 4145
rect 55372 3389 55412 3676
rect 58444 3800 58484 3809
rect 54316 3380 54356 3389
rect 54316 2633 54356 3340
rect 55371 3380 55413 3389
rect 55371 3340 55372 3380
rect 55412 3340 55413 3380
rect 55371 3331 55413 3340
rect 55084 3212 55124 3221
rect 54988 2960 55028 2969
rect 54507 2876 54549 2885
rect 54507 2836 54508 2876
rect 54548 2836 54549 2876
rect 54507 2827 54549 2836
rect 54508 2633 54548 2827
rect 54892 2792 54932 2801
rect 54315 2624 54357 2633
rect 54315 2584 54316 2624
rect 54356 2584 54357 2624
rect 54315 2575 54357 2584
rect 54507 2624 54549 2633
rect 54507 2584 54508 2624
rect 54548 2584 54549 2624
rect 54507 2575 54549 2584
rect 54892 2624 54932 2752
rect 54892 2575 54932 2584
rect 54316 2465 54356 2575
rect 54315 2456 54357 2465
rect 54315 2416 54316 2456
rect 54356 2416 54357 2456
rect 54315 2407 54357 2416
rect 54795 1700 54837 1709
rect 54795 1660 54796 1700
rect 54836 1660 54837 1700
rect 54795 1651 54837 1660
rect 54796 1289 54836 1651
rect 54795 1280 54837 1289
rect 54795 1240 54796 1280
rect 54836 1240 54837 1280
rect 54795 1231 54837 1240
rect 54988 860 55028 2920
rect 55084 1616 55124 3172
rect 55468 2456 55508 2465
rect 55508 2416 55604 2456
rect 55468 2407 55508 2416
rect 55564 2288 55604 2416
rect 55564 2239 55604 2248
rect 58444 2036 58484 3760
rect 58636 2624 58676 4096
rect 62380 4061 62420 4684
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 66796 4388 66836 4397
rect 66796 4145 66836 4348
rect 68523 4220 68565 4229
rect 68523 4180 68524 4220
rect 68564 4180 68565 4220
rect 68523 4171 68565 4180
rect 66508 4136 66548 4145
rect 62379 4052 62421 4061
rect 62379 4012 62380 4052
rect 62420 4012 62421 4052
rect 62379 4003 62421 4012
rect 66508 3977 66548 4096
rect 66795 4136 66837 4145
rect 66795 4096 66796 4136
rect 66836 4096 66837 4136
rect 66795 4087 66837 4096
rect 68524 4086 68564 4171
rect 66507 3968 66549 3977
rect 66507 3928 66508 3968
rect 66548 3928 66549 3968
rect 66507 3919 66549 3928
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 66219 3632 66261 3641
rect 66219 3592 66220 3632
rect 66260 3592 66261 3632
rect 66219 3583 66261 3592
rect 72459 3632 72501 3641
rect 72459 3592 72460 3632
rect 72500 3592 72501 3632
rect 72459 3583 72501 3592
rect 72939 3632 72981 3641
rect 72939 3592 72940 3632
rect 72980 3592 72981 3632
rect 72939 3583 72981 3592
rect 79179 3632 79221 3641
rect 79179 3592 79180 3632
rect 79220 3592 79221 3632
rect 79179 3583 79221 3592
rect 85323 3632 85365 3641
rect 85323 3592 85324 3632
rect 85364 3592 85365 3632
rect 85323 3583 85365 3592
rect 90700 3632 90740 3641
rect 64587 3464 64629 3473
rect 64587 3424 64588 3464
rect 64628 3424 64629 3464
rect 64587 3415 64629 3424
rect 65836 3464 65876 3473
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 64588 2801 64628 3415
rect 64684 3380 64724 3389
rect 64587 2792 64629 2801
rect 64587 2752 64588 2792
rect 64628 2752 64629 2792
rect 64587 2743 64629 2752
rect 64684 2792 64724 3340
rect 61323 2708 61365 2717
rect 61323 2668 61324 2708
rect 61364 2668 61365 2708
rect 61323 2659 61365 2668
rect 58636 2575 58676 2584
rect 61324 2574 61364 2659
rect 61708 2624 61748 2633
rect 58444 1987 58484 1996
rect 59116 2456 59156 2465
rect 55084 1567 55124 1576
rect 55468 1700 55508 1709
rect 55468 1532 55508 1660
rect 55468 1483 55508 1492
rect 55948 1700 55988 1709
rect 55948 1112 55988 1660
rect 59116 1121 59156 2416
rect 55948 1063 55988 1072
rect 59115 1112 59157 1121
rect 59115 1072 59116 1112
rect 59156 1072 59157 1112
rect 59115 1063 59157 1072
rect 54988 811 55028 820
rect 52492 727 52532 736
rect 59116 701 59156 1063
rect 61708 953 61748 2584
rect 63532 2624 63572 2633
rect 62571 1952 62613 1961
rect 62571 1912 62572 1952
rect 62612 1912 62613 1952
rect 62571 1903 62613 1912
rect 62572 1818 62612 1903
rect 63532 1877 63572 2584
rect 64012 2624 64052 2633
rect 64203 2624 64245 2633
rect 64052 2584 64204 2624
rect 64244 2584 64245 2624
rect 64012 2575 64052 2584
rect 64203 2575 64245 2584
rect 64299 2540 64341 2549
rect 64299 2500 64300 2540
rect 64340 2500 64341 2540
rect 64299 2491 64341 2500
rect 64300 2456 64340 2491
rect 64300 2405 64340 2416
rect 64588 1952 64628 2743
rect 64684 2129 64724 2752
rect 65356 3212 65396 3221
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 64683 2120 64725 2129
rect 64683 2080 64684 2120
rect 64724 2080 64725 2120
rect 64683 2071 64725 2080
rect 64588 1903 64628 1912
rect 63531 1868 63573 1877
rect 63531 1828 63532 1868
rect 63572 1828 63573 1868
rect 63531 1819 63573 1828
rect 64012 1700 64052 1709
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 62860 1364 62900 1373
rect 62667 1280 62709 1289
rect 62667 1240 62668 1280
rect 62708 1240 62709 1280
rect 62667 1231 62709 1240
rect 62668 1112 62708 1231
rect 61707 944 61749 953
rect 61707 904 61708 944
rect 61748 904 61749 944
rect 61707 895 61749 904
rect 59115 692 59157 701
rect 59115 652 59116 692
rect 59156 652 59157 692
rect 59115 643 59157 652
rect 62668 692 62708 1072
rect 62668 643 62708 652
rect 62764 1196 62804 1205
rect 62764 617 62804 1156
rect 62763 608 62805 617
rect 62763 568 62764 608
rect 62804 568 62805 608
rect 62763 559 62805 568
rect 50187 524 50229 533
rect 50187 484 50188 524
rect 50228 484 50229 524
rect 50187 475 50229 484
rect 62860 524 62900 1324
rect 63532 1196 63572 1207
rect 63532 1121 63572 1156
rect 62956 1112 62996 1121
rect 62956 944 62996 1072
rect 63051 1112 63093 1121
rect 63051 1072 63052 1112
rect 63092 1072 63093 1112
rect 63051 1063 63093 1072
rect 63531 1112 63573 1121
rect 63531 1072 63532 1112
rect 63572 1072 63573 1112
rect 63531 1063 63573 1072
rect 62956 895 62996 904
rect 62860 475 62900 484
rect 63052 449 63092 1063
rect 64012 944 64052 1660
rect 64012 895 64052 904
rect 64204 1364 64244 1373
rect 63051 440 63093 449
rect 63051 400 63052 440
rect 63092 400 63093 440
rect 63051 391 63093 400
rect 49996 307 50036 316
rect 45484 223 45524 232
rect 27820 55 27860 64
rect 64204 104 64244 1324
rect 64684 1364 64724 1373
rect 64300 1112 64340 1123
rect 64300 1037 64340 1072
rect 64588 1112 64628 1121
rect 64299 1028 64341 1037
rect 64299 988 64300 1028
rect 64340 988 64341 1028
rect 64299 979 64341 988
rect 64588 272 64628 1072
rect 64684 524 64724 1324
rect 65260 1364 65300 1373
rect 65260 860 65300 1324
rect 65356 944 65396 3172
rect 65836 2960 65876 3424
rect 66220 3464 66260 3583
rect 66220 3389 66260 3424
rect 69196 3548 69236 3557
rect 66219 3380 66261 3389
rect 66219 3340 66220 3380
rect 66260 3340 66261 3380
rect 66219 3331 66261 3340
rect 66603 3380 66645 3389
rect 66603 3340 66604 3380
rect 66644 3340 66645 3380
rect 66603 3331 66645 3340
rect 65836 2045 65876 2920
rect 66604 2456 66644 3331
rect 66988 3296 67028 3305
rect 66988 2465 67028 3256
rect 69196 2801 69236 3508
rect 69772 3548 69812 3557
rect 69195 2792 69237 2801
rect 69195 2752 69196 2792
rect 69236 2752 69237 2792
rect 69195 2743 69237 2752
rect 67851 2708 67893 2717
rect 67851 2668 67852 2708
rect 67892 2668 67893 2708
rect 67851 2659 67893 2668
rect 66604 2407 66644 2416
rect 66987 2456 67029 2465
rect 66987 2416 66988 2456
rect 67028 2416 67029 2456
rect 66987 2407 67029 2416
rect 65835 2036 65877 2045
rect 65835 1996 65836 2036
rect 65876 1996 65877 2036
rect 65835 1987 65877 1996
rect 67852 1952 67892 2659
rect 69196 2036 69236 2743
rect 69772 2633 69812 3508
rect 71308 3548 71348 3557
rect 71308 3473 71348 3508
rect 71307 3464 71349 3473
rect 71307 3424 71308 3464
rect 71348 3424 71349 3464
rect 71307 3415 71349 3424
rect 69771 2624 69813 2633
rect 69771 2584 69772 2624
rect 69812 2584 69813 2624
rect 69771 2575 69813 2584
rect 71308 2549 71348 3415
rect 72460 3380 72500 3583
rect 72844 3464 72884 3475
rect 72844 3389 72884 3424
rect 72460 3331 72500 3340
rect 72843 3380 72885 3389
rect 72843 3340 72844 3380
rect 72884 3340 72885 3380
rect 72843 3331 72885 3340
rect 72940 3212 72980 3583
rect 79180 3464 79220 3583
rect 79180 3415 79220 3424
rect 80332 3464 80372 3473
rect 78603 3380 78645 3389
rect 78603 3340 78604 3380
rect 78644 3340 78645 3380
rect 78603 3331 78645 3340
rect 72940 2708 72980 3172
rect 78604 2885 78644 3331
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 80332 2969 80372 3424
rect 84555 3464 84597 3473
rect 84555 3424 84556 3464
rect 84596 3424 84597 3464
rect 84555 3415 84597 3424
rect 83788 3212 83828 3221
rect 80331 2960 80373 2969
rect 80331 2920 80332 2960
rect 80372 2920 80373 2960
rect 80331 2911 80373 2920
rect 78603 2876 78645 2885
rect 78603 2836 78604 2876
rect 78644 2836 78645 2876
rect 78603 2827 78645 2836
rect 74763 2792 74805 2801
rect 74763 2752 74764 2792
rect 74804 2752 74805 2792
rect 74763 2743 74805 2752
rect 76875 2792 76917 2801
rect 76875 2752 76876 2792
rect 76916 2752 76917 2792
rect 76875 2743 76917 2752
rect 72940 2659 72980 2668
rect 74283 2708 74325 2717
rect 74283 2668 74284 2708
rect 74324 2668 74325 2708
rect 74283 2659 74325 2668
rect 71307 2540 71349 2549
rect 71307 2500 71308 2540
rect 71348 2500 71349 2540
rect 71307 2491 71349 2500
rect 74284 2540 74324 2659
rect 74764 2658 74804 2743
rect 75628 2633 75668 2718
rect 75627 2624 75669 2633
rect 75627 2584 75628 2624
rect 75668 2584 75669 2624
rect 75627 2575 75669 2584
rect 76876 2624 76916 2743
rect 76876 2549 76916 2584
rect 78604 2624 78644 2827
rect 80332 2717 80372 2911
rect 81771 2876 81813 2885
rect 81771 2836 81772 2876
rect 81812 2836 81908 2876
rect 81771 2827 81813 2836
rect 81868 2801 81908 2836
rect 81579 2792 81621 2801
rect 81579 2752 81580 2792
rect 81620 2752 81621 2792
rect 81868 2792 81921 2801
rect 81868 2752 81880 2792
rect 81920 2752 81921 2792
rect 81579 2743 81621 2752
rect 81879 2743 81921 2752
rect 80331 2708 80373 2717
rect 80331 2668 80332 2708
rect 80372 2668 80373 2708
rect 80331 2659 80373 2668
rect 81484 2633 81524 2718
rect 78604 2575 78644 2584
rect 81483 2624 81525 2633
rect 81483 2584 81484 2624
rect 81524 2584 81525 2624
rect 81483 2575 81525 2584
rect 81580 2549 81620 2743
rect 83403 2624 83445 2633
rect 83403 2584 83404 2624
rect 83444 2584 83445 2624
rect 83403 2575 83445 2584
rect 74284 2491 74324 2500
rect 76875 2540 76917 2549
rect 76875 2500 76876 2540
rect 76916 2500 76917 2540
rect 76875 2491 76917 2500
rect 77260 2540 77300 2549
rect 69196 1987 69236 1996
rect 67852 1903 67892 1912
rect 71308 1616 71348 1625
rect 70732 1532 70772 1541
rect 69388 1448 69428 1457
rect 65739 1364 65781 1373
rect 65739 1324 65740 1364
rect 65780 1324 65781 1364
rect 65739 1315 65781 1324
rect 66892 1364 66932 1373
rect 65356 895 65396 904
rect 65452 1112 65492 1121
rect 65260 811 65300 820
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 64684 475 64724 484
rect 65452 356 65492 1072
rect 65740 1112 65780 1315
rect 66603 1196 66645 1205
rect 66603 1156 66604 1196
rect 66644 1156 66645 1196
rect 66603 1147 66645 1156
rect 66795 1196 66837 1205
rect 66795 1156 66796 1196
rect 66836 1156 66837 1196
rect 66795 1147 66837 1156
rect 65740 785 65780 1072
rect 66604 869 66644 1147
rect 66796 1112 66836 1147
rect 66796 1061 66836 1072
rect 66892 944 66932 1324
rect 69388 1289 69428 1408
rect 69387 1280 69429 1289
rect 69387 1240 69388 1280
rect 69428 1240 69429 1280
rect 69387 1231 69429 1240
rect 66892 895 66932 904
rect 67276 1196 67316 1205
rect 67276 869 67316 1156
rect 68044 1196 68084 1205
rect 68044 869 68084 1156
rect 69772 1196 69812 1207
rect 69772 1121 69812 1156
rect 70156 1196 70196 1205
rect 68620 1112 68660 1121
rect 68620 953 68660 1072
rect 68812 1112 68852 1121
rect 68619 944 68661 953
rect 68619 904 68620 944
rect 68660 904 68661 944
rect 68619 895 68661 904
rect 66603 860 66645 869
rect 66603 820 66604 860
rect 66644 820 66645 860
rect 66603 811 66645 820
rect 67275 860 67317 869
rect 67275 820 67276 860
rect 67316 820 67317 860
rect 67275 811 67317 820
rect 68043 860 68085 869
rect 68043 820 68044 860
rect 68084 820 68085 860
rect 68043 811 68085 820
rect 65739 776 65781 785
rect 65739 736 65740 776
rect 65780 736 65781 776
rect 65739 727 65781 736
rect 66700 692 66740 703
rect 66700 617 66740 652
rect 66699 608 66741 617
rect 66699 568 66700 608
rect 66740 568 66741 608
rect 66699 559 66741 568
rect 65452 307 65492 316
rect 64588 223 64628 232
rect 64204 55 64244 64
rect 67276 104 67316 811
rect 68044 533 68084 811
rect 68812 617 68852 1072
rect 69771 1112 69813 1121
rect 69771 1072 69772 1112
rect 69812 1072 69813 1112
rect 69771 1063 69813 1072
rect 70156 860 70196 1156
rect 70444 1196 70484 1205
rect 70444 1037 70484 1156
rect 70443 1028 70485 1037
rect 70443 988 70444 1028
rect 70484 988 70485 1028
rect 70443 979 70485 988
rect 70156 811 70196 820
rect 70539 692 70581 701
rect 70539 652 70540 692
rect 70580 652 70581 692
rect 70539 643 70581 652
rect 68811 608 68853 617
rect 68811 568 68812 608
rect 68852 568 68853 608
rect 68811 559 68853 568
rect 70540 558 70580 643
rect 68043 524 68085 533
rect 68043 484 68044 524
rect 68084 484 68085 524
rect 68043 475 68085 484
rect 70732 188 70772 1492
rect 71308 1028 71348 1576
rect 73036 1448 73076 1457
rect 71308 979 71348 988
rect 71500 1364 71540 1373
rect 70924 944 70964 953
rect 70924 524 70964 904
rect 71500 860 71540 1324
rect 72268 1364 72308 1373
rect 71500 811 71540 820
rect 72076 1196 72116 1205
rect 72076 785 72116 1156
rect 72268 944 72308 1324
rect 72939 1364 72981 1373
rect 72939 1324 72940 1364
rect 72980 1324 72981 1364
rect 72939 1315 72981 1324
rect 72844 1280 72884 1289
rect 72459 1196 72501 1205
rect 72459 1156 72460 1196
rect 72500 1156 72501 1196
rect 72459 1147 72501 1156
rect 72651 1196 72693 1205
rect 72651 1156 72652 1196
rect 72692 1156 72693 1196
rect 72651 1147 72693 1156
rect 72460 1062 72500 1147
rect 72652 953 72692 1147
rect 72268 895 72308 904
rect 72651 944 72693 953
rect 72651 904 72652 944
rect 72692 904 72693 944
rect 72651 895 72693 904
rect 72075 776 72117 785
rect 72075 736 72076 776
rect 72116 736 72117 776
rect 72075 727 72117 736
rect 70924 475 70964 484
rect 72844 356 72884 1240
rect 72940 1196 72980 1315
rect 72940 1147 72980 1156
rect 72844 307 72884 316
rect 72940 776 72980 785
rect 70732 139 70772 148
rect 67276 55 67316 64
rect 72940 104 72980 736
rect 73036 692 73076 1408
rect 75531 1280 75573 1289
rect 75531 1240 75532 1280
rect 75572 1240 75573 1280
rect 74764 1205 74804 1236
rect 75531 1231 75573 1240
rect 73612 1196 73652 1205
rect 73612 776 73652 1156
rect 74763 1196 74805 1205
rect 74763 1156 74764 1196
rect 74804 1156 74805 1196
rect 74763 1147 74805 1156
rect 74764 1112 74804 1147
rect 75532 1146 75572 1231
rect 74764 1037 74804 1072
rect 75915 1112 75957 1121
rect 75915 1072 75916 1112
rect 75956 1072 75957 1112
rect 75915 1063 75957 1072
rect 76300 1112 76340 1121
rect 74763 1028 74805 1037
rect 74763 988 74764 1028
rect 74804 988 74805 1028
rect 74763 979 74805 988
rect 75916 978 75956 1063
rect 74859 944 74901 953
rect 74859 904 74860 944
rect 74900 904 74901 944
rect 74859 895 74901 904
rect 74379 860 74421 869
rect 74379 820 74380 860
rect 74420 820 74421 860
rect 74379 811 74421 820
rect 74860 860 74900 895
rect 73612 727 73652 736
rect 74380 726 74420 811
rect 74860 809 74900 820
rect 75148 860 75188 869
rect 73036 643 73076 652
rect 75148 617 75188 820
rect 76300 701 76340 1072
rect 76683 860 76725 869
rect 76683 820 76684 860
rect 76724 820 76725 860
rect 76683 811 76725 820
rect 76299 692 76341 701
rect 76299 652 76300 692
rect 76340 652 76341 692
rect 76299 643 76341 652
rect 75147 608 75189 617
rect 75147 568 75148 608
rect 75188 568 75189 608
rect 75147 559 75189 568
rect 76300 272 76340 643
rect 76684 449 76724 811
rect 77260 524 77300 2500
rect 81579 2540 81621 2549
rect 81579 2500 81580 2540
rect 81620 2500 81621 2540
rect 81579 2491 81621 2500
rect 83404 2490 83444 2575
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 79948 1868 79988 1877
rect 79852 1616 79892 1625
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 79756 1532 79796 1541
rect 79180 1280 79220 1289
rect 78603 1196 78645 1205
rect 78603 1156 78604 1196
rect 78644 1156 78645 1196
rect 78603 1147 78645 1156
rect 78604 1028 78644 1147
rect 78604 979 78644 988
rect 78220 944 78260 953
rect 78220 785 78260 904
rect 78219 776 78261 785
rect 78219 736 78220 776
rect 78260 736 78261 776
rect 78219 727 78261 736
rect 77260 475 77300 484
rect 79180 524 79220 1240
rect 79756 776 79796 1492
rect 79756 727 79796 736
rect 79852 608 79892 1576
rect 79948 1037 79988 1828
rect 81484 1448 81524 1457
rect 80524 1364 80564 1373
rect 79947 1028 79989 1037
rect 79947 988 79948 1028
rect 79988 988 79989 1028
rect 79947 979 79989 988
rect 80524 869 80564 1324
rect 81484 1289 81524 1408
rect 82828 1364 82868 1373
rect 81100 1280 81140 1289
rect 80811 1112 80853 1121
rect 80811 1072 80812 1112
rect 80852 1072 80853 1112
rect 80811 1063 80853 1072
rect 80812 953 80852 1063
rect 80811 944 80853 953
rect 80811 904 80812 944
rect 80852 904 80853 944
rect 80811 895 80853 904
rect 80523 860 80565 869
rect 80523 820 80524 860
rect 80564 820 80565 860
rect 80523 811 80565 820
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 79852 559 79892 568
rect 81100 533 81140 1240
rect 81483 1280 81525 1289
rect 81483 1240 81484 1280
rect 81524 1240 81525 1280
rect 81483 1231 81525 1240
rect 81868 1112 81908 1121
rect 81868 953 81908 1072
rect 82252 1112 82292 1121
rect 81867 944 81909 953
rect 81867 904 81868 944
rect 81908 904 81909 944
rect 81867 895 81909 904
rect 82252 944 82292 1072
rect 81868 701 81908 895
rect 81867 692 81909 701
rect 81867 652 81868 692
rect 81908 652 81909 692
rect 81867 643 81909 652
rect 79180 475 79220 484
rect 81099 524 81141 533
rect 81099 484 81100 524
rect 81140 484 81141 524
rect 81099 475 81141 484
rect 76683 440 76725 449
rect 76683 400 76684 440
rect 76724 400 76725 440
rect 76683 391 76725 400
rect 76300 223 76340 232
rect 82252 272 82292 904
rect 82636 1112 82676 1121
rect 82636 533 82676 1072
rect 82828 776 82868 1324
rect 82828 727 82868 736
rect 83020 1112 83060 1121
rect 83020 608 83060 1072
rect 83788 776 83828 3172
rect 84556 2456 84596 3415
rect 85324 2801 85364 3583
rect 90700 3473 90740 3592
rect 90699 3464 90741 3473
rect 90699 3424 90700 3464
rect 90740 3424 90741 3464
rect 90699 3415 90741 3424
rect 92812 3464 92852 3473
rect 86475 2876 86517 2885
rect 86475 2836 86476 2876
rect 86516 2836 86517 2876
rect 86475 2827 86517 2836
rect 84556 2407 84596 2416
rect 84748 2792 84788 2801
rect 84748 2456 84788 2752
rect 84939 2792 84981 2801
rect 84939 2752 84940 2792
rect 84980 2752 84981 2792
rect 84939 2743 84981 2752
rect 85323 2792 85365 2801
rect 85323 2752 85324 2792
rect 85364 2752 85365 2792
rect 85323 2743 85365 2752
rect 84940 2549 84980 2743
rect 85324 2708 85364 2743
rect 85324 2658 85364 2668
rect 86476 2624 86516 2827
rect 90700 2801 90740 3415
rect 91467 3380 91509 3389
rect 91467 3340 91468 3380
rect 91508 3340 91509 3380
rect 91467 3331 91509 3340
rect 91468 2885 91508 3331
rect 92812 2969 92852 3424
rect 97131 3380 97173 3389
rect 97131 3340 97132 3380
rect 97172 3340 97173 3380
rect 97131 3331 97173 3340
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 92811 2960 92853 2969
rect 92811 2920 92812 2960
rect 92852 2920 92853 2960
rect 92811 2911 92853 2920
rect 91467 2876 91509 2885
rect 91467 2836 91468 2876
rect 91508 2836 91509 2876
rect 91467 2827 91509 2836
rect 92812 2876 92852 2911
rect 90699 2792 90741 2801
rect 90699 2752 90700 2792
rect 90740 2752 90741 2792
rect 90699 2743 90741 2752
rect 91468 2742 91508 2827
rect 92812 2796 92852 2836
rect 96363 2792 96405 2801
rect 96363 2752 96364 2792
rect 96404 2752 96405 2792
rect 96363 2743 96405 2752
rect 88011 2708 88053 2717
rect 88011 2668 88012 2708
rect 88052 2668 88053 2708
rect 88011 2659 88053 2668
rect 93675 2708 93717 2717
rect 93675 2668 93676 2708
rect 93716 2668 93717 2708
rect 93675 2659 93717 2668
rect 93867 2708 93909 2717
rect 93867 2668 93868 2708
rect 93908 2668 93909 2708
rect 93867 2659 93909 2668
rect 86476 2575 86516 2584
rect 88012 2574 88052 2659
rect 89547 2624 89589 2633
rect 89547 2584 89548 2624
rect 89588 2584 89589 2624
rect 89547 2575 89589 2584
rect 84939 2540 84981 2549
rect 84939 2500 84940 2540
rect 84980 2500 84981 2540
rect 84939 2491 84981 2500
rect 85228 2540 85268 2549
rect 84748 2407 84788 2416
rect 83788 727 83828 736
rect 84172 1112 84212 1121
rect 84172 860 84212 1072
rect 84556 1112 84596 1123
rect 84556 1037 84596 1072
rect 84555 1028 84597 1037
rect 84555 988 84556 1028
rect 84596 988 84597 1028
rect 84555 979 84597 988
rect 83499 692 83541 701
rect 83499 652 83500 692
rect 83540 652 83541 692
rect 83499 643 83541 652
rect 82635 524 82677 533
rect 82635 484 82636 524
rect 82676 484 82677 524
rect 82635 475 82677 484
rect 82252 223 82292 232
rect 83020 188 83060 568
rect 83500 449 83540 643
rect 84172 617 84212 820
rect 85228 860 85268 2500
rect 89548 2490 89588 2575
rect 93676 2574 93716 2659
rect 91083 2540 91125 2549
rect 91083 2500 91084 2540
rect 91124 2500 91125 2540
rect 91083 2491 91125 2500
rect 91084 2406 91124 2491
rect 93868 2372 93908 2659
rect 95115 2624 95157 2633
rect 95115 2584 95116 2624
rect 95156 2584 95157 2624
rect 95115 2575 95157 2584
rect 96364 2624 96404 2743
rect 96364 2575 96404 2584
rect 96747 2624 96789 2633
rect 96747 2584 96748 2624
rect 96788 2584 96789 2624
rect 96747 2575 96789 2584
rect 97132 2624 97172 3331
rect 97132 2575 97172 2584
rect 95116 2490 95156 2575
rect 96748 2490 96788 2575
rect 97996 2540 98036 2549
rect 93868 2323 93908 2332
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 94828 1532 94868 1541
rect 88396 1448 88436 1457
rect 85228 811 85268 820
rect 85324 1364 85364 1373
rect 85324 692 85364 1324
rect 85708 1280 85748 1289
rect 84171 608 84213 617
rect 84171 568 84172 608
rect 84212 568 84213 608
rect 84171 559 84213 568
rect 83499 440 83541 449
rect 83499 400 83500 440
rect 83540 400 83541 440
rect 83499 391 83541 400
rect 85324 440 85364 652
rect 85612 1112 85652 1121
rect 85612 692 85652 1072
rect 85612 643 85652 652
rect 85324 391 85364 400
rect 83020 139 83060 148
rect 85708 188 85748 1240
rect 87627 1280 87669 1289
rect 87627 1240 87628 1280
rect 87668 1240 87669 1280
rect 87627 1231 87669 1240
rect 87819 1280 87861 1289
rect 87819 1240 87820 1280
rect 87860 1240 87861 1280
rect 87819 1231 87861 1240
rect 86859 1196 86901 1205
rect 86859 1156 86860 1196
rect 86900 1156 86901 1196
rect 86859 1147 86901 1156
rect 86956 1196 86996 1205
rect 86476 1112 86516 1121
rect 86476 869 86516 1072
rect 86860 1112 86900 1147
rect 86860 1061 86900 1072
rect 86475 860 86517 869
rect 86475 820 86476 860
rect 86516 820 86517 860
rect 86475 811 86517 820
rect 86956 701 86996 1156
rect 87628 1121 87668 1231
rect 87627 1112 87669 1121
rect 87627 1072 87628 1112
rect 87668 1072 87669 1112
rect 87627 1063 87669 1072
rect 87820 701 87860 1231
rect 88012 1196 88052 1205
rect 88012 701 88052 1156
rect 88396 944 88436 1408
rect 88396 895 88436 904
rect 88780 1364 88820 1373
rect 86955 692 86997 701
rect 86955 652 86956 692
rect 86996 652 86997 692
rect 86955 643 86997 652
rect 87819 692 87861 701
rect 87819 652 87820 692
rect 87860 652 87861 692
rect 87819 643 87861 652
rect 88011 692 88053 701
rect 88011 652 88012 692
rect 88052 652 88053 692
rect 88011 643 88053 652
rect 88012 449 88052 643
rect 88780 533 88820 1324
rect 89932 1280 89972 1289
rect 89164 1196 89204 1205
rect 89164 608 89204 1156
rect 89548 1196 89588 1205
rect 89548 1028 89588 1156
rect 89548 979 89588 988
rect 89932 860 89972 1240
rect 89932 811 89972 820
rect 90316 1280 90356 1289
rect 90316 617 90356 1240
rect 92620 1280 92660 1289
rect 91084 1112 91124 1121
rect 90699 1028 90741 1037
rect 90699 988 90700 1028
rect 90740 988 90741 1028
rect 90699 979 90741 988
rect 90700 894 90740 979
rect 91084 692 91124 1072
rect 91084 643 91124 652
rect 91468 1112 91508 1121
rect 89164 559 89204 568
rect 90315 608 90357 617
rect 90315 568 90316 608
rect 90356 568 90357 608
rect 90315 559 90357 568
rect 88779 524 88821 533
rect 88779 484 88780 524
rect 88820 484 88821 524
rect 88779 475 88821 484
rect 88011 440 88053 449
rect 88011 400 88012 440
rect 88052 400 88053 440
rect 88011 391 88053 400
rect 91468 440 91508 1072
rect 91468 391 91508 400
rect 91852 1112 91892 1121
rect 85708 139 85748 148
rect 91852 188 91892 1072
rect 92043 1028 92085 1037
rect 92043 988 92044 1028
rect 92084 988 92085 1028
rect 92043 979 92085 988
rect 92044 894 92084 979
rect 92620 869 92660 1240
rect 93195 1280 93237 1289
rect 93195 1240 93196 1280
rect 93236 1240 93237 1280
rect 93004 1205 93044 1236
rect 93195 1231 93237 1240
rect 94540 1280 94580 1289
rect 93003 1196 93045 1205
rect 93003 1156 93004 1196
rect 93044 1156 93045 1196
rect 93003 1147 93045 1156
rect 93004 1112 93044 1147
rect 93196 1146 93236 1231
rect 93004 953 93044 1072
rect 93579 1112 93621 1121
rect 93579 1072 93580 1112
rect 93620 1072 93621 1112
rect 93579 1063 93621 1072
rect 93964 1112 94004 1121
rect 93580 978 93620 1063
rect 93003 944 93045 953
rect 93003 904 93004 944
rect 93044 904 93045 944
rect 93003 895 93045 904
rect 92619 860 92661 869
rect 92619 820 92620 860
rect 92660 820 92661 860
rect 92619 811 92661 820
rect 92620 356 92660 811
rect 93964 701 94004 1072
rect 94540 860 94580 1240
rect 94540 811 94580 820
rect 94732 1112 94772 1121
rect 93963 692 94005 701
rect 93963 652 93964 692
rect 94004 652 94005 692
rect 93963 643 94005 652
rect 94732 533 94772 1072
rect 94828 776 94868 1492
rect 97228 1532 97268 1541
rect 94828 727 94868 736
rect 94924 1448 94964 1457
rect 94924 608 94964 1408
rect 96268 1112 96308 1121
rect 95500 860 95540 869
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
rect 94924 559 94964 568
rect 94731 524 94773 533
rect 94731 484 94732 524
rect 94772 484 94773 524
rect 94731 475 94773 484
rect 92620 307 92660 316
rect 91852 139 91892 148
rect 72940 55 72980 64
rect 95500 104 95540 820
rect 96268 617 96308 1072
rect 96651 1112 96693 1121
rect 96651 1072 96652 1112
rect 96692 1072 96693 1112
rect 96651 1063 96693 1072
rect 96652 978 96692 1063
rect 97228 776 97268 1492
rect 97996 944 98036 2500
rect 99148 1112 99188 1121
rect 99148 953 99188 1072
rect 97996 895 98036 904
rect 99147 944 99189 953
rect 99147 904 99148 944
rect 99188 904 99189 944
rect 99147 895 99189 904
rect 97228 727 97268 736
rect 96267 608 96309 617
rect 96267 568 96268 608
rect 96308 568 96309 608
rect 96267 559 96309 568
rect 95500 55 95540 64
<< via4 >>
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 26092 4096 26132 4136
rect 28012 4012 28052 4052
rect 38956 4180 38996 4220
rect 38668 3928 38708 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 11116 3676 11156 3716
rect 17164 3676 17204 3716
rect 9580 3508 9620 3548
rect 5932 3424 5972 3464
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 2284 2584 2324 2624
rect 3916 2584 3956 2624
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 1228 904 1268 944
rect 1996 1072 2036 1112
rect 2764 1072 2804 1112
rect 1612 568 1652 608
rect 6892 3172 6932 3212
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 4300 1072 4340 1112
rect 4684 904 4724 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 6508 820 6548 860
rect 8044 2668 8084 2708
rect 7180 2584 7220 2624
rect 15820 3508 15860 3548
rect 11500 3340 11540 3380
rect 13036 3172 13076 3212
rect 19372 3508 19412 3548
rect 25324 3508 25364 3548
rect 31660 3508 31700 3548
rect 17548 3340 17588 3380
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 19372 3172 19412 3212
rect 18700 2920 18740 2960
rect 17164 2836 17204 2876
rect 14284 2668 14324 2708
rect 15820 2668 15860 2708
rect 12748 2584 12788 2624
rect 18700 2584 18740 2624
rect 9580 2500 9620 2540
rect 23788 3340 23828 3380
rect 29836 3340 29876 3380
rect 24844 2920 24884 2960
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 7564 1324 7604 1364
rect 6892 1240 6932 1280
rect 6892 988 6932 1028
rect 10060 1240 10100 1280
rect 8332 1156 8372 1196
rect 9868 1072 9908 1112
rect 10060 1072 10100 1112
rect 8332 988 8372 1028
rect 10252 904 10292 944
rect 7564 736 7604 776
rect 7180 568 7220 608
rect 11404 1240 11444 1280
rect 12556 1240 12596 1280
rect 11212 904 11252 944
rect 11404 904 11444 944
rect 12940 1072 12980 1112
rect 12076 988 12116 1028
rect 12268 988 12308 1028
rect 13708 736 13748 776
rect 13324 400 13364 440
rect 16012 1156 16052 1196
rect 16492 904 16532 944
rect 16396 568 16436 608
rect 14380 232 14420 272
rect 18700 1240 18740 1280
rect 17548 1072 17588 1112
rect 18316 1072 18356 1112
rect 17548 904 17588 944
rect 19372 736 19412 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 19276 400 19316 440
rect 19660 64 19700 104
rect 23404 2836 23444 2876
rect 20428 2752 20468 2792
rect 21868 2584 21908 2624
rect 26572 2752 26612 2792
rect 24844 2668 24884 2708
rect 23404 2500 23444 2540
rect 30892 2668 30932 2708
rect 28108 2584 28148 2624
rect 29548 2416 29588 2456
rect 20620 820 20660 860
rect 22156 1156 22196 1196
rect 22540 568 22580 608
rect 22924 484 22964 524
rect 20620 232 20660 272
rect 23788 904 23828 944
rect 24844 1240 24884 1280
rect 24460 1072 24500 1112
rect 25516 1072 25556 1112
rect 25900 988 25940 1028
rect 24460 904 24500 944
rect 28204 1156 28244 1196
rect 26668 820 26708 860
rect 26188 484 26228 524
rect 28588 568 28628 608
rect 22924 64 22964 104
rect 29740 484 29780 524
rect 30508 904 30548 944
rect 31084 1240 31124 1280
rect 31468 1072 31508 1112
rect 35692 3424 35732 3464
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 32236 2752 32276 2792
rect 33772 2584 33812 2624
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 31852 988 31892 1028
rect 32620 820 32660 860
rect 32620 568 32660 608
rect 34156 1156 34196 1196
rect 35308 2920 35348 2960
rect 35308 2500 35348 2540
rect 38764 2836 38804 2876
rect 36844 2668 36884 2708
rect 35692 2416 35732 2456
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 35020 736 35060 776
rect 34444 652 34484 692
rect 34348 400 34388 440
rect 35020 400 35060 440
rect 37036 1240 37076 1280
rect 36460 904 36500 944
rect 37324 904 37364 944
rect 36076 736 36116 776
rect 41356 3508 41396 3548
rect 40204 3004 40244 3044
rect 44620 3004 44660 3044
rect 40588 2920 40628 2960
rect 40204 2584 40244 2624
rect 44044 2836 44084 2876
rect 41644 2752 41684 2792
rect 42220 2752 42260 2792
rect 42988 2668 43028 2708
rect 41644 2584 41684 2624
rect 41836 2584 41876 2624
rect 42220 2584 42260 2624
rect 40588 2416 40628 2456
rect 38860 568 38900 608
rect 36076 484 36116 524
rect 40300 1156 40340 1196
rect 40780 1072 40820 1112
rect 40396 652 40436 692
rect 45004 1828 45044 1868
rect 47596 3508 47636 3548
rect 46540 3004 46580 3044
rect 46636 2836 46676 2876
rect 46540 2752 46580 2792
rect 46636 2500 46676 2540
rect 46156 2080 46196 2120
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 48076 2836 48116 2876
rect 48364 2836 48404 2876
rect 49324 2668 49364 2708
rect 48460 2584 48500 2624
rect 47884 1996 47924 2036
rect 45388 1660 45428 1700
rect 46060 1660 46100 1700
rect 42028 736 42068 776
rect 43276 1240 43316 1280
rect 42316 568 42356 608
rect 42700 988 42740 1028
rect 43564 904 43604 944
rect 42700 820 42740 860
rect 43948 568 43988 608
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 50380 1912 50420 1952
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 47980 1324 48020 1364
rect 48364 1324 48404 1364
rect 45388 904 45428 944
rect 45100 484 45140 524
rect 44428 316 44468 356
rect 48076 1156 48116 1196
rect 47020 1072 47060 1112
rect 46636 652 46676 692
rect 49132 1072 49172 1112
rect 48940 988 48980 1028
rect 48076 736 48116 776
rect 49516 1240 49556 1280
rect 49708 1156 49748 1196
rect 50188 988 50228 1028
rect 49516 904 49556 944
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 55372 3340 55412 3380
rect 54508 2836 54548 2876
rect 54316 2584 54356 2624
rect 54508 2584 54548 2624
rect 54316 2416 54356 2456
rect 54796 1660 54836 1700
rect 54796 1240 54836 1280
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 68524 4180 68564 4220
rect 62380 4012 62420 4052
rect 66796 4096 66836 4136
rect 66508 3928 66548 3968
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 66220 3592 66260 3632
rect 72460 3592 72500 3632
rect 72940 3592 72980 3632
rect 79180 3592 79220 3632
rect 85324 3592 85364 3632
rect 64588 3424 64628 3464
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 64588 2752 64628 2792
rect 61324 2668 61364 2708
rect 59116 1072 59156 1112
rect 62572 1912 62612 1952
rect 64204 2584 64244 2624
rect 64300 2500 64340 2540
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 64684 2080 64724 2120
rect 63532 1828 63572 1868
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 62668 1240 62708 1280
rect 61708 904 61748 944
rect 59116 652 59156 692
rect 62764 568 62804 608
rect 50188 484 50228 524
rect 63052 1072 63092 1112
rect 63532 1072 63572 1112
rect 63052 400 63092 440
rect 64300 988 64340 1028
rect 66220 3340 66260 3380
rect 66604 3340 66644 3380
rect 69196 2752 69236 2792
rect 67852 2668 67892 2708
rect 66988 2416 67028 2456
rect 65836 1996 65876 2036
rect 71308 3424 71348 3464
rect 69772 2584 69812 2624
rect 72844 3340 72884 3380
rect 78604 3340 78644 3380
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 84556 3424 84596 3464
rect 80332 2920 80372 2960
rect 78604 2836 78644 2876
rect 74764 2752 74804 2792
rect 76876 2752 76916 2792
rect 74284 2668 74324 2708
rect 71308 2500 71348 2540
rect 75628 2584 75668 2624
rect 81772 2836 81812 2876
rect 81580 2752 81620 2792
rect 81880 2752 81920 2792
rect 80332 2668 80372 2708
rect 81484 2584 81524 2624
rect 83404 2584 83444 2624
rect 76876 2500 76916 2540
rect 65740 1324 65780 1364
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 66604 1156 66644 1196
rect 66796 1156 66836 1196
rect 69388 1240 69428 1280
rect 68620 904 68660 944
rect 66604 820 66644 860
rect 67276 820 67316 860
rect 68044 820 68084 860
rect 65740 736 65780 776
rect 66700 568 66740 608
rect 69772 1072 69812 1112
rect 70444 988 70484 1028
rect 70540 652 70580 692
rect 68812 568 68852 608
rect 68044 484 68084 524
rect 72940 1324 72980 1364
rect 72460 1156 72500 1196
rect 72652 1156 72692 1196
rect 72652 904 72692 944
rect 72076 736 72116 776
rect 75532 1240 75572 1280
rect 74764 1156 74804 1196
rect 75916 1072 75956 1112
rect 74764 988 74804 1028
rect 74860 904 74900 944
rect 74380 820 74420 860
rect 76684 820 76724 860
rect 76300 652 76340 692
rect 75148 568 75188 608
rect 81580 2500 81620 2540
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 78604 1156 78644 1196
rect 78220 736 78260 776
rect 79948 988 79988 1028
rect 80812 1072 80852 1112
rect 80812 904 80852 944
rect 80524 820 80564 860
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 81484 1240 81524 1280
rect 81868 904 81908 944
rect 81868 652 81908 692
rect 81100 484 81140 524
rect 76684 400 76724 440
rect 90700 3424 90740 3464
rect 86476 2836 86516 2876
rect 84940 2752 84980 2792
rect 85324 2752 85364 2792
rect 91468 3340 91508 3380
rect 97132 3340 97172 3380
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 92812 2920 92852 2960
rect 91468 2836 91508 2876
rect 90700 2752 90740 2792
rect 96364 2752 96404 2792
rect 88012 2668 88052 2708
rect 93676 2668 93716 2708
rect 93868 2668 93908 2708
rect 89548 2584 89588 2624
rect 84940 2500 84980 2540
rect 84556 988 84596 1028
rect 83500 652 83540 692
rect 82636 484 82676 524
rect 91084 2500 91124 2540
rect 95116 2584 95156 2624
rect 96748 2584 96788 2624
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 84172 568 84212 608
rect 83500 400 83540 440
rect 87628 1240 87668 1280
rect 87820 1240 87860 1280
rect 86860 1156 86900 1196
rect 86476 820 86516 860
rect 87628 1072 87668 1112
rect 86956 652 86996 692
rect 87820 652 87860 692
rect 88012 652 88052 692
rect 90700 988 90740 1028
rect 90316 568 90356 608
rect 88780 484 88820 524
rect 88012 400 88052 440
rect 92044 988 92084 1028
rect 93196 1240 93236 1280
rect 93004 1156 93044 1196
rect 93580 1072 93620 1112
rect 93004 904 93044 944
rect 92620 820 92660 860
rect 93964 652 94004 692
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
rect 94732 484 94772 524
rect 96652 1072 96692 1112
rect 99148 904 99188 944
rect 96268 568 96308 608
<< metal5 >>
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 38947 4180 38956 4220
rect 38996 4180 68524 4220
rect 68564 4180 68573 4220
rect 26083 4096 26092 4136
rect 26132 4096 66796 4136
rect 66836 4096 66845 4136
rect 28003 4012 28012 4052
rect 28052 4012 62380 4052
rect 62420 4012 62429 4052
rect 38659 3928 38668 3968
rect 38708 3928 66508 3968
rect 66548 3928 66557 3968
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 11107 3676 11116 3716
rect 11156 3676 17164 3716
rect 17204 3676 17213 3716
rect 66211 3592 66220 3632
rect 66260 3592 72460 3632
rect 72500 3592 72509 3632
rect 72931 3592 72940 3632
rect 72980 3592 79180 3632
rect 79220 3592 85324 3632
rect 85364 3592 85373 3632
rect 9571 3508 9580 3548
rect 9620 3508 15820 3548
rect 15860 3508 15869 3548
rect 19363 3508 19372 3548
rect 19412 3508 25324 3548
rect 25364 3508 31660 3548
rect 31700 3508 31709 3548
rect 41347 3508 41356 3548
rect 41396 3508 47596 3548
rect 47636 3508 47645 3548
rect 5923 3424 5932 3464
rect 5972 3424 11360 3464
rect 11320 3380 11360 3424
rect 32740 3424 35692 3464
rect 35732 3424 35741 3464
rect 64579 3424 64588 3464
rect 64628 3424 71308 3464
rect 71348 3424 71357 3464
rect 84547 3424 84556 3464
rect 84596 3424 90700 3464
rect 90740 3424 90749 3464
rect 32740 3380 32780 3424
rect 11320 3340 11500 3380
rect 11540 3340 17548 3380
rect 17588 3340 23788 3380
rect 23828 3340 29836 3380
rect 29876 3340 32780 3380
rect 55363 3340 55372 3380
rect 55412 3340 66220 3380
rect 66260 3340 66269 3380
rect 66595 3340 66604 3380
rect 66644 3340 72844 3380
rect 72884 3340 78604 3380
rect 78644 3340 78653 3380
rect 91459 3340 91468 3380
rect 91508 3340 97132 3380
rect 97172 3340 97181 3380
rect 6883 3172 6892 3212
rect 6932 3172 13036 3212
rect 13076 3172 19372 3212
rect 19412 3172 19421 3212
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 40195 3004 40204 3044
rect 40244 3004 44620 3044
rect 44660 3004 46540 3044
rect 46580 3004 46589 3044
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 18691 2920 18700 2960
rect 18740 2920 24844 2960
rect 24884 2920 24893 2960
rect 35299 2920 35308 2960
rect 35348 2920 40588 2960
rect 40628 2920 40637 2960
rect 80323 2920 80332 2960
rect 80372 2920 81920 2960
rect 81880 2876 81920 2920
rect 90140 2920 92812 2960
rect 92852 2920 92861 2960
rect 90140 2876 90180 2920
rect 17155 2836 17164 2876
rect 17204 2836 23404 2876
rect 23444 2836 23453 2876
rect 38755 2836 38764 2876
rect 38804 2836 44044 2876
rect 44084 2836 44093 2876
rect 46627 2836 46636 2876
rect 46676 2836 48076 2876
rect 48116 2836 48364 2876
rect 48404 2836 54508 2876
rect 54548 2836 54557 2876
rect 78595 2836 78604 2876
rect 78644 2836 81772 2876
rect 81812 2836 81821 2876
rect 81880 2836 86476 2876
rect 86516 2836 90180 2876
rect 90596 2836 91468 2876
rect 91508 2836 91517 2876
rect 90596 2792 90636 2836
rect 20419 2752 20428 2792
rect 20468 2752 26572 2792
rect 26612 2752 32236 2792
rect 32276 2752 32285 2792
rect 41635 2752 41644 2792
rect 41684 2752 42220 2792
rect 42260 2752 42269 2792
rect 46531 2752 46540 2792
rect 46580 2752 64588 2792
rect 64628 2752 64637 2792
rect 69187 2752 69196 2792
rect 69236 2752 74764 2792
rect 74804 2752 74813 2792
rect 76867 2752 76876 2792
rect 76916 2752 81580 2792
rect 81620 2752 81629 2792
rect 81871 2752 81880 2792
rect 81920 2752 84940 2792
rect 84980 2752 84989 2792
rect 85315 2752 85324 2792
rect 85364 2752 90636 2792
rect 90691 2752 90700 2792
rect 90740 2752 96364 2792
rect 96404 2752 96413 2792
rect 3500 2668 8044 2708
rect 8084 2668 14284 2708
rect 14324 2668 14333 2708
rect 15811 2668 15820 2708
rect 15860 2668 19044 2708
rect 24835 2668 24844 2708
rect 24884 2668 30892 2708
rect 30932 2668 36844 2708
rect 36884 2668 42988 2708
rect 43028 2668 49324 2708
rect 49364 2668 61324 2708
rect 61364 2668 67852 2708
rect 67892 2668 74284 2708
rect 74324 2668 80332 2708
rect 80372 2668 80381 2708
rect 81476 2668 88012 2708
rect 88052 2668 93676 2708
rect 93716 2668 93725 2708
rect 93859 2668 93868 2708
rect 93908 2668 95652 2708
rect 3500 2624 3540 2668
rect 19004 2624 19044 2668
rect 81476 2624 81516 2668
rect 95612 2624 95652 2668
rect 2275 2584 2284 2624
rect 2324 2584 3540 2624
rect 3907 2584 3916 2624
rect 3956 2584 6320 2624
rect 7171 2584 7180 2624
rect 7220 2584 12748 2624
rect 12788 2584 18700 2624
rect 18740 2584 18749 2624
rect 19004 2584 21868 2624
rect 21908 2584 28108 2624
rect 28148 2584 33772 2624
rect 33812 2584 40204 2624
rect 40244 2584 40253 2624
rect 40436 2584 41644 2624
rect 41684 2584 41693 2624
rect 41804 2584 41836 2624
rect 41876 2584 41885 2624
rect 42211 2584 42220 2624
rect 42260 2584 48460 2624
rect 48500 2584 54316 2624
rect 54356 2584 54365 2624
rect 54499 2584 54508 2624
rect 54548 2584 55980 2624
rect 64195 2584 64204 2624
rect 64244 2584 69772 2624
rect 69812 2584 75628 2624
rect 75668 2584 81484 2624
rect 81524 2584 81533 2624
rect 81880 2584 83404 2624
rect 83444 2584 89548 2624
rect 89588 2584 95116 2624
rect 95156 2584 95165 2624
rect 95612 2584 96748 2624
rect 96788 2584 96797 2624
rect 6280 2456 6320 2584
rect 9428 2500 9580 2540
rect 9620 2500 9629 2540
rect 23364 2500 23404 2540
rect 23444 2500 23453 2540
rect 35299 2500 35308 2540
rect 35348 2500 35357 2540
rect 9428 2456 9468 2500
rect 6280 2416 9468 2456
rect 23404 2456 23444 2500
rect 35308 2456 35348 2500
rect 40436 2456 40476 2584
rect 41804 2456 41844 2584
rect 46600 2500 46636 2540
rect 46676 2500 46685 2540
rect 46600 2456 46640 2500
rect 55940 2456 55980 2584
rect 81880 2540 81920 2584
rect 63692 2500 64300 2540
rect 64340 2500 64349 2540
rect 71299 2500 71308 2540
rect 71348 2500 71484 2540
rect 63692 2456 63732 2500
rect 71444 2456 71484 2500
rect 76840 2500 76876 2540
rect 76916 2500 76925 2540
rect 81571 2500 81580 2540
rect 81620 2500 81920 2540
rect 84931 2500 84940 2540
rect 84980 2500 84989 2540
rect 91052 2500 91084 2540
rect 91124 2500 91133 2540
rect 76840 2456 76880 2500
rect 23404 2416 29548 2456
rect 29588 2416 35348 2456
rect 35683 2416 35692 2456
rect 35732 2416 40476 2456
rect 40579 2416 40588 2456
rect 40628 2416 46640 2456
rect 54307 2416 54316 2456
rect 54356 2416 55460 2456
rect 55940 2416 63732 2456
rect 64240 2416 66988 2456
rect 67028 2416 67037 2456
rect 71444 2416 76880 2456
rect 84940 2456 84980 2500
rect 91052 2456 91092 2500
rect 84940 2416 91092 2456
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 55420 2288 55460 2416
rect 64240 2288 64280 2416
rect 55420 2248 64280 2288
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 46147 2080 46156 2120
rect 46196 2080 64684 2120
rect 64724 2080 64733 2120
rect 47875 1996 47884 2036
rect 47924 1996 65836 2036
rect 65876 1996 65885 2036
rect 50371 1912 50380 1952
rect 50420 1912 62572 1952
rect 62612 1912 62621 1952
rect 44995 1828 45004 1868
rect 45044 1828 63532 1868
rect 63572 1828 63581 1868
rect 45379 1660 45388 1700
rect 45428 1660 46060 1700
rect 46100 1660 54796 1700
rect 54836 1660 54845 1700
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 6692 1324 7564 1364
rect 7604 1324 7613 1364
rect 47971 1324 47980 1364
rect 48020 1324 48364 1364
rect 48404 1324 65740 1364
rect 65780 1324 65789 1364
rect 72931 1324 72940 1364
rect 72980 1324 76500 1364
rect 6692 1280 6732 1324
rect 76460 1280 76500 1324
rect 2500 1240 6732 1280
rect 6883 1240 6892 1280
rect 6932 1240 10060 1280
rect 10100 1240 10109 1280
rect 11395 1240 11404 1280
rect 11444 1240 12556 1280
rect 12596 1240 18700 1280
rect 18740 1240 24844 1280
rect 24884 1240 31084 1280
rect 31124 1240 37036 1280
rect 37076 1240 43276 1280
rect 43316 1240 49516 1280
rect 49556 1240 49565 1280
rect 54787 1240 54796 1280
rect 54836 1240 62668 1280
rect 62708 1240 62717 1280
rect 69379 1240 69388 1280
rect 69428 1240 75532 1280
rect 75572 1240 75581 1280
rect 76460 1240 78644 1280
rect 81475 1240 81484 1280
rect 81524 1240 87628 1280
rect 87668 1240 87677 1280
rect 87811 1240 87820 1280
rect 87860 1240 93196 1280
rect 93236 1240 93245 1280
rect 2500 1112 2540 1240
rect 78604 1196 78644 1240
rect 80978 1219 81102 1238
rect 80978 1196 80997 1219
rect 3956 1156 8332 1196
rect 8372 1156 8381 1196
rect 9884 1156 16012 1196
rect 16052 1156 22156 1196
rect 22196 1156 28204 1196
rect 28244 1156 34156 1196
rect 34196 1156 40300 1196
rect 40340 1156 40349 1196
rect 48067 1156 48076 1196
rect 48116 1156 49708 1196
rect 49748 1156 66604 1196
rect 66644 1156 66653 1196
rect 66787 1156 66796 1196
rect 66836 1156 72460 1196
rect 72500 1156 72509 1196
rect 72643 1156 72652 1196
rect 72692 1156 74764 1196
rect 74804 1156 74813 1196
rect 78595 1156 78604 1196
rect 78644 1156 80997 1196
rect 3956 1112 3996 1156
rect 9884 1112 9924 1156
rect 40394 1135 40518 1154
rect 1987 1072 1996 1112
rect 2036 1072 2540 1112
rect 2755 1072 2764 1112
rect 2804 1072 3996 1112
rect 4291 1072 4300 1112
rect 4340 1072 9868 1112
rect 9908 1072 9924 1112
rect 10051 1072 10060 1112
rect 10100 1072 12940 1112
rect 12980 1072 17548 1112
rect 17588 1072 17597 1112
rect 18092 1072 18316 1112
rect 18356 1072 24460 1112
rect 24500 1072 24509 1112
rect 25507 1072 25516 1112
rect 25556 1072 31468 1112
rect 31508 1072 31517 1112
rect 18092 1028 18132 1072
rect 40394 1049 40413 1135
rect 40499 1112 40518 1135
rect 80978 1133 80997 1156
rect 81083 1133 81102 1219
rect 80978 1114 81102 1133
rect 81880 1156 86860 1196
rect 86900 1156 93004 1196
rect 93044 1156 93053 1196
rect 40499 1072 40780 1112
rect 40820 1072 47020 1112
rect 47060 1072 49132 1112
rect 49172 1072 49181 1112
rect 49556 1072 59116 1112
rect 59156 1072 59165 1112
rect 63043 1072 63052 1112
rect 63092 1072 63532 1112
rect 63572 1072 69772 1112
rect 69812 1072 75916 1112
rect 75956 1072 80812 1112
rect 80852 1072 80861 1112
rect 40499 1049 40518 1072
rect 40394 1030 40518 1049
rect 49556 1028 49596 1072
rect 81880 1028 81920 1156
rect 87619 1072 87628 1112
rect 87668 1072 93580 1112
rect 93620 1072 93629 1112
rect 93676 1072 96652 1112
rect 96692 1072 96701 1112
rect 84626 1051 84750 1070
rect 84626 1028 84645 1051
rect 2500 988 6892 1028
rect 6932 988 6941 1028
rect 8323 988 8332 1028
rect 8372 988 12076 1028
rect 12116 988 12125 1028
rect 12259 988 12268 1028
rect 12308 988 18132 1028
rect 25891 988 25900 1028
rect 25940 988 31852 1028
rect 31892 988 31901 1028
rect 42691 988 42700 1028
rect 42740 988 48940 1028
rect 48980 988 49596 1028
rect 50179 988 50188 1028
rect 50228 988 64300 1028
rect 64340 988 70444 1028
rect 70484 988 73100 1028
rect 74755 988 74764 1028
rect 74804 988 79948 1028
rect 79988 988 81920 1028
rect 84547 988 84556 1028
rect 84596 988 84645 1028
rect 2500 944 2540 988
rect 73060 944 73100 988
rect 84626 965 84645 988
rect 84731 1028 84750 1051
rect 93676 1028 93716 1072
rect 84731 988 90700 1028
rect 90740 988 90749 1028
rect 92035 988 92044 1028
rect 92084 988 93716 1028
rect 84731 965 84750 988
rect 84626 946 84750 965
rect 1219 904 1228 944
rect 1268 904 2540 944
rect 4675 904 4684 944
rect 4724 904 10252 944
rect 10292 904 11212 944
rect 11252 904 11261 944
rect 11320 904 11404 944
rect 11444 904 11453 944
rect 16483 904 16492 944
rect 16532 904 17548 944
rect 17588 904 23788 944
rect 23828 904 23837 944
rect 24451 904 24460 944
rect 24500 904 30508 944
rect 30548 904 36460 944
rect 36500 904 36828 944
rect 37315 904 37324 944
rect 37364 904 43564 944
rect 43604 904 45388 944
rect 45428 904 45437 944
rect 49507 904 49516 944
rect 49556 904 61708 944
rect 61748 904 68620 944
rect 68660 904 72652 944
rect 72692 904 72701 944
rect 73060 904 74804 944
rect 74851 904 74860 944
rect 74900 904 80604 944
rect 80803 904 80812 944
rect 80852 904 81868 944
rect 81908 904 81917 944
rect 92995 904 93004 944
rect 93044 904 99148 944
rect 99188 904 99197 944
rect 11320 860 11360 904
rect 36788 860 36828 904
rect 74764 860 74804 904
rect 80564 860 80604 904
rect 6499 820 6508 860
rect 6548 820 11360 860
rect 20611 820 20620 860
rect 20660 820 26668 860
rect 26708 820 32620 860
rect 32660 820 32669 860
rect 36788 820 42700 860
rect 42740 820 42749 860
rect 66595 820 66604 860
rect 66644 820 67276 860
rect 67316 820 67325 860
rect 68035 820 68044 860
rect 68084 820 74380 860
rect 74420 820 74429 860
rect 74764 820 76684 860
rect 76724 820 76733 860
rect 80515 820 80524 860
rect 80564 820 86476 860
rect 86516 820 92620 860
rect 92660 820 92669 860
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 7555 736 7564 776
rect 7604 736 13708 776
rect 13748 736 19372 776
rect 19412 736 19421 776
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 35834 799 35958 818
rect 35834 776 35853 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 35011 736 35020 776
rect 35060 736 35853 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 35834 713 35853 736
rect 35939 713 35958 799
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 36067 736 36076 776
rect 36116 736 42028 776
rect 42068 736 48076 776
rect 48116 736 48125 776
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 35834 694 35958 713
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 65731 736 65740 776
rect 65780 736 72076 776
rect 72116 736 78220 776
rect 78260 736 78269 776
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
rect 28588 652 34444 692
rect 34484 652 34493 692
rect 40387 652 40396 692
rect 40436 652 46636 692
rect 46676 652 46685 692
rect 59107 652 59116 692
rect 59156 652 64280 692
rect 70531 652 70540 692
rect 70580 652 76300 692
rect 76340 652 76349 692
rect 81859 652 81868 692
rect 81908 652 83500 692
rect 83540 652 83549 692
rect 83756 652 86956 692
rect 86996 652 87820 692
rect 87860 652 87869 692
rect 88003 652 88012 692
rect 88052 652 93964 692
rect 94004 652 94013 692
rect 28588 608 28628 652
rect 1603 568 1612 608
rect 1652 568 7180 608
rect 7220 568 7229 608
rect 16387 568 16396 608
rect 16436 568 22540 608
rect 22580 568 28588 608
rect 28628 568 28637 608
rect 32611 568 32620 608
rect 32660 568 38860 608
rect 38900 568 42260 608
rect 42307 568 42316 608
rect 42356 568 43948 608
rect 43988 568 62764 608
rect 62804 568 62813 608
rect 7180 440 7220 568
rect 42220 524 42260 568
rect 64240 524 64280 652
rect 83756 608 83796 652
rect 66691 568 66700 608
rect 66740 568 68812 608
rect 68852 568 75148 608
rect 75188 568 75668 608
rect 75628 524 75668 568
rect 81880 568 83796 608
rect 84163 568 84172 608
rect 84212 568 90316 608
rect 90356 568 96268 608
rect 96308 568 96317 608
rect 81880 524 81920 568
rect 22915 484 22924 524
rect 22964 484 26188 524
rect 26228 484 26237 524
rect 29731 484 29740 524
rect 29780 484 36076 524
rect 36116 484 36125 524
rect 42220 484 45100 524
rect 45140 484 50188 524
rect 50228 484 50237 524
rect 64240 484 68044 524
rect 68084 484 68093 524
rect 75628 484 81100 524
rect 81140 484 81920 524
rect 82388 484 82636 524
rect 82676 484 88780 524
rect 88820 484 94732 524
rect 94772 484 94781 524
rect 62738 463 62862 482
rect 7180 400 13324 440
rect 13364 400 19276 440
rect 19316 400 19325 440
rect 34339 400 34348 440
rect 34388 400 35020 440
rect 35060 400 35069 440
rect 44498 379 44622 398
rect 44498 356 44517 379
rect 44419 316 44428 356
rect 44468 316 44517 356
rect 44498 293 44517 316
rect 44603 293 44622 379
rect 62738 377 62757 463
rect 62843 440 62862 463
rect 82388 440 82428 484
rect 62843 400 63052 440
rect 63092 400 63101 440
rect 76675 400 76684 440
rect 76724 400 82428 440
rect 83491 400 83500 440
rect 83540 400 88012 440
rect 88052 400 88061 440
rect 62843 377 62862 400
rect 62738 358 62862 377
rect 44498 274 44622 293
rect 14371 232 14380 272
rect 14420 232 20620 272
rect 20660 232 20669 272
rect 19651 64 19660 104
rect 19700 64 22924 104
rect 22964 64 22973 104
<< via5 >>
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 40413 1049 40499 1135
rect 80997 1133 81083 1219
rect 84645 965 84731 1051
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 35853 713 35939 799
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
rect 44517 293 44603 379
rect 62757 377 62843 463
<< metal6 >>
rect 3076 9115 3516 9198
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3666 3516 4493
rect 3076 3286 3106 3666
rect 3486 3286 3516 3666
rect 3076 3067 3516 3286
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 8359 4756 9116
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 4906 4756 5249
rect 4316 4526 4346 4906
rect 4726 4526 4756 4906
rect 4316 3823 4756 4526
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 9115 18636 9198
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3666 18636 4493
rect 18196 3286 18226 3666
rect 18606 3286 18636 3666
rect 18196 3067 18636 3286
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 8359 19876 9116
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 4906 19876 5249
rect 19436 4526 19466 4906
rect 19846 4526 19876 4906
rect 19436 3823 19876 4526
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 9115 33756 9198
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3666 33756 4493
rect 33316 3286 33346 3666
rect 33726 3286 33756 3666
rect 33316 3067 33756 3286
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 8359 34996 9116
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 4906 34996 5249
rect 34556 4526 34586 4906
rect 34966 4526 34996 4906
rect 34556 3823 34996 4526
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 48436 9115 48876 9198
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3666 48876 4493
rect 48436 3286 48466 3666
rect 48846 3286 48876 3666
rect 48436 3067 48876 3286
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 35732 799 36060 1010
rect 40292 928 40620 1010
rect 35732 713 35853 799
rect 35939 713 36060 799
rect 35732 592 36060 713
rect 48436 712 48876 1469
rect 49676 8359 50116 9116
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 4906 50116 5249
rect 49676 4526 49706 4906
rect 50086 4526 50116 4906
rect 49676 3823 50116 4526
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 9115 63996 9198
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3666 63996 4493
rect 63556 3286 63586 3666
rect 63966 3286 63996 3666
rect 63556 3067 63996 3286
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 8359 65236 9116
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 4906 65236 5249
rect 64796 4526 64826 4906
rect 65206 4526 65236 4906
rect 64796 3823 65236 4526
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 9115 79116 9198
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3666 79116 4493
rect 78676 3286 78706 3666
rect 79086 3286 79116 3666
rect 78676 3067 79116 3286
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 8359 80356 9116
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 4906 80356 5249
rect 79916 4526 79946 4906
rect 80326 4526 80356 4906
rect 79916 3823 80356 4526
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 93796 9115 94236 9198
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3666 94236 4493
rect 93796 3286 93826 3666
rect 94206 3286 94236 3666
rect 93796 3067 94236 3286
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 84524 965 84645 1010
rect 84731 965 84852 1010
rect 84524 844 84852 965
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 712 94236 1469
rect 95036 8359 95476 9116
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 4906 95476 5249
rect 95036 4526 95066 4906
rect 95446 4526 95476 4906
rect 95036 3823 95476 4526
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
rect 44396 172 44724 210
<< via6 >>
rect 3106 3286 3486 3666
rect 4346 4526 4726 4906
rect 18226 3286 18606 3666
rect 19466 4526 19846 4906
rect 33346 3286 33726 3666
rect 34586 4526 34966 4906
rect 48466 3286 48846 3666
rect 35706 1010 36086 1390
rect 40266 1135 40646 1390
rect 40266 1049 40413 1135
rect 40413 1049 40499 1135
rect 40499 1049 40646 1135
rect 40266 1010 40646 1049
rect 49706 4526 50086 4906
rect 63586 3286 63966 3666
rect 64826 4526 65206 4906
rect 78706 3286 79086 3666
rect 79946 4526 80326 4906
rect 93826 3286 94206 3666
rect 80850 1219 81230 1390
rect 80850 1133 80997 1219
rect 80997 1133 81083 1219
rect 81083 1133 81230 1219
rect 80850 1010 81230 1133
rect 84498 1051 84878 1390
rect 84498 1010 84645 1051
rect 84645 1010 84731 1051
rect 84731 1010 84878 1051
rect 95066 4526 95446 4906
rect 44370 379 44750 590
rect 44370 293 44517 379
rect 44517 293 44603 379
rect 44603 293 44750 379
rect 44370 210 44750 293
rect 62610 463 62990 590
rect 62610 377 62757 463
rect 62757 377 62843 463
rect 62843 377 62990 463
rect 62610 210 62990 377
<< metal7 >>
rect 532 4906 99404 4936
rect 532 4526 4346 4906
rect 4726 4526 19466 4906
rect 19846 4526 34586 4906
rect 34966 4526 49706 4906
rect 50086 4526 64826 4906
rect 65206 4526 79946 4906
rect 80326 4526 95066 4906
rect 95446 4526 99404 4906
rect 532 4496 99404 4526
rect 532 3666 99404 3696
rect 532 3286 3106 3666
rect 3486 3286 18226 3666
rect 18606 3286 33346 3666
rect 33726 3286 48466 3666
rect 48846 3286 63586 3666
rect 63966 3286 78706 3666
rect 79086 3286 93826 3666
rect 94206 3286 99404 3666
rect 532 3256 99404 3286
rect 35696 1390 40656 1400
rect 35696 1010 35706 1390
rect 36086 1010 40266 1390
rect 40646 1010 40656 1390
rect 35696 1000 40656 1010
rect 80840 1390 84888 1400
rect 80840 1010 80850 1390
rect 81230 1010 84498 1390
rect 84878 1010 84888 1390
rect 80840 1000 84888 1010
rect 44360 590 63000 600
rect 44360 210 44370 590
rect 44750 210 62610 590
rect 62990 210 63000 590
rect 44360 200 63000 210
use sg13g2_inv_1  _095_
timestamp 1676382929
transform -1 0 22560 0 -1 5292
box -48 -56 336 834
use sg13g2_nor2_1  _096_
timestamp 1676627187
transform -1 0 49536 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _097_
timestamp 1676627187
transform -1 0 44832 0 -1 6804
box -48 -56 432 834
use sg13g2_nor4_1  _098_
timestamp 1676643125
transform 1 0 46368 0 -1 6804
box -48 -56 624 834
use sg13g2_nor2b_1  _099_
timestamp 1685181386
transform 1 0 66816 0 -1 5292
box -54 -56 528 834
use sg13g2_and4_1  _100_
timestamp 1676985977
transform -1 0 62208 0 1 5292
box -48 -56 816 834
use sg13g2_nand4_1  _101_
timestamp 1685201930
transform -1 0 61440 0 1 5292
box -48 -56 624 834
use sg13g2_and2_1  _102_
timestamp 1676901763
transform -1 0 56544 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _103_
timestamp 1676557249
transform -1 0 56928 0 1 5292
box -48 -56 432 834
use sg13g2_and2_1  _104_
timestamp 1676901763
transform -1 0 48672 0 -1 6804
box -48 -56 528 834
use sg13g2_and2_1  _105_
timestamp 1676901763
transform 1 0 45696 0 -1 6804
box -48 -56 528 834
use sg13g2_nand2_1  _106_
timestamp 1676557249
transform -1 0 50784 0 1 5292
box -48 -56 432 834
use sg13g2_nor2b_1  _107_
timestamp 1685181386
transform 1 0 73728 0 -1 5292
box -54 -56 528 834
use sg13g2_and3_1  _108_
timestamp 1676971669
transform 1 0 61632 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _109_
timestamp 1683988354
transform 1 0 61152 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _110_
timestamp 1676627187
transform 1 0 55872 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2b_1  _111_
timestamp 1676567195
transform 1 0 56256 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _112_
timestamp 1685181386
transform 1 0 40992 0 1 5292
box -54 -56 528 834
use sg13g2_nand2_1  _113_
timestamp 1676557249
transform -1 0 50880 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _114_
timestamp 1676627187
transform -1 0 57216 0 -1 3780
box -48 -56 432 834
use sg13g2_or2_1  _115_
timestamp 1684236171
transform -1 0 56832 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _116_
timestamp 1685181386
transform -1 0 42144 0 -1 6804
box -54 -56 528 834
use sg13g2_nand2_1  _117_
timestamp 1676557249
transform 1 0 50112 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _118_
timestamp 1676627187
transform 1 0 56160 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _119_
timestamp 1684236171
transform 1 0 56544 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _120_
timestamp 1676557249
transform 1 0 50880 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _121_
timestamp 1676627187
transform 1 0 56928 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _122_
timestamp 1684236171
transform 1 0 57024 0 1 756
box -48 -56 528 834
use sg13g2_nor2b_1  _123_
timestamp 1685181386
transform -1 0 48000 0 -1 6804
box -54 -56 528 834
use sg13g2_nand2_1  _124_
timestamp 1676557249
transform -1 0 52512 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _125_
timestamp 1676627187
transform -1 0 58176 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _126_
timestamp 1684236171
transform 1 0 57312 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _127_
timestamp 1676557249
transform 1 0 52512 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _128_
timestamp 1676627187
transform -1 0 58464 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _129_
timestamp 1684236171
transform 1 0 57600 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _130_
timestamp 1676557249
transform 1 0 51840 0 1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _131_
timestamp 1676627187
transform -1 0 58464 0 1 5292
box -48 -56 432 834
use sg13g2_or2_1  _132_
timestamp 1684236171
transform 1 0 57984 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _133_
timestamp 1676557249
transform 1 0 52512 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _134_
timestamp 1676627187
transform -1 0 59040 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _135_
timestamp 1684236171
transform 1 0 58464 0 1 2268
box -48 -56 528 834
use sg13g2_nor2b_1  _136_
timestamp 1685181386
transform -1 0 49152 0 -1 6804
box -54 -56 528 834
use sg13g2_nand2_1  _137_
timestamp 1676557249
transform -1 0 53856 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _138_
timestamp 1676627187
transform -1 0 59712 0 1 3780
box -48 -56 432 834
use sg13g2_or2_1  _139_
timestamp 1684236171
transform 1 0 58848 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _140_
timestamp 1676557249
transform -1 0 55200 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _141_
timestamp 1676627187
transform 1 0 59040 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _142_
timestamp 1684236171
transform 1 0 59424 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _143_
timestamp 1676557249
transform -1 0 55584 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _144_
timestamp 1676627187
transform 1 0 59904 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _145_
timestamp 1684236171
transform -1 0 60384 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _146_
timestamp 1676557249
transform -1 0 53568 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _147_
timestamp 1676627187
transform -1 0 61248 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _148_
timestamp 1684236171
transform -1 0 60864 0 1 756
box -48 -56 528 834
use sg13g2_nand2_1  _149_
timestamp 1676557249
transform 1 0 54240 0 1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _150_
timestamp 1676627187
transform -1 0 61152 0 -1 5292
box -48 -56 432 834
use sg13g2_or2_1  _151_
timestamp 1684236171
transform 1 0 60288 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _152_
timestamp 1676557249
transform -1 0 58848 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _153_
timestamp 1676627187
transform 1 0 60384 0 1 2268
box -48 -56 432 834
use sg13g2_or2_1  _154_
timestamp 1684236171
transform 1 0 60768 0 1 2268
box -48 -56 528 834
use sg13g2_nand2_1  _155_
timestamp 1676557249
transform -1 0 58464 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _156_
timestamp 1676627187
transform -1 0 62112 0 1 2268
box -48 -56 432 834
use sg13g2_or2_1  _157_
timestamp 1684236171
transform 1 0 61248 0 1 2268
box -48 -56 528 834
use sg13g2_and2_1  _158_
timestamp 1676901763
transform 1 0 61728 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _159_
timestamp 1676557249
transform -1 0 62592 0 1 3780
box -48 -56 432 834
use sg13g2_nor2b_1  _160_
timestamp 1685181386
transform -1 0 73728 0 -1 5292
box -54 -56 528 834
use sg13g2_and2_1  _161_
timestamp 1676901763
transform -1 0 66720 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _162_
timestamp 1676557249
transform -1 0 67104 0 1 3780
box -48 -56 432 834
use sg13g2_and3_1  _163_
timestamp 1676971669
transform 1 0 45600 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _164_
timestamp 1683988354
transform -1 0 46464 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _165_
timestamp 1676627187
transform -1 0 62976 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _166_
timestamp 1676557249
transform 1 0 62496 0 -1 2268
box -48 -56 432 834
use sg13g2_and3_1  _167_
timestamp 1676971669
transform -1 0 42336 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _168_
timestamp 1683988354
transform -1 0 42720 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _169_
timestamp 1676627187
transform -1 0 63360 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _170_
timestamp 1676557249
transform -1 0 63168 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  _171_
timestamp 1676971669
transform -1 0 41760 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _172_
timestamp 1683988354
transform -1 0 43296 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _173_
timestamp 1676627187
transform -1 0 63744 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _174_
timestamp 1676557249
transform -1 0 63456 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _175_
timestamp 1676971669
transform -1 0 44640 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _176_
timestamp 1683988354
transform -1 0 45216 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _177_
timestamp 1676627187
transform -1 0 64128 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _178_
timestamp 1676557249
transform -1 0 63648 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  _179_
timestamp 1676971669
transform -1 0 46944 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _180_
timestamp 1683988354
transform -1 0 46464 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _181_
timestamp 1676627187
transform -1 0 64512 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _182_
timestamp 1676557249
transform -1 0 64128 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _183_
timestamp 1676971669
transform -1 0 42144 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _184_
timestamp 1683988354
transform -1 0 41664 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _185_
timestamp 1676627187
transform -1 0 64896 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _186_
timestamp 1676557249
transform -1 0 64512 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _187_
timestamp 1676971669
transform -1 0 42432 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _188_
timestamp 1683988354
transform -1 0 42816 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _189_
timestamp 1676627187
transform -1 0 65280 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _190_
timestamp 1676557249
transform -1 0 64896 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _191_
timestamp 1676971669
transform -1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _192_
timestamp 1683988354
transform -1 0 44736 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _193_
timestamp 1676627187
transform -1 0 65664 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _194_
timestamp 1676557249
transform -1 0 65184 0 -1 2268
box -48 -56 432 834
use sg13g2_and3_1  _195_
timestamp 1676971669
transform -1 0 52896 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _196_
timestamp 1683988354
transform -1 0 49056 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _197_
timestamp 1676627187
transform -1 0 66048 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _198_
timestamp 1676557249
transform -1 0 65568 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _199_
timestamp 1676971669
transform 1 0 47808 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _200_
timestamp 1683988354
transform -1 0 51648 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _201_
timestamp 1676627187
transform -1 0 66432 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _202_
timestamp 1676557249
transform -1 0 65952 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _203_
timestamp 1676971669
transform -1 0 55872 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _204_
timestamp 1683988354
transform -1 0 55488 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _205_
timestamp 1676627187
transform -1 0 66816 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _206_
timestamp 1676557249
transform -1 0 66336 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _207_
timestamp 1676971669
transform -1 0 49152 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _208_
timestamp 1683988354
transform -1 0 48576 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _209_
timestamp 1676627187
transform -1 0 67200 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _210_
timestamp 1676557249
transform -1 0 66720 0 -1 2268
box -48 -56 432 834
use sg13g2_and3_1  _211_
timestamp 1676971669
transform -1 0 54048 0 1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _212_
timestamp 1683988354
transform -1 0 49728 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _213_
timestamp 1676627187
transform -1 0 67584 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _214_
timestamp 1676557249
transform -1 0 67104 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _215_
timestamp 1676971669
transform -1 0 59040 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _216_
timestamp 1683988354
transform 1 0 58944 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _217_
timestamp 1676627187
transform -1 0 67968 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _218_
timestamp 1676557249
transform -1 0 67488 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _219_
timestamp 1676971669
transform -1 0 58368 0 -1 5292
box -48 -56 720 834
use sg13g2_nand3_1  _220_
timestamp 1683988354
transform 1 0 58464 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _221_
timestamp 1676627187
transform -1 0 68352 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _222_
timestamp 1676557249
transform 1 0 67296 0 1 2268
box -48 -56 432 834
use sg13g2_and2_1  _223_
timestamp 1676901763
transform -1 0 61728 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _224_
timestamp 1676557249
transform -1 0 61920 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _225_
timestamp 1676627187
transform 1 0 68352 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _226_
timestamp 1676557249
transform -1 0 67968 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _227_
timestamp 1676627187
transform -1 0 74592 0 -1 5292
box -48 -56 432 834
use sg13g2_and2_1  _228_
timestamp 1676901763
transform 1 0 68352 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _229_
timestamp 1676557249
transform -1 0 69216 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _230_
timestamp 1676627187
transform 1 0 68736 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _231_
timestamp 1676557249
transform -1 0 68928 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _232_
timestamp 1676627187
transform -1 0 69504 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _233_
timestamp 1676557249
transform -1 0 69312 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _234_
timestamp 1676627187
transform -1 0 69888 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _235_
timestamp 1676557249
transform -1 0 69696 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _236_
timestamp 1676627187
transform -1 0 70272 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _237_
timestamp 1676557249
transform -1 0 70080 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _238_
timestamp 1676627187
transform -1 0 70656 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _239_
timestamp 1676557249
transform -1 0 70464 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _240_
timestamp 1676627187
transform -1 0 71040 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _241_
timestamp 1676557249
transform -1 0 70848 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _242_
timestamp 1676627187
transform -1 0 71424 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _243_
timestamp 1676557249
transform -1 0 71232 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _244_
timestamp 1676627187
transform -1 0 71808 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _245_
timestamp 1676557249
transform -1 0 71616 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _246_
timestamp 1676627187
transform -1 0 72192 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _247_
timestamp 1676557249
transform -1 0 72000 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _248_
timestamp 1676627187
transform -1 0 72576 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _249_
timestamp 1676557249
transform -1 0 72384 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _250_
timestamp 1676627187
transform -1 0 72960 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _251_
timestamp 1676557249
transform -1 0 72768 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _252_
timestamp 1676627187
transform -1 0 73344 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _253_
timestamp 1676557249
transform -1 0 73152 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _254_
timestamp 1676627187
transform -1 0 73728 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _255_
timestamp 1676557249
transform -1 0 73248 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _256_
timestamp 1676627187
transform -1 0 74112 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _257_
timestamp 1676557249
transform -1 0 73632 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _258_
timestamp 1676627187
transform -1 0 74496 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _259_
timestamp 1676557249
transform -1 0 74016 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _260_
timestamp 1676627187
transform -1 0 74880 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _261_
timestamp 1676557249
transform 1 0 74016 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _262_
timestamp 1676627187
transform -1 0 82464 0 -1 5292
box -48 -56 432 834
use sg13g2_and3_1  _263_
timestamp 1676971669
transform 1 0 74496 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _264_
timestamp 1683988354
transform -1 0 74496 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _265_
timestamp 1676627187
transform -1 0 75264 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _266_
timestamp 1676557249
transform -1 0 75072 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _267_
timestamp 1676627187
transform -1 0 75648 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _268_
timestamp 1676557249
transform -1 0 75264 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _269_
timestamp 1676627187
transform -1 0 76032 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _270_
timestamp 1676557249
transform -1 0 75648 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _271_
timestamp 1676627187
transform -1 0 76416 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _272_
timestamp 1676557249
transform -1 0 75936 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _273_
timestamp 1676627187
transform -1 0 76800 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _274_
timestamp 1676557249
transform -1 0 76320 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _275_
timestamp 1676627187
transform -1 0 77184 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _276_
timestamp 1676557249
transform -1 0 76704 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _277_
timestamp 1676627187
transform -1 0 77568 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _278_
timestamp 1676557249
transform -1 0 77088 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _279_
timestamp 1676627187
transform -1 0 77952 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _280_
timestamp 1676557249
transform 1 0 76992 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _281_
timestamp 1676627187
transform -1 0 78336 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _282_
timestamp 1676557249
transform 1 0 77376 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _283_
timestamp 1676627187
transform -1 0 78720 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _284_
timestamp 1676557249
transform -1 0 78240 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _285_
timestamp 1676627187
transform -1 0 79104 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _286_
timestamp 1676557249
transform -1 0 78624 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _287_
timestamp 1676627187
transform -1 0 79488 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _288_
timestamp 1676557249
transform 1 0 78528 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _289_
timestamp 1676627187
transform -1 0 79872 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _290_
timestamp 1676557249
transform 1 0 78912 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _291_
timestamp 1676627187
transform -1 0 80256 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _292_
timestamp 1676557249
transform 1 0 79296 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _293_
timestamp 1676627187
transform -1 0 80640 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _294_
timestamp 1676557249
transform 1 0 79680 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _295_
timestamp 1676627187
transform 1 0 79872 0 -1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _296_
timestamp 1676557249
transform 1 0 80064 0 -1 3780
box -48 -56 432 834
use sg13g2_and2_1  _297_
timestamp 1676901763
transform 1 0 80640 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _298_
timestamp 1676557249
transform 1 0 80256 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _299_
timestamp 1676627187
transform -1 0 81216 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _300_
timestamp 1676557249
transform -1 0 81120 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _301_
timestamp 1676627187
transform -1 0 81600 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _302_
timestamp 1676557249
transform -1 0 81408 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _303_
timestamp 1676627187
transform -1 0 81984 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _304_
timestamp 1676557249
transform -1 0 81792 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _305_
timestamp 1676627187
transform -1 0 82368 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _306_
timestamp 1676557249
transform 1 0 81600 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _307_
timestamp 1676627187
transform -1 0 82752 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _308_
timestamp 1676557249
transform -1 0 82464 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _309_
timestamp 1676627187
transform -1 0 83136 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _310_
timestamp 1676557249
transform -1 0 82848 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _311_
timestamp 1676627187
transform -1 0 83520 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _312_
timestamp 1676557249
transform -1 0 83232 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _313_
timestamp 1676627187
transform -1 0 83904 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _314_
timestamp 1676557249
transform 1 0 83136 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _315_
timestamp 1676627187
transform -1 0 84288 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _316_
timestamp 1676557249
transform 1 0 83520 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _317_
timestamp 1676627187
transform -1 0 84672 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _318_
timestamp 1676557249
transform 1 0 83904 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _319_
timestamp 1676627187
transform -1 0 85056 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _320_
timestamp 1676557249
transform 1 0 84288 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _321_
timestamp 1676627187
transform -1 0 85440 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _322_
timestamp 1676557249
transform 1 0 84672 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _323_
timestamp 1676627187
transform -1 0 85824 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _324_
timestamp 1676557249
transform 1 0 85056 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _325_
timestamp 1676627187
transform -1 0 86208 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _326_
timestamp 1676557249
transform 1 0 85440 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _327_
timestamp 1676627187
transform -1 0 86592 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _328_
timestamp 1676557249
transform 1 0 85824 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _329_
timestamp 1676627187
transform -1 0 86976 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _330_
timestamp 1676557249
transform 1 0 86208 0 1 2268
box -48 -56 432 834
use sg13g2_and2_1  _331_
timestamp 1676901763
transform 1 0 86496 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _332_
timestamp 1676557249
transform -1 0 87360 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _333_
timestamp 1676627187
transform 1 0 86976 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _334_
timestamp 1676557249
transform -1 0 87168 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _335_
timestamp 1676627187
transform -1 0 87744 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _336_
timestamp 1676557249
transform -1 0 87552 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _337_
timestamp 1676627187
transform -1 0 88128 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _338_
timestamp 1676557249
transform -1 0 87936 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _339_
timestamp 1676627187
transform -1 0 88512 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _340_
timestamp 1676557249
transform -1 0 88320 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _341_
timestamp 1676627187
transform -1 0 88896 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _342_
timestamp 1676557249
transform -1 0 88704 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _343_
timestamp 1676627187
transform -1 0 89280 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _344_
timestamp 1676557249
transform -1 0 89088 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _345_
timestamp 1676627187
transform -1 0 89664 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _346_
timestamp 1676557249
transform -1 0 89472 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _347_
timestamp 1676627187
transform -1 0 90048 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _348_
timestamp 1676557249
transform -1 0 89856 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _349_
timestamp 1676627187
transform -1 0 90432 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _350_
timestamp 1676557249
transform -1 0 90240 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _351_
timestamp 1676627187
transform -1 0 90816 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _352_
timestamp 1676557249
transform -1 0 90624 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _353_
timestamp 1676627187
transform -1 0 91200 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _354_
timestamp 1676557249
transform -1 0 91008 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _355_
timestamp 1676627187
transform -1 0 91584 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _356_
timestamp 1676557249
transform -1 0 91392 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _357_
timestamp 1676627187
transform -1 0 91968 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _358_
timestamp 1676557249
transform -1 0 91776 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _359_
timestamp 1676627187
transform -1 0 92352 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _360_
timestamp 1676557249
transform -1 0 92160 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _361_
timestamp 1676627187
transform -1 0 92736 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _362_
timestamp 1676557249
transform -1 0 92544 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _363_
timestamp 1676627187
transform -1 0 93120 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _364_
timestamp 1676557249
transform 1 0 92544 0 -1 3780
box -48 -56 432 834
use sg13g2_and2_1  _365_
timestamp 1676901763
transform 1 0 91872 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _366_
timestamp 1676557249
transform 1 0 91488 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _367_
timestamp 1676627187
transform 1 0 93120 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _368_
timestamp 1676557249
transform -1 0 92832 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _369_
timestamp 1676627187
transform 1 0 93504 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _370_
timestamp 1676557249
transform -1 0 93216 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _371_
timestamp 1676627187
transform 1 0 93888 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _372_
timestamp 1676557249
transform -1 0 93600 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _373_
timestamp 1676627187
transform 1 0 94272 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _374_
timestamp 1676557249
transform -1 0 93888 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _375_
timestamp 1676627187
transform 1 0 94656 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _376_
timestamp 1676557249
transform -1 0 94368 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _377_
timestamp 1676627187
transform 1 0 95040 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _378_
timestamp 1676557249
transform -1 0 94752 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _379_
timestamp 1676627187
transform 1 0 95424 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _380_
timestamp 1676557249
transform -1 0 95136 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _381_
timestamp 1676627187
transform 1 0 95808 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _382_
timestamp 1676557249
transform -1 0 95424 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _383_
timestamp 1676627187
transform 1 0 96192 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _384_
timestamp 1676557249
transform -1 0 95808 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _385_
timestamp 1676627187
transform 1 0 96576 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _386_
timestamp 1676557249
transform -1 0 96288 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _387_
timestamp 1676627187
transform 1 0 96960 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _388_
timestamp 1676557249
transform -1 0 96672 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _389_
timestamp 1676627187
transform 1 0 97344 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _390_
timestamp 1676557249
transform -1 0 97056 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _391_
timestamp 1676627187
transform 1 0 97728 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _392_
timestamp 1676557249
transform -1 0 97440 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _393_
timestamp 1676627187
transform 1 0 98112 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _394_
timestamp 1676557249
transform -1 0 97824 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _395_
timestamp 1676627187
transform 1 0 98496 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _396_
timestamp 1676557249
transform 1 0 97824 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _397_
timestamp 1676627187
transform -1 0 99264 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _398_
timestamp 1676557249
transform 1 0 97824 0 -1 2268
box -48 -56 432 834
use sg13g2_and3_1  _399_
timestamp 1676971669
transform -1 0 19392 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _400_
timestamp 1683988354
transform -1 0 19296 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _401_
timestamp 1676627187
transform 1 0 6720 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _402_
timestamp 1676557249
transform -1 0 7200 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _403_
timestamp 1676627187
transform 1 0 7104 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _404_
timestamp 1676557249
transform -1 0 7584 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _405_
timestamp 1676627187
transform 1 0 7488 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _406_
timestamp 1676557249
transform -1 0 7968 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _407_
timestamp 1676627187
transform 1 0 7872 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _408_
timestamp 1676557249
transform -1 0 8352 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _409_
timestamp 1676627187
transform 1 0 8256 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _410_
timestamp 1676557249
transform -1 0 8736 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _411_
timestamp 1676627187
transform 1 0 8640 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _412_
timestamp 1676557249
transform -1 0 9120 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _413_
timestamp 1676627187
transform 1 0 9024 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _414_
timestamp 1676557249
transform -1 0 9504 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _415_
timestamp 1676627187
transform 1 0 9408 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _416_
timestamp 1676557249
transform -1 0 9888 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _417_
timestamp 1676627187
transform 1 0 9792 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _418_
timestamp 1676557249
transform -1 0 10272 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _419_
timestamp 1676627187
transform 1 0 10176 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _420_
timestamp 1676557249
transform -1 0 10656 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _421_
timestamp 1676627187
transform 1 0 10560 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _422_
timestamp 1676557249
transform -1 0 11040 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _423_
timestamp 1676627187
transform 1 0 10944 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _424_
timestamp 1676557249
transform -1 0 11424 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _425_
timestamp 1676627187
transform 1 0 11328 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _426_
timestamp 1676557249
transform -1 0 11808 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _427_
timestamp 1676627187
transform 1 0 11712 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _428_
timestamp 1676557249
transform -1 0 12192 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _429_
timestamp 1676627187
transform 1 0 12096 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _430_
timestamp 1676557249
transform -1 0 12576 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _431_
timestamp 1676627187
transform 1 0 12480 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _432_
timestamp 1676557249
transform 1 0 12480 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  _433_
timestamp 1676971669
transform -1 0 18720 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _434_
timestamp 1683988354
transform -1 0 19872 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _435_
timestamp 1676627187
transform 1 0 12864 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _436_
timestamp 1676557249
transform -1 0 13344 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _437_
timestamp 1676627187
transform 1 0 13248 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _438_
timestamp 1676557249
transform -1 0 13728 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _439_
timestamp 1676627187
transform 1 0 13632 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _440_
timestamp 1676557249
transform -1 0 14112 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _441_
timestamp 1676627187
transform 1 0 14016 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _442_
timestamp 1676557249
transform 1 0 14016 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _443_
timestamp 1676627187
transform 1 0 14400 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _444_
timestamp 1676557249
transform 1 0 14208 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _445_
timestamp 1676627187
transform 1 0 14784 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _446_
timestamp 1676557249
transform 1 0 14592 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _447_
timestamp 1676627187
transform 1 0 15168 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _448_
timestamp 1676557249
transform 1 0 14976 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _449_
timestamp 1676627187
transform 1 0 15552 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _450_
timestamp 1676557249
transform 1 0 15360 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _451_
timestamp 1676627187
transform 1 0 15936 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _452_
timestamp 1676557249
transform 1 0 15744 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _453_
timestamp 1676627187
transform 1 0 16320 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _454_
timestamp 1676557249
transform 1 0 16128 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _455_
timestamp 1676627187
transform 1 0 16704 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _456_
timestamp 1676557249
transform 1 0 16512 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _457_
timestamp 1676627187
transform 1 0 17088 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _458_
timestamp 1676557249
transform 1 0 16896 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _459_
timestamp 1676627187
transform 1 0 17472 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _460_
timestamp 1676557249
transform 1 0 17280 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _461_
timestamp 1676627187
transform 1 0 17856 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _462_
timestamp 1676557249
transform 1 0 17664 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _463_
timestamp 1676627187
transform 1 0 18240 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _464_
timestamp 1676557249
transform 1 0 18048 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _465_
timestamp 1676627187
transform 1 0 18624 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _466_
timestamp 1676557249
transform 1 0 18432 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _467_
timestamp 1676971669
transform 1 0 24096 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _468_
timestamp 1683988354
transform -1 0 25248 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _469_
timestamp 1676627187
transform 1 0 19008 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _470_
timestamp 1676557249
transform -1 0 19680 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _471_
timestamp 1676627187
transform 1 0 19392 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _472_
timestamp 1676557249
transform -1 0 19968 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _473_
timestamp 1676627187
transform 1 0 19776 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _474_
timestamp 1676557249
transform -1 0 20256 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _475_
timestamp 1676627187
transform 1 0 20160 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _476_
timestamp 1676557249
transform 1 0 20160 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _477_
timestamp 1676627187
transform 1 0 20544 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _478_
timestamp 1676557249
transform -1 0 21024 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _479_
timestamp 1676627187
transform 1 0 20928 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _480_
timestamp 1676557249
transform -1 0 21408 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _481_
timestamp 1676627187
transform 1 0 21312 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _482_
timestamp 1676557249
transform -1 0 21792 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _483_
timestamp 1676627187
transform 1 0 21696 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _484_
timestamp 1676557249
transform -1 0 22176 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _485_
timestamp 1676627187
transform 1 0 22080 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _486_
timestamp 1676557249
transform 1 0 22080 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _487_
timestamp 1676627187
transform 1 0 22464 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _488_
timestamp 1676557249
transform 1 0 22464 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _489_
timestamp 1676627187
transform 1 0 22848 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _490_
timestamp 1676557249
transform 1 0 22848 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _491_
timestamp 1676627187
transform 1 0 23232 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _492_
timestamp 1676557249
transform -1 0 23712 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _493_
timestamp 1676627187
transform 1 0 23616 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _494_
timestamp 1676557249
transform 1 0 23520 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _495_
timestamp 1676627187
transform 1 0 24000 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _496_
timestamp 1676557249
transform 1 0 23904 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _497_
timestamp 1676627187
transform 1 0 24384 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _498_
timestamp 1676557249
transform 1 0 24288 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _499_
timestamp 1676627187
transform 1 0 24768 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _500_
timestamp 1676557249
transform 1 0 24576 0 -1 2268
box -48 -56 432 834
use sg13g2_nand3_1  _501_
timestamp 1683988354
transform -1 0 62784 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _502_
timestamp 1676627187
transform -1 0 26208 0 1 3780
box -48 -56 432 834
use sg13g2_nand2b_1  _503_
timestamp 1676567195
transform -1 0 28128 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _504_
timestamp 1676627187
transform -1 0 26208 0 -1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _505_
timestamp 1676557249
transform -1 0 25632 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _506_
timestamp 1676627187
transform 1 0 25440 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _507_
timestamp 1676557249
transform -1 0 26016 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _508_
timestamp 1676627187
transform 1 0 25824 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _509_
timestamp 1676557249
transform -1 0 26400 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _510_
timestamp 1676627187
transform 1 0 26208 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _511_
timestamp 1676557249
transform 1 0 26304 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _512_
timestamp 1676627187
transform 1 0 26592 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _513_
timestamp 1676557249
transform 1 0 26688 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _514_
timestamp 1676627187
transform 1 0 26976 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _515_
timestamp 1676557249
transform 1 0 27072 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _516_
timestamp 1676627187
transform 1 0 27360 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _517_
timestamp 1676557249
transform -1 0 27936 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _518_
timestamp 1676627187
transform 1 0 27744 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _519_
timestamp 1676557249
transform 1 0 27840 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _520_
timestamp 1676627187
transform 1 0 28128 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _521_
timestamp 1676557249
transform -1 0 28704 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _522_
timestamp 1676627187
transform 1 0 28512 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _523_
timestamp 1676557249
transform -1 0 29088 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _524_
timestamp 1676627187
transform 1 0 28896 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _525_
timestamp 1676557249
transform -1 0 29472 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _526_
timestamp 1676627187
transform 1 0 29280 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _527_
timestamp 1676557249
transform -1 0 29856 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _528_
timestamp 1676627187
transform 1 0 29664 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _529_
timestamp 1676557249
transform 1 0 29568 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _530_
timestamp 1676627187
transform 1 0 30048 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _531_
timestamp 1676557249
transform 1 0 29952 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _532_
timestamp 1676627187
transform 1 0 30432 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _533_
timestamp 1676557249
transform 1 0 30336 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _534_
timestamp 1676627187
transform -1 0 31200 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _535_
timestamp 1676557249
transform 1 0 30624 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  _536_
timestamp 1676971669
transform -1 0 32544 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _537_
timestamp 1683988354
transform -1 0 33024 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _538_
timestamp 1676627187
transform -1 0 32256 0 -1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _539_
timestamp 1676557249
transform -1 0 31968 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _540_
timestamp 1676627187
transform 1 0 31392 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _541_
timestamp 1676557249
transform -1 0 31584 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _542_
timestamp 1676627187
transform 1 0 31776 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _543_
timestamp 1676557249
transform 1 0 31584 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _544_
timestamp 1676627187
transform 1 0 32160 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _545_
timestamp 1676557249
transform 1 0 31968 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _546_
timestamp 1676627187
transform 1 0 32544 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _547_
timestamp 1676557249
transform 1 0 32352 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _548_
timestamp 1676627187
transform 1 0 32928 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _549_
timestamp 1676557249
transform 1 0 32736 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _550_
timestamp 1676627187
transform 1 0 33312 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _551_
timestamp 1676557249
transform 1 0 33120 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _552_
timestamp 1676627187
transform 1 0 33696 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _553_
timestamp 1676557249
transform 1 0 33504 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _554_
timestamp 1676627187
transform 1 0 34080 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _555_
timestamp 1676557249
transform 1 0 33888 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _556_
timestamp 1676627187
transform 1 0 34464 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _557_
timestamp 1676557249
transform 1 0 34272 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _558_
timestamp 1676627187
transform 1 0 34848 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _559_
timestamp 1676557249
transform 1 0 34656 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _560_
timestamp 1676627187
transform 1 0 35232 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _561_
timestamp 1676557249
transform 1 0 35040 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _562_
timestamp 1676627187
transform 1 0 35616 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _563_
timestamp 1676557249
transform 1 0 35424 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _564_
timestamp 1676627187
transform 1 0 36000 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _565_
timestamp 1676557249
transform 1 0 35808 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _566_
timestamp 1676627187
transform 1 0 36384 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _567_
timestamp 1676557249
transform 1 0 36192 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _568_
timestamp 1676627187
transform -1 0 37152 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _569_
timestamp 1676557249
transform 1 0 36576 0 -1 3780
box -48 -56 432 834
use sg13g2_and3_1  _570_
timestamp 1676971669
transform 1 0 36960 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _571_
timestamp 1683988354
transform -1 0 38208 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _572_
timestamp 1676627187
transform 1 0 37248 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _573_
timestamp 1676557249
transform -1 0 37920 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _574_
timestamp 1676627187
transform 1 0 37632 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _575_
timestamp 1676557249
transform -1 0 38592 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _576_
timestamp 1676627187
transform 1 0 38016 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _577_
timestamp 1676557249
transform 1 0 38112 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _578_
timestamp 1676627187
transform 1 0 38400 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _579_
timestamp 1676557249
transform 1 0 38496 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _580_
timestamp 1676627187
transform 1 0 38784 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _581_
timestamp 1676557249
transform 1 0 38784 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _582_
timestamp 1676627187
transform 1 0 39168 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _583_
timestamp 1676557249
transform 1 0 39168 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _584_
timestamp 1676627187
transform 1 0 39552 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _585_
timestamp 1676557249
transform 1 0 39552 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _586_
timestamp 1676627187
transform 1 0 39936 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _587_
timestamp 1676557249
transform 1 0 39936 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _588_
timestamp 1676627187
transform 1 0 40320 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _589_
timestamp 1676557249
transform 1 0 40224 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _590_
timestamp 1676627187
transform 1 0 40704 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _591_
timestamp 1676557249
transform 1 0 40704 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _592_
timestamp 1676627187
transform 1 0 41088 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _593_
timestamp 1676557249
transform 1 0 41088 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _594_
timestamp 1676627187
transform 1 0 41472 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _595_
timestamp 1676557249
transform 1 0 41568 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _596_
timestamp 1676627187
transform 1 0 41856 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _597_
timestamp 1676557249
transform 1 0 41952 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _598_
timestamp 1676627187
transform 1 0 42240 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _599_
timestamp 1676557249
transform 1 0 41856 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _600_
timestamp 1676627187
transform 1 0 42624 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _601_
timestamp 1676557249
transform 1 0 42720 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _602_
timestamp 1676627187
transform -1 0 43392 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _603_
timestamp 1676557249
transform 1 0 42720 0 1 2268
box -48 -56 432 834
use sg13g2_and3_1  _604_
timestamp 1676971669
transform 1 0 38112 0 1 3780
box -48 -56 720 834
use sg13g2_nand3_1  _605_
timestamp 1683988354
transform 1 0 37632 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _606_
timestamp 1676627187
transform 1 0 43488 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _607_
timestamp 1676557249
transform 1 0 43584 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _608_
timestamp 1676627187
transform 1 0 43872 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _609_
timestamp 1676557249
transform 1 0 43968 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _610_
timestamp 1676627187
transform 1 0 44256 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _611_
timestamp 1676557249
transform 1 0 44352 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _612_
timestamp 1676627187
transform 1 0 44640 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _613_
timestamp 1676557249
transform 1 0 44736 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _614_
timestamp 1676627187
transform 1 0 45024 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _615_
timestamp 1676557249
transform 1 0 45120 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _616_
timestamp 1676627187
transform 1 0 45408 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _617_
timestamp 1676557249
transform 1 0 45504 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _618_
timestamp 1676627187
transform 1 0 45792 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _619_
timestamp 1676557249
transform 1 0 45888 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _620_
timestamp 1676627187
transform 1 0 46176 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _621_
timestamp 1676557249
transform 1 0 46272 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _622_
timestamp 1676627187
transform 1 0 46560 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _623_
timestamp 1676557249
transform -1 0 47136 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _624_
timestamp 1676627187
transform 1 0 46944 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _625_
timestamp 1676557249
transform -1 0 47520 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _626_
timestamp 1676627187
transform 1 0 47328 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _627_
timestamp 1676557249
transform -1 0 47904 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _628_
timestamp 1676627187
transform 1 0 47712 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _629_
timestamp 1676557249
transform 1 0 47808 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _630_
timestamp 1676627187
transform 1 0 48096 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _631_
timestamp 1676557249
transform 1 0 48192 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _632_
timestamp 1676627187
transform 1 0 48480 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _633_
timestamp 1676557249
transform 1 0 48576 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _634_
timestamp 1676627187
transform 1 0 48864 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _635_
timestamp 1676557249
transform 1 0 48864 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _636_
timestamp 1676627187
transform -1 0 49632 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _637_
timestamp 1676557249
transform 1 0 49056 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _638_
timestamp 1676627187
transform -1 0 50976 0 -1 5292
box -48 -56 432 834
use sg13g2_or2_1  _639_
timestamp 1684236171
transform -1 0 50592 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _640_
timestamp 1676627187
transform 1 0 50016 0 -1 3780
box -48 -56 432 834
use sg13g2_or2_1  _641_
timestamp 1684236171
transform -1 0 50880 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _642_
timestamp 1676627187
transform 1 0 50304 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _643_
timestamp 1684236171
transform -1 0 51168 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _644_
timestamp 1676627187
transform 1 0 51168 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _645_
timestamp 1684236171
transform -1 0 51648 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _646_
timestamp 1676627187
transform -1 0 52416 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _647_
timestamp 1684236171
transform -1 0 52032 0 -1 2268
box -48 -56 528 834
use sg13g2_nor2_1  _648_
timestamp 1676627187
transform -1 0 52800 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _649_
timestamp 1684236171
transform -1 0 52416 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _650_
timestamp 1676627187
transform -1 0 52992 0 -1 5292
box -48 -56 432 834
use sg13g2_or2_1  _651_
timestamp 1684236171
transform -1 0 52608 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _652_
timestamp 1676627187
transform -1 0 53472 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _653_
timestamp 1684236171
transform -1 0 53088 0 -1 2268
box -48 -56 528 834
use sg13g2_nor2_1  _654_
timestamp 1676627187
transform -1 0 53952 0 1 3780
box -48 -56 432 834
use sg13g2_or2_1  _655_
timestamp 1684236171
transform -1 0 53568 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _656_
timestamp 1676627187
transform 1 0 53472 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _657_
timestamp 1684236171
transform -1 0 54336 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _658_
timestamp 1676627187
transform 1 0 54240 0 -1 2268
box -48 -56 432 834
use sg13g2_or2_1  _659_
timestamp 1684236171
transform -1 0 55296 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _660_
timestamp 1676627187
transform -1 0 55680 0 1 756
box -48 -56 432 834
use sg13g2_or2_1  _661_
timestamp 1684236171
transform -1 0 54816 0 1 756
box -48 -56 528 834
use sg13g2_nor2_1  _662_
timestamp 1676627187
transform -1 0 55488 0 -1 5292
box -48 -56 432 834
use sg13g2_or2_1  _663_
timestamp 1684236171
transform -1 0 55104 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _664_
timestamp 1676627187
transform 1 0 54624 0 1 2268
box -48 -56 432 834
use sg13g2_or2_1  _665_
timestamp 1684236171
transform -1 0 55488 0 1 2268
box -48 -56 528 834
use sg13g2_nor2_1  _666_
timestamp 1676627187
transform -1 0 56352 0 1 2268
box -48 -56 432 834
use sg13g2_or2_1  _667_
timestamp 1684236171
transform -1 0 55968 0 1 2268
box -48 -56 528 834
use sg13g2_nor2_1  _668_
timestamp 1676627187
transform -1 0 7296 0 1 3780
box -48 -56 432 834
use sg13g2_or2_1  _669_
timestamp 1684236171
transform -1 0 7776 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _670_
timestamp 1676627187
transform -1 0 1344 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _671_
timestamp 1676557249
transform -1 0 1824 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _672_
timestamp 1676627187
transform -1 0 1728 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _673_
timestamp 1676557249
transform -1 0 1920 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _674_
timestamp 1676627187
transform -1 0 2112 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _675_
timestamp 1676557249
transform 1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _676_
timestamp 1676627187
transform -1 0 2496 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _677_
timestamp 1676557249
transform 1 0 2016 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _678_
timestamp 1676627187
transform -1 0 2880 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _679_
timestamp 1676557249
transform 1 0 2400 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _680_
timestamp 1676627187
transform -1 0 3264 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _681_
timestamp 1676557249
transform 1 0 2880 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _682_
timestamp 1676627187
transform -1 0 3648 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _683_
timestamp 1676557249
transform 1 0 3264 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _684_
timestamp 1676627187
transform -1 0 4032 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _685_
timestamp 1676557249
transform 1 0 3648 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _686_
timestamp 1676627187
transform -1 0 4416 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _687_
timestamp 1676557249
transform 1 0 4128 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _688_
timestamp 1676627187
transform -1 0 4800 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _689_
timestamp 1676557249
transform 1 0 4512 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _690_
timestamp 1676627187
transform -1 0 5184 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _691_
timestamp 1676557249
transform 1 0 4896 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _692_
timestamp 1676627187
transform -1 0 5568 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _693_
timestamp 1676557249
transform 1 0 5280 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _694_
timestamp 1676627187
transform -1 0 5952 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _695_
timestamp 1676557249
transform 1 0 5664 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _696_
timestamp 1676627187
transform -1 0 6336 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _697_
timestamp 1676557249
transform 1 0 6048 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _698_
timestamp 1676627187
transform -1 0 7104 0 -1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _699_
timestamp 1676557249
transform 1 0 6528 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _700_
timestamp 1676627187
transform -1 0 6720 0 1 756
box -48 -56 432 834
use sg13g2_nand2_1  _701_
timestamp 1676557249
transform 1 0 6912 0 1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_0_0
timestamp 1679577901
transform 1 0 576 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_256
timestamp 1677580104
transform 1 0 25152 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_258
timestamp 1677579658
transform 1 0 25344 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_319
timestamp 1677580104
transform 1 0 31200 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_381
timestamp 1677579658
transform 1 0 37152 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_446
timestamp 1677579658
transform 1 0 43392 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_532
timestamp 1677580104
transform 1 0 51648 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_534
timestamp 1677579658
transform 1 0 51840 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_544
timestamp 1679581782
transform 1 0 52800 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_574
timestamp 1679577901
transform 1 0 55680 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_578
timestamp 1677579658
transform 1 0 56064 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_593
timestamp 1677579658
transform 1 0 57504 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_603
timestamp 1679577901
transform 1 0 58464 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_607
timestamp 1677580104
transform 1 0 58848 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_632
timestamp 1679581782
transform 1 0 61248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_639
timestamp 1679581782
transform 1 0 61920 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_834
timestamp 1677580104
transform 1 0 80640 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_1028
timestamp 1677579658
transform 1 0 99264 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_7
timestamp 1677580104
transform 1 0 1248 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_13
timestamp 1679581782
transform 1 0 1824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_20
timestamp 1679581782
transform 1 0 2496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_27
timestamp 1679581782
transform 1 0 3168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_34
timestamp 1679581782
transform 1 0 3840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_41
timestamp 1679581782
transform 1 0 4512 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_48
timestamp 1677579658
transform 1 0 5184 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_53
timestamp 1679581782
transform 1 0 5664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_60
timestamp 1679577901
transform 1 0 6336 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_68
timestamp 1679581782
transform 1 0 7104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_75
timestamp 1679581782
transform 1 0 7776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_82
timestamp 1679581782
transform 1 0 8448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_89
timestamp 1679581782
transform 1 0 9120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_96
timestamp 1679581782
transform 1 0 9792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_103
timestamp 1679581782
transform 1 0 10464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_110
timestamp 1679581782
transform 1 0 11136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_117
timestamp 1679581782
transform 1 0 11808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_124
timestamp 1679581782
transform 1 0 12480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_131
timestamp 1679581782
transform 1 0 13152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_138
timestamp 1679581782
transform 1 0 13824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_145
timestamp 1679581782
transform 1 0 14496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_152
timestamp 1679581782
transform 1 0 15168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_159
timestamp 1679581782
transform 1 0 15840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_166
timestamp 1679581782
transform 1 0 16512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_173
timestamp 1679581782
transform 1 0 17184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_180
timestamp 1679581782
transform 1 0 17856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_187
timestamp 1679581782
transform 1 0 18528 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_194
timestamp 1677579658
transform 1 0 19200 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_199
timestamp 1679581782
transform 1 0 19680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_206
timestamp 1679581782
transform 1 0 20352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_213
timestamp 1679581782
transform 1 0 21024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_220
timestamp 1679581782
transform 1 0 21696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_227
timestamp 1679581782
transform 1 0 22368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_234
timestamp 1679581782
transform 1 0 23040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_241
timestamp 1679581782
transform 1 0 23712 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_248
timestamp 1677580104
transform 1 0 24384 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_254
timestamp 1679581782
transform 1 0 24960 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_261
timestamp 1677580104
transform 1 0 25632 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_267
timestamp 1679581782
transform 1 0 26208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_274
timestamp 1679581782
transform 1 0 26880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_281
timestamp 1679581782
transform 1 0 27552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_288
timestamp 1679581782
transform 1 0 28224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_295
timestamp 1679581782
transform 1 0 28896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_302
timestamp 1679581782
transform 1 0 29568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_309
timestamp 1679581782
transform 1 0 30240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_316
timestamp 1679581782
transform 1 0 30912 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_323
timestamp 1677580104
transform 1 0 31584 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_325
timestamp 1677579658
transform 1 0 31776 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_330
timestamp 1679581782
transform 1 0 32256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_337
timestamp 1679581782
transform 1 0 32928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_344
timestamp 1679581782
transform 1 0 33600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_351
timestamp 1679581782
transform 1 0 34272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_358
timestamp 1679581782
transform 1 0 34944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_365
timestamp 1679581782
transform 1 0 35616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_372
timestamp 1679581782
transform 1 0 36288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_379
timestamp 1679581782
transform 1 0 36960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_386
timestamp 1679581782
transform 1 0 37632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_393
timestamp 1679581782
transform 1 0 38304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_400
timestamp 1679581782
transform 1 0 38976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_407
timestamp 1679581782
transform 1 0 39648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_414
timestamp 1679581782
transform 1 0 40320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_421
timestamp 1679581782
transform 1 0 40992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_428
timestamp 1679581782
transform 1 0 41664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_435
timestamp 1679581782
transform 1 0 42336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_442
timestamp 1679577901
transform 1 0 43008 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_446
timestamp 1677580104
transform 1 0 43392 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_452
timestamp 1679581782
transform 1 0 43968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_459
timestamp 1679581782
transform 1 0 44640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_466
timestamp 1679581782
transform 1 0 45312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_473
timestamp 1679581782
transform 1 0 45984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_480
timestamp 1679581782
transform 1 0 46656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_487
timestamp 1679581782
transform 1 0 47328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_494
timestamp 1679581782
transform 1 0 48000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_501
timestamp 1679581782
transform 1 0 48672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_508
timestamp 1679581782
transform 1 0 49344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_515
timestamp 1679581782
transform 1 0 50016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_522
timestamp 1679577901
transform 1 0 50688 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_526
timestamp 1677579658
transform 1 0 51072 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_540
timestamp 1677580104
transform 1 0 52416 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_551
timestamp 1679581782
transform 1 0 53472 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_558
timestamp 1677579658
transform 1 0 54144 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_563
timestamp 1679581782
transform 1 0 54624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_570
timestamp 1679581782
transform 1 0 55296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_577
timestamp 1679581782
transform 1 0 55968 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_584
timestamp 1677580104
transform 1 0 56640 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_586
timestamp 1677579658
transform 1 0 56832 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_600
timestamp 1679577901
transform 1 0 58176 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_604
timestamp 1677579658
transform 1 0 58560 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_616
timestamp 1677580104
transform 1 0 59712 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_622
timestamp 1679581782
transform 1 0 60288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_629
timestamp 1679581782
transform 1 0 60960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_636
timestamp 1679581782
transform 1 0 61632 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_643
timestamp 1677580104
transform 1 0 62304 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_649
timestamp 1679581782
transform 1 0 62880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_656
timestamp 1679581782
transform 1 0 63552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_663
timestamp 1679577901
transform 1 0 64224 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_667
timestamp 1677580104
transform 1 0 64608 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_673
timestamp 1679581782
transform 1 0 65184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_680
timestamp 1679577901
transform 1 0 65856 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_684
timestamp 1677579658
transform 1 0 66240 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_689
timestamp 1679581782
transform 1 0 66720 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_696
timestamp 1677580104
transform 1 0 67392 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_702
timestamp 1679581782
transform 1 0 67968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_709
timestamp 1679581782
transform 1 0 68640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_716
timestamp 1679581782
transform 1 0 69312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_723
timestamp 1679581782
transform 1 0 69984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_730
timestamp 1679581782
transform 1 0 70656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_737
timestamp 1679581782
transform 1 0 71328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_744
timestamp 1679581782
transform 1 0 72000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_751
timestamp 1679581782
transform 1 0 72672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_758
timestamp 1679581782
transform 1 0 73344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_765
timestamp 1679581782
transform 1 0 74016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_772
timestamp 1679581782
transform 1 0 74688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_779
timestamp 1679581782
transform 1 0 75360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_786
timestamp 1679581782
transform 1 0 76032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_793
timestamp 1679581782
transform 1 0 76704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_800
timestamp 1679581782
transform 1 0 77376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_807
timestamp 1679581782
transform 1 0 78048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_814
timestamp 1679581782
transform 1 0 78720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_821
timestamp 1679577901
transform 1 0 79392 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_825
timestamp 1677579658
transform 1 0 79776 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_830
timestamp 1679577901
transform 1 0 80256 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_834
timestamp 1677579658
transform 1 0 80640 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_839
timestamp 1679581782
transform 1 0 81120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_846
timestamp 1679581782
transform 1 0 81792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_853
timestamp 1679581782
transform 1 0 82464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_860
timestamp 1679581782
transform 1 0 83136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_867
timestamp 1679581782
transform 1 0 83808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_874
timestamp 1679581782
transform 1 0 84480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_881
timestamp 1679581782
transform 1 0 85152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_888
timestamp 1679581782
transform 1 0 85824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_895
timestamp 1679581782
transform 1 0 86496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_902
timestamp 1679581782
transform 1 0 87168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_909
timestamp 1679581782
transform 1 0 87840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_916
timestamp 1679581782
transform 1 0 88512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_923
timestamp 1679581782
transform 1 0 89184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_930
timestamp 1679581782
transform 1 0 89856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_937
timestamp 1679581782
transform 1 0 90528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_944
timestamp 1679581782
transform 1 0 91200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_951
timestamp 1679577901
transform 1 0 91872 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_955
timestamp 1677580104
transform 1 0 92256 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_961
timestamp 1679581782
transform 1 0 92832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_968
timestamp 1679581782
transform 1 0 93504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_975
timestamp 1679581782
transform 1 0 94176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_982
timestamp 1679581782
transform 1 0 94848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_989
timestamp 1679581782
transform 1 0 95520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_996
timestamp 1679581782
transform 1 0 96192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1003
timestamp 1679581782
transform 1 0 96864 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_1010
timestamp 1677580104
transform 1 0 97536 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_1012
timestamp 1677579658
transform 1 0 97728 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_1017
timestamp 1679581782
transform 1 0 98208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_1024
timestamp 1679577901
transform 1 0 98880 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_1028
timestamp 1677579658
transform 1 0 99264 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 576 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_7
timestamp 1677580104
transform 1 0 1248 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_9
timestamp 1677579658
transform 1 0 1440 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_14
timestamp 1677579658
transform 1 0 1920 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_23
timestamp 1677579658
transform 1 0 2784 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_36
timestamp 1679581782
transform 1 0 4032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_43
timestamp 1679581782
transform 1 0 4704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_50
timestamp 1679581782
transform 1 0 5376 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_61
timestamp 1677579658
transform 1 0 6432 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_123
timestamp 1677579658
transform 1 0 12384 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_128
timestamp 1679581782
transform 1 0 12864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_135
timestamp 1679577901
transform 1 0 13536 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_139
timestamp 1677579658
transform 1 0 13920 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_193
timestamp 1679577901
transform 1 0 19104 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_197
timestamp 1677579658
transform 1 0 19488 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_202
timestamp 1677580104
transform 1 0 19968 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_208
timestamp 1679581782
transform 1 0 20544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_215
timestamp 1679577901
transform 1 0 21216 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_219
timestamp 1677580104
transform 1 0 21600 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_225
timestamp 1679581782
transform 1 0 22176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_232
timestamp 1679577901
transform 1 0 22848 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_236
timestamp 1677579658
transform 1 0 23232 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_241
timestamp 1679581782
transform 1 0 23712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_248
timestamp 1679581782
transform 1 0 24384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_255
timestamp 1679581782
transform 1 0 25056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_262
timestamp 1679577901
transform 1 0 25728 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_266
timestamp 1677580104
transform 1 0 26112 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_272
timestamp 1679581782
transform 1 0 26688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_279
timestamp 1679577901
transform 1 0 27360 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_283
timestamp 1677579658
transform 1 0 27744 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_288
timestamp 1679581782
transform 1 0 28224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_295
timestamp 1679577901
transform 1 0 28896 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_299
timestamp 1677580104
transform 1 0 29280 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_312
timestamp 1677579658
transform 1 0 30528 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_317
timestamp 1679577901
transform 1 0 31008 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_321
timestamp 1677580104
transform 1 0 31392 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_327
timestamp 1679581782
transform 1 0 31968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_334
timestamp 1679581782
transform 1 0 32640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_341
timestamp 1679581782
transform 1 0 33312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_348
timestamp 1679581782
transform 1 0 33984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_355
timestamp 1679581782
transform 1 0 34656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_362
timestamp 1679581782
transform 1 0 35328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_369
timestamp 1679581782
transform 1 0 36000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_376
timestamp 1679581782
transform 1 0 36672 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_383
timestamp 1677580104
transform 1 0 37344 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_389
timestamp 1677580104
transform 1 0 37920 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_399
timestamp 1679581782
transform 1 0 38880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_406
timestamp 1679577901
transform 1 0 39552 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_414
timestamp 1679581782
transform 1 0 40320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_421
timestamp 1679577901
transform 1 0 40992 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_425
timestamp 1677580104
transform 1 0 41376 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_435
timestamp 1679577901
transform 1 0 42336 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_443
timestamp 1679581782
transform 1 0 43104 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_450
timestamp 1677580104
transform 1 0 43776 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_456
timestamp 1679577901
transform 1 0 44352 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_464
timestamp 1679581782
transform 1 0 45120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_471
timestamp 1679577901
transform 1 0 45792 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_475
timestamp 1677579658
transform 1 0 46176 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_487
timestamp 1679577901
transform 1 0 47328 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_491
timestamp 1677579658
transform 1 0 47712 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_504
timestamp 1677579658
transform 1 0 48960 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_509
timestamp 1679581782
transform 1 0 49440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_516
timestamp 1679581782
transform 1 0 50112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_523
timestamp 1679581782
transform 1 0 50784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_530
timestamp 1679581782
transform 1 0 51456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_537
timestamp 1679581782
transform 1 0 52128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_544
timestamp 1679581782
transform 1 0 52800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_551
timestamp 1679581782
transform 1 0 53472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_558
timestamp 1679577901
transform 1 0 54144 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_562
timestamp 1677579658
transform 1 0 54528 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_581
timestamp 1679581782
transform 1 0 56352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_588
timestamp 1679581782
transform 1 0 57024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_595
timestamp 1679581782
transform 1 0 57696 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_602
timestamp 1677579658
transform 1 0 58368 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_608
timestamp 1679581782
transform 1 0 58944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_615
timestamp 1679581782
transform 1 0 59616 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_622
timestamp 1677579658
transform 1 0 60288 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_652
timestamp 1677579658
transform 1 0 63168 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_657
timestamp 1679581782
transform 1 0 63648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_664
timestamp 1679581782
transform 1 0 64320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_671
timestamp 1679581782
transform 1 0 64992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_678
timestamp 1679581782
transform 1 0 65664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_685
timestamp 1679581782
transform 1 0 66336 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_692
timestamp 1677580104
transform 1 0 67008 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_694
timestamp 1677579658
transform 1 0 67200 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_699
timestamp 1679581782
transform 1 0 67680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_706
timestamp 1679581782
transform 1 0 68352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_713
timestamp 1679581782
transform 1 0 69024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_720
timestamp 1679581782
transform 1 0 69696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_727
timestamp 1679581782
transform 1 0 70368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_734
timestamp 1679581782
transform 1 0 71040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_741
timestamp 1679581782
transform 1 0 71712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_748
timestamp 1679577901
transform 1 0 72384 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_752
timestamp 1677579658
transform 1 0 72768 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_769
timestamp 1677580104
transform 1 0 74400 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_771
timestamp 1677579658
transform 1 0 74592 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_776
timestamp 1679577901
transform 1 0 75072 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_780
timestamp 1677579658
transform 1 0 75456 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_785
timestamp 1679581782
transform 1 0 75936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_792
timestamp 1679577901
transform 1 0 76608 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_800
timestamp 1679581782
transform 1 0 77376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_807
timestamp 1679577901
transform 1 0 78048 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_811
timestamp 1677579658
transform 1 0 78432 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_848
timestamp 1679581782
transform 1 0 81984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_855
timestamp 1679577901
transform 1 0 82656 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_859
timestamp 1677579658
transform 1 0 83040 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_864
timestamp 1679581782
transform 1 0 83520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_871
timestamp 1679577901
transform 1 0 84192 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_875
timestamp 1677579658
transform 1 0 84576 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_896
timestamp 1679581782
transform 1 0 86592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_903
timestamp 1679581782
transform 1 0 87264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_910
timestamp 1679581782
transform 1 0 87936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_917
timestamp 1679581782
transform 1 0 88608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_924
timestamp 1679581782
transform 1 0 89280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_931
timestamp 1679581782
transform 1 0 89952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_938
timestamp 1679581782
transform 1 0 90624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_945
timestamp 1679581782
transform 1 0 91296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_952
timestamp 1679581782
transform 1 0 91968 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_959
timestamp 1677580104
transform 1 0 92640 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_965
timestamp 1677580104
transform 1 0 93216 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_967
timestamp 1677579658
transform 1 0 93408 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_972
timestamp 1679581782
transform 1 0 93888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_979
timestamp 1679577901
transform 1 0 94560 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_983
timestamp 1677579658
transform 1 0 94944 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_988
timestamp 1679581782
transform 1 0 95424 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_995
timestamp 1677580104
transform 1 0 96096 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_1017
timestamp 1679581782
transform 1 0 98208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_1024
timestamp 1679577901
transform 1 0 98880 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_7
timestamp 1679577901
transform 1 0 1248 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_11
timestamp 1677580104
transform 1 0 1632 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_17
timestamp 1679581782
transform 1 0 2208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_24
timestamp 1679581782
transform 1 0 2880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_31
timestamp 1679577901
transform 1 0 3552 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_35
timestamp 1677580104
transform 1 0 3936 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_49
timestamp 1679577901
transform 1 0 5280 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_57
timestamp 1679581782
transform 1 0 6048 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_64
timestamp 1677579658
transform 1 0 6720 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_77
timestamp 1679577901
transform 1 0 7968 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_3_125
timestamp 1679577901
transform 1 0 12576 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_141
timestamp 1677579658
transform 1 0 14112 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_195
timestamp 1679577901
transform 1 0 19296 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_199
timestamp 1677580104
transform 1 0 19680 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_205
timestamp 1679577901
transform 1 0 20256 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_221
timestamp 1677580104
transform 1 0 21792 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_223
timestamp 1677579658
transform 1 0 21984 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_236
timestamp 1677580104
transform 1 0 23232 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_238
timestamp 1677579658
transform 1 0 23424 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_251
timestamp 1679577901
transform 1 0 24672 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_255
timestamp 1677580104
transform 1 0 25056 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_269
timestamp 1677580104
transform 1 0 26400 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_271
timestamp 1677579658
transform 1 0 26592 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_280
timestamp 1677579658
transform 1 0 27456 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_285
timestamp 1679577901
transform 1 0 27936 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_301
timestamp 1677579658
transform 1 0 29472 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_314
timestamp 1679577901
transform 1 0 30720 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_318
timestamp 1677579658
transform 1 0 31104 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_379
timestamp 1679581782
transform 1 0 36960 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_386
timestamp 1677579658
transform 1 0 37632 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_396
timestamp 1677580104
transform 1 0 38592 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_410
timestamp 1677580104
transform 1 0 39936 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_412
timestamp 1677579658
transform 1 0 40128 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_417
timestamp 1677579658
transform 1 0 40608 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_426
timestamp 1679577901
transform 1 0 41472 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_443
timestamp 1679581782
transform 1 0 43104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_450
timestamp 1679577901
transform 1 0 43776 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_454
timestamp 1677580104
transform 1 0 44160 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_460
timestamp 1679577901
transform 1 0 44736 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_3_476
timestamp 1679577901
transform 1 0 46272 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_480
timestamp 1677579658
transform 1 0 46656 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_493
timestamp 1679581782
transform 1 0 47904 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_500
timestamp 1677580104
transform 1 0 48576 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_502
timestamp 1677579658
transform 1 0 48768 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_507
timestamp 1679581782
transform 1 0 49248 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_514
timestamp 1677579658
transform 1 0 49920 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_528
timestamp 1679581782
transform 1 0 51264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_535
timestamp 1679577901
transform 1 0 51936 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_539
timestamp 1677580104
transform 1 0 52320 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_545
timestamp 1677580104
transform 1 0 52896 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_547
timestamp 1677579658
transform 1 0 53088 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_552
timestamp 1679581782
transform 1 0 53568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_559
timestamp 1679577901
transform 1 0 54240 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_563
timestamp 1677580104
transform 1 0 54624 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_573
timestamp 1679581782
transform 1 0 55584 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_580
timestamp 1677579658
transform 1 0 56256 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_590
timestamp 1679581782
transform 1 0 57216 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_597
timestamp 1677580104
transform 1 0 57888 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_634
timestamp 1677579658
transform 1 0 61440 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_639
timestamp 1679581782
transform 1 0 61920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_646
timestamp 1679577901
transform 1 0 62592 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_650
timestamp 1677579658
transform 1 0 62976 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_655
timestamp 1677580104
transform 1 0 63456 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_657
timestamp 1677579658
transform 1 0 63648 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_670
timestamp 1677580104
transform 1 0 64896 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_672
timestamp 1677579658
transform 1 0 65088 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_685
timestamp 1679577901
transform 1 0 66336 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_704
timestamp 1679577901
transform 1 0 68160 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_756
timestamp 1679581782
transform 1 0 73152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_763
timestamp 1679581782
transform 1 0 73824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_770
timestamp 1679577901
transform 1 0 74496 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_782
timestamp 1677580104
transform 1 0 75648 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_784
timestamp 1677579658
transform 1 0 75840 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_797
timestamp 1677580104
transform 1 0 77088 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_799
timestamp 1677579658
transform 1 0 77280 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_804
timestamp 1677579658
transform 1 0 77760 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_813
timestamp 1677580104
transform 1 0 78624 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_815
timestamp 1677579658
transform 1 0 78816 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_832
timestamp 1679577901
transform 1 0 80448 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_836
timestamp 1677580104
transform 1 0 80832 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_846
timestamp 1677580104
transform 1 0 81792 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_848
timestamp 1677579658
transform 1 0 81984 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_861
timestamp 1677580104
transform 1 0 83232 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_863
timestamp 1677579658
transform 1 0 83424 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_876
timestamp 1679581782
transform 1 0 84672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_883
timestamp 1679581782
transform 1 0 85344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_890
timestamp 1679581782
transform 1 0 86016 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_897
timestamp 1677579658
transform 1 0 86688 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_962
timestamp 1677580104
transform 1 0 92928 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_964
timestamp 1677579658
transform 1 0 93120 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_969
timestamp 1679577901
transform 1 0 93600 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_985
timestamp 1677580104
transform 1 0 95136 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_987
timestamp 1677579658
transform 1 0 95328 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_992
timestamp 1677579658
transform 1 0 95808 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_997
timestamp 1679581782
transform 1 0 96288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1004
timestamp 1679581782
transform 1 0 96960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1011
timestamp 1679581782
transform 1 0 97632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1018
timestamp 1679581782
transform 1 0 98304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_1025
timestamp 1679577901
transform 1 0 98976 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 1920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 2592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 3936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 4608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 5952 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_63
timestamp 1677580104
transform 1 0 6624 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_65
timestamp 1677579658
transform 1 0 6816 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_75
timestamp 1679581782
transform 1 0 7776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_82
timestamp 1679581782
transform 1 0 8448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_89
timestamp 1679581782
transform 1 0 9120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_96
timestamp 1679581782
transform 1 0 9792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_103
timestamp 1679581782
transform 1 0 10464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_110
timestamp 1679581782
transform 1 0 11136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_117
timestamp 1679581782
transform 1 0 11808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_124
timestamp 1679581782
transform 1 0 12480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_131
timestamp 1679581782
transform 1 0 13152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_138
timestamp 1679581782
transform 1 0 13824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_145
timestamp 1679581782
transform 1 0 14496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_152
timestamp 1679581782
transform 1 0 15168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_159
timestamp 1679581782
transform 1 0 15840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_166
timestamp 1679581782
transform 1 0 16512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_173
timestamp 1679581782
transform 1 0 17184 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_180
timestamp 1677580104
transform 1 0 17856 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_201
timestamp 1679581782
transform 1 0 19872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_208
timestamp 1679581782
transform 1 0 20544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_215
timestamp 1679581782
transform 1 0 21216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_222
timestamp 1679581782
transform 1 0 21888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_229
timestamp 1679581782
transform 1 0 22560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_236
timestamp 1679581782
transform 1 0 23232 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_243
timestamp 1677580104
transform 1 0 23904 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_257
timestamp 1679577901
transform 1 0 25248 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_261
timestamp 1677580104
transform 1 0 25632 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_267
timestamp 1679581782
transform 1 0 26208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_274
timestamp 1679581782
transform 1 0 26880 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_281
timestamp 1677579658
transform 1 0 27552 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679581782
transform 1 0 28128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679581782
transform 1 0 28800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679581782
transform 1 0 29472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_308
timestamp 1679581782
transform 1 0 30144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_315
timestamp 1679581782
transform 1 0 30816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_322
timestamp 1679577901
transform 1 0 31488 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_338
timestamp 1679581782
transform 1 0 33024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_345
timestamp 1679581782
transform 1 0 33696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_352
timestamp 1679581782
transform 1 0 34368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_359
timestamp 1679581782
transform 1 0 35040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_366
timestamp 1679581782
transform 1 0 35712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_373
timestamp 1679577901
transform 1 0 36384 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_377
timestamp 1677580104
transform 1 0 36768 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_398
timestamp 1679581782
transform 1 0 38784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_405
timestamp 1679581782
transform 1 0 39456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_412
timestamp 1679581782
transform 1 0 40128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_419
timestamp 1679577901
transform 1 0 40800 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_445
timestamp 1679581782
transform 1 0 43296 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_452
timestamp 1677580104
transform 1 0 43968 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_454
timestamp 1677579658
transform 1 0 44160 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_465
timestamp 1679581782
transform 1 0 45216 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_472
timestamp 1677579658
transform 1 0 45888 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_478
timestamp 1679581782
transform 1 0 46464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_485
timestamp 1679581782
transform 1 0 47136 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_492
timestamp 1677580104
transform 1 0 47808 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_494
timestamp 1677579658
transform 1 0 48000 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_505
timestamp 1679581782
transform 1 0 49056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_512
timestamp 1679577901
transform 1 0 49728 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_524
timestamp 1677580104
transform 1 0 50880 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_526
timestamp 1677579658
transform 1 0 51072 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_532
timestamp 1679577901
transform 1 0 51648 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_536
timestamp 1677579658
transform 1 0 52032 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_545
timestamp 1677580104
transform 1 0 52896 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_556
timestamp 1679581782
transform 1 0 53952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_563
timestamp 1679577901
transform 1 0 54624 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_572
timestamp 1679581782
transform 1 0 55488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_579
timestamp 1679581782
transform 1 0 56160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_586
timestamp 1679581782
transform 1 0 56832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_593
timestamp 1679577901
transform 1 0 57504 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_597
timestamp 1677579658
transform 1 0 57888 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_616
timestamp 1679581782
transform 1 0 59712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_623
timestamp 1679581782
transform 1 0 60384 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_630
timestamp 1677580104
transform 1 0 61056 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_646
timestamp 1679581782
transform 1 0 62592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_653
timestamp 1679581782
transform 1 0 63264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_660
timestamp 1679581782
transform 1 0 63936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_667
timestamp 1679581782
transform 1 0 64608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_674
timestamp 1679581782
transform 1 0 65280 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_681
timestamp 1677580104
transform 1 0 65952 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_683
timestamp 1677579658
transform 1 0 66144 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_693
timestamp 1679581782
transform 1 0 67104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_700
timestamp 1679577901
transform 1 0 67776 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_704
timestamp 1677580104
transform 1 0 68160 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_715
timestamp 1679581782
transform 1 0 69216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_722
timestamp 1679581782
transform 1 0 69888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_729
timestamp 1679581782
transform 1 0 70560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_736
timestamp 1679581782
transform 1 0 71232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_743
timestamp 1679581782
transform 1 0 71904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_750
timestamp 1679581782
transform 1 0 72576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_757
timestamp 1679581782
transform 1 0 73248 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_764
timestamp 1677579658
transform 1 0 73920 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_777
timestamp 1679581782
transform 1 0 75168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_784
timestamp 1679581782
transform 1 0 75840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_791
timestamp 1679581782
transform 1 0 76512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_798
timestamp 1679581782
transform 1 0 77184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_805
timestamp 1679581782
transform 1 0 77856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_812
timestamp 1679581782
transform 1 0 78528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_819
timestamp 1679581782
transform 1 0 79200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_826
timestamp 1679577901
transform 1 0 79872 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_839
timestamp 1679581782
transform 1 0 81120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_846
timestamp 1679581782
transform 1 0 81792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_853
timestamp 1679581782
transform 1 0 82464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_860
timestamp 1679581782
transform 1 0 83136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_867
timestamp 1679581782
transform 1 0 83808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_874
timestamp 1679581782
transform 1 0 84480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_881
timestamp 1679581782
transform 1 0 85152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_888
timestamp 1679581782
transform 1 0 85824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_904
timestamp 1679581782
transform 1 0 87360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_911
timestamp 1679581782
transform 1 0 88032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_918
timestamp 1679581782
transform 1 0 88704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_925
timestamp 1679581782
transform 1 0 89376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_932
timestamp 1679581782
transform 1 0 90048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_939
timestamp 1679581782
transform 1 0 90720 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_946
timestamp 1677579658
transform 1 0 91392 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_956
timestamp 1679581782
transform 1 0 92352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_963
timestamp 1679581782
transform 1 0 93024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_970
timestamp 1679581782
transform 1 0 93696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_977
timestamp 1679581782
transform 1 0 94368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_984
timestamp 1679581782
transform 1 0 95040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_991
timestamp 1679581782
transform 1 0 95712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_998
timestamp 1679581782
transform 1 0 96384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1005
timestamp 1679581782
transform 1 0 97056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1012
timestamp 1679581782
transform 1 0 97728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1019
timestamp 1679581782
transform 1 0 98400 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_1026
timestamp 1677580104
transform 1 0 99072 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_1028
timestamp 1677579658
transform 1 0 99264 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 1920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 2592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 3936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 4608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 5952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 6624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 7968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679581782
transform 1 0 8640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679581782
transform 1 0 9312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679581782
transform 1 0 9984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 10656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679581782
transform 1 0 11328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 12000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679581782
transform 1 0 12672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679581782
transform 1 0 13344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679581782
transform 1 0 14016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 14688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 16704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679581782
transform 1 0 17376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679581782
transform 1 0 18048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679581782
transform 1 0 18720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679581782
transform 1 0 19392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679581782
transform 1 0 20064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 20736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679581782
transform 1 0 21408 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_224
timestamp 1677580104
transform 1 0 22080 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_229
timestamp 1679581782
transform 1 0 22560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_236
timestamp 1679581782
transform 1 0 23232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_243
timestamp 1679581782
transform 1 0 23904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_250
timestamp 1679581782
transform 1 0 24576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_257
timestamp 1679581782
transform 1 0 25248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_264
timestamp 1679581782
transform 1 0 25920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_271
timestamp 1679581782
transform 1 0 26592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_278
timestamp 1679581782
transform 1 0 27264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_285
timestamp 1679581782
transform 1 0 27936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_292
timestamp 1679581782
transform 1 0 28608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_299
timestamp 1679581782
transform 1 0 29280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_306
timestamp 1679581782
transform 1 0 29952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_313
timestamp 1679581782
transform 1 0 30624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_320
timestamp 1679581782
transform 1 0 31296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_327
timestamp 1679581782
transform 1 0 31968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_334
timestamp 1679581782
transform 1 0 32640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_341
timestamp 1679581782
transform 1 0 33312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_348
timestamp 1679581782
transform 1 0 33984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_355
timestamp 1679581782
transform 1 0 34656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_362
timestamp 1679581782
transform 1 0 35328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_369
timestamp 1679581782
transform 1 0 36000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_376
timestamp 1679581782
transform 1 0 36672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_383
timestamp 1679581782
transform 1 0 37344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_390
timestamp 1679581782
transform 1 0 38016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_397
timestamp 1679581782
transform 1 0 38688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_404
timestamp 1679581782
transform 1 0 39360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_411
timestamp 1679581782
transform 1 0 40032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_418
timestamp 1679577901
transform 1 0 40704 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_436
timestamp 1679581782
transform 1 0 42432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_443
timestamp 1679581782
transform 1 0 43104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_450
timestamp 1679581782
transform 1 0 43776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_457
timestamp 1679581782
transform 1 0 44448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_464
timestamp 1679577901
transform 1 0 45120 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_468
timestamp 1677579658
transform 1 0 45504 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_483
timestamp 1679581782
transform 1 0 46944 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_490
timestamp 1677580104
transform 1 0 47616 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_506
timestamp 1677579658
transform 1 0 49152 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_512
timestamp 1679577901
transform 1 0 49728 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_525
timestamp 1679581782
transform 1 0 50976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_532
timestamp 1679577901
transform 1 0 51648 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_536
timestamp 1677579658
transform 1 0 52032 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_546
timestamp 1679577901
transform 1 0 52992 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_550
timestamp 1677579658
transform 1 0 53376 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_555
timestamp 1679581782
transform 1 0 53856 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_562
timestamp 1677579658
transform 1 0 54528 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_572
timestamp 1679577901
transform 1 0 55488 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_592
timestamp 1677580104
transform 1 0 57408 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_594
timestamp 1677579658
transform 1 0 57600 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_609
timestamp 1679581782
transform 1 0 59040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_616
timestamp 1679577901
transform 1 0 59712 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_620
timestamp 1677580104
transform 1 0 60096 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_695
timestamp 1679581782
transform 1 0 67296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_702
timestamp 1679581782
transform 1 0 67968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_709
timestamp 1679581782
transform 1 0 68640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_716
timestamp 1679581782
transform 1 0 69312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_723
timestamp 1679581782
transform 1 0 69984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_730
timestamp 1679581782
transform 1 0 70656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_737
timestamp 1679581782
transform 1 0 71328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_744
timestamp 1679581782
transform 1 0 72000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_751
timestamp 1679577901
transform 1 0 72672 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_755
timestamp 1677580104
transform 1 0 73056 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_771
timestamp 1679581782
transform 1 0 74592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_778
timestamp 1679581782
transform 1 0 75264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_785
timestamp 1679581782
transform 1 0 75936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_792
timestamp 1679581782
transform 1 0 76608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_799
timestamp 1679581782
transform 1 0 77280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_806
timestamp 1679581782
transform 1 0 77952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_813
timestamp 1679581782
transform 1 0 78624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_820
timestamp 1679581782
transform 1 0 79296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_827
timestamp 1679581782
transform 1 0 79968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_834
timestamp 1679581782
transform 1 0 80640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_841
timestamp 1679581782
transform 1 0 81312 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_848
timestamp 1677579658
transform 1 0 81984 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_853
timestamp 1679581782
transform 1 0 82464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_860
timestamp 1679581782
transform 1 0 83136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_867
timestamp 1679581782
transform 1 0 83808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_874
timestamp 1679581782
transform 1 0 84480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_881
timestamp 1679581782
transform 1 0 85152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_888
timestamp 1679581782
transform 1 0 85824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_895
timestamp 1679581782
transform 1 0 86496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_902
timestamp 1679581782
transform 1 0 87168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_909
timestamp 1679581782
transform 1 0 87840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_916
timestamp 1679581782
transform 1 0 88512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_923
timestamp 1679581782
transform 1 0 89184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_930
timestamp 1679581782
transform 1 0 89856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_937
timestamp 1679581782
transform 1 0 90528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_944
timestamp 1679581782
transform 1 0 91200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_951
timestamp 1679581782
transform 1 0 91872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_958
timestamp 1679581782
transform 1 0 92544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_965
timestamp 1679581782
transform 1 0 93216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_972
timestamp 1679581782
transform 1 0 93888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_979
timestamp 1679581782
transform 1 0 94560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_986
timestamp 1679581782
transform 1 0 95232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_993
timestamp 1679581782
transform 1 0 95904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1000
timestamp 1679581782
transform 1 0 96576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1007
timestamp 1679581782
transform 1 0 97248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1014
timestamp 1679581782
transform 1 0 97920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1021
timestamp 1679581782
transform 1 0 98592 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_1028
timestamp 1677579658
transform 1 0 99264 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 1920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 2592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 3936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 4608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 5952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 6624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 7968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 8640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 9984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 10656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 12672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 14688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 16704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 18720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 20736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679581782
transform 1 0 22080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679581782
transform 1 0 22752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679581782
transform 1 0 23424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679581782
transform 1 0 24096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679581782
transform 1 0 24768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 25440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679581782
transform 1 0 26112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679581782
transform 1 0 26784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1679581782
transform 1 0 27456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1679581782
transform 1 0 28128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1679581782
transform 1 0 28800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1679581782
transform 1 0 29472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679581782
transform 1 0 30144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_315
timestamp 1679581782
transform 1 0 30816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_322
timestamp 1679581782
transform 1 0 31488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_329
timestamp 1679581782
transform 1 0 32160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679581782
transform 1 0 32832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679581782
transform 1 0 33504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679581782
transform 1 0 34176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_357
timestamp 1679581782
transform 1 0 34848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_364
timestamp 1679581782
transform 1 0 35520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_371
timestamp 1679581782
transform 1 0 36192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_378
timestamp 1679581782
transform 1 0 36864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_385
timestamp 1679581782
transform 1 0 37536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_392
timestamp 1679581782
transform 1 0 38208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_399
timestamp 1679581782
transform 1 0 38880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_406
timestamp 1679581782
transform 1 0 39552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679581782
transform 1 0 40224 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_420
timestamp 1677579658
transform 1 0 40896 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_433
timestamp 1679581782
transform 1 0 42144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_440
timestamp 1679581782
transform 1 0 42816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_447
timestamp 1679577901
transform 1 0 43488 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_451
timestamp 1677579658
transform 1 0 43872 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_466
timestamp 1679581782
transform 1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_478
timestamp 1679581782
transform 1 0 46464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_485
timestamp 1679581782
transform 1 0 47136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_492
timestamp 1679581782
transform 1 0 47808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_499
timestamp 1679581782
transform 1 0 48480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_506
timestamp 1679581782
transform 1 0 49152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_513
timestamp 1679577901
transform 1 0 49824 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_517
timestamp 1677580104
transform 1 0 50208 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_523
timestamp 1679581782
transform 1 0 50784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_530
timestamp 1679577901
transform 1 0 51456 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_545
timestamp 1679577901
transform 1 0 52896 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_549
timestamp 1677579658
transform 1 0 53280 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_557
timestamp 1677580104
transform 1 0 54048 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_563
timestamp 1679577901
transform 1 0 54624 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_567
timestamp 1677580104
transform 1 0 55008 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_576
timestamp 1677580104
transform 1 0 55872 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_587
timestamp 1679581782
transform 1 0 56928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_594
timestamp 1679577901
transform 1 0 57600 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_598
timestamp 1677579658
transform 1 0 57984 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_603
timestamp 1679581782
transform 1 0 58464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_610
timestamp 1679581782
transform 1 0 59136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_617
timestamp 1679581782
transform 1 0 59808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_624
timestamp 1679577901
transform 1 0 60480 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_642
timestamp 1679581782
transform 1 0 62208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_649
timestamp 1679581782
transform 1 0 62880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_656
timestamp 1679581782
transform 1 0 63552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_663
timestamp 1679581782
transform 1 0 64224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_670
timestamp 1679581782
transform 1 0 64896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_677
timestamp 1679581782
transform 1 0 65568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_684
timestamp 1679581782
transform 1 0 66240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_691
timestamp 1679581782
transform 1 0 66912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_698
timestamp 1679581782
transform 1 0 67584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_705
timestamp 1679581782
transform 1 0 68256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_712
timestamp 1679581782
transform 1 0 68928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_719
timestamp 1679581782
transform 1 0 69600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_726
timestamp 1679581782
transform 1 0 70272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_733
timestamp 1679581782
transform 1 0 70944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_740
timestamp 1679581782
transform 1 0 71616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_747
timestamp 1679581782
transform 1 0 72288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_754
timestamp 1679581782
transform 1 0 72960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_761
timestamp 1679581782
transform 1 0 73632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_768
timestamp 1679581782
transform 1 0 74304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_775
timestamp 1679581782
transform 1 0 74976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_782
timestamp 1679581782
transform 1 0 75648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_789
timestamp 1679581782
transform 1 0 76320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_796
timestamp 1679581782
transform 1 0 76992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_803
timestamp 1679581782
transform 1 0 77664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_810
timestamp 1679581782
transform 1 0 78336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_817
timestamp 1679581782
transform 1 0 79008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_824
timestamp 1679581782
transform 1 0 79680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_831
timestamp 1679581782
transform 1 0 80352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_838
timestamp 1679581782
transform 1 0 81024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_845
timestamp 1679581782
transform 1 0 81696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_852
timestamp 1679581782
transform 1 0 82368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_859
timestamp 1679581782
transform 1 0 83040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_866
timestamp 1679581782
transform 1 0 83712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_873
timestamp 1679581782
transform 1 0 84384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_880
timestamp 1679581782
transform 1 0 85056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_887
timestamp 1679581782
transform 1 0 85728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_894
timestamp 1679581782
transform 1 0 86400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_901
timestamp 1679581782
transform 1 0 87072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_908
timestamp 1679581782
transform 1 0 87744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_915
timestamp 1679581782
transform 1 0 88416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_922
timestamp 1679581782
transform 1 0 89088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_929
timestamp 1679581782
transform 1 0 89760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_936
timestamp 1679581782
transform 1 0 90432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_943
timestamp 1679581782
transform 1 0 91104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_950
timestamp 1679581782
transform 1 0 91776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_957
timestamp 1679581782
transform 1 0 92448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_964
timestamp 1679581782
transform 1 0 93120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_971
timestamp 1679581782
transform 1 0 93792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_978
timestamp 1679581782
transform 1 0 94464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_985
timestamp 1679581782
transform 1 0 95136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_992
timestamp 1679581782
transform 1 0 95808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_999
timestamp 1679581782
transform 1 0 96480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1006
timestamp 1679581782
transform 1 0 97152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1013
timestamp 1679581782
transform 1 0 97824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1020
timestamp 1679581782
transform 1 0 98496 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1027
timestamp 1677580104
transform 1 0 99168 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 9984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 10656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 12672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 20064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 22080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 22752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 23424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 24096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 24768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 25440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 26112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 26784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 27456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 28128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 28800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 29472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 30816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 31488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 32160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 32832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 33504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 34176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 34848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 35520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679581782
transform 1 0 36192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679581782
transform 1 0 36864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 37536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 38208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 38880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 39552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 40224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679581782
transform 1 0 40896 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_427
timestamp 1677579658
transform 1 0 41568 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_433
timestamp 1679581782
transform 1 0 42144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_440
timestamp 1679581782
transform 1 0 42816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_447
timestamp 1679581782
transform 1 0 43488 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_454
timestamp 1677580104
transform 1 0 44160 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_456
timestamp 1677579658
transform 1 0 44352 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_461
timestamp 1679581782
transform 1 0 44832 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_468
timestamp 1677580104
transform 1 0 45504 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_475
timestamp 1677580104
transform 1 0 46176 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_483
timestamp 1679577901
transform 1 0 46944 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_487
timestamp 1677580104
transform 1 0 47328 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_494
timestamp 1677580104
transform 1 0 48000 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_510
timestamp 1679581782
transform 1 0 49536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_517
timestamp 1679581782
transform 1 0 50208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_524
timestamp 1679581782
transform 1 0 50880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_531
timestamp 1679581782
transform 1 0 51552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_538
timestamp 1679581782
transform 1 0 52224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_545
timestamp 1679581782
transform 1 0 52896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_552
timestamp 1679581782
transform 1 0 53568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_559
timestamp 1679581782
transform 1 0 54240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_566
timestamp 1679581782
transform 1 0 54912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_573
timestamp 1679581782
transform 1 0 55584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_580
timestamp 1679581782
transform 1 0 56256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_587
timestamp 1679581782
transform 1 0 56928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_594
timestamp 1679581782
transform 1 0 57600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_601
timestamp 1679581782
transform 1 0 58272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_608
timestamp 1679581782
transform 1 0 58944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_615
timestamp 1679581782
transform 1 0 59616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_622
timestamp 1679581782
transform 1 0 60288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_629
timestamp 1679581782
transform 1 0 60960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_636
timestamp 1679581782
transform 1 0 61632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_643
timestamp 1679581782
transform 1 0 62304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_650
timestamp 1679581782
transform 1 0 62976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_657
timestamp 1679581782
transform 1 0 63648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_664
timestamp 1679581782
transform 1 0 64320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_671
timestamp 1679581782
transform 1 0 64992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_678
timestamp 1679581782
transform 1 0 65664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_685
timestamp 1679581782
transform 1 0 66336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_692
timestamp 1679581782
transform 1 0 67008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_699
timestamp 1679581782
transform 1 0 67680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_706
timestamp 1679581782
transform 1 0 68352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_713
timestamp 1679581782
transform 1 0 69024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_720
timestamp 1679581782
transform 1 0 69696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_727
timestamp 1679581782
transform 1 0 70368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_734
timestamp 1679581782
transform 1 0 71040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_741
timestamp 1679581782
transform 1 0 71712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_748
timestamp 1679581782
transform 1 0 72384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_755
timestamp 1679581782
transform 1 0 73056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_762
timestamp 1679581782
transform 1 0 73728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_769
timestamp 1679581782
transform 1 0 74400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_776
timestamp 1679581782
transform 1 0 75072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_783
timestamp 1679581782
transform 1 0 75744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_790
timestamp 1679581782
transform 1 0 76416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_797
timestamp 1679581782
transform 1 0 77088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_804
timestamp 1679581782
transform 1 0 77760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_811
timestamp 1679581782
transform 1 0 78432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_818
timestamp 1679581782
transform 1 0 79104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_825
timestamp 1679581782
transform 1 0 79776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_832
timestamp 1679581782
transform 1 0 80448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_839
timestamp 1679581782
transform 1 0 81120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_846
timestamp 1679581782
transform 1 0 81792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_853
timestamp 1679581782
transform 1 0 82464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_860
timestamp 1679581782
transform 1 0 83136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_867
timestamp 1679581782
transform 1 0 83808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_874
timestamp 1679581782
transform 1 0 84480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_881
timestamp 1679581782
transform 1 0 85152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_888
timestamp 1679581782
transform 1 0 85824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_895
timestamp 1679581782
transform 1 0 86496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_902
timestamp 1679581782
transform 1 0 87168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_909
timestamp 1679581782
transform 1 0 87840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_916
timestamp 1679581782
transform 1 0 88512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_923
timestamp 1679581782
transform 1 0 89184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_930
timestamp 1679581782
transform 1 0 89856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_937
timestamp 1679581782
transform 1 0 90528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_944
timestamp 1679581782
transform 1 0 91200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_951
timestamp 1679581782
transform 1 0 91872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_958
timestamp 1679581782
transform 1 0 92544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_965
timestamp 1679581782
transform 1 0 93216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_972
timestamp 1679581782
transform 1 0 93888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_979
timestamp 1679581782
transform 1 0 94560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_986
timestamp 1679581782
transform 1 0 95232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_993
timestamp 1679581782
transform 1 0 95904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1000
timestamp 1679581782
transform 1 0 96576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1007
timestamp 1679581782
transform 1 0 97248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1014
timestamp 1679581782
transform 1 0 97920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1021
timestamp 1679581782
transform 1 0 98592 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677579658
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 1920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 2592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 3936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 4608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 5952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 6624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 7968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 8640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 9984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 10656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 12672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 14688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 16704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 18048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679581782
transform 1 0 18720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 19392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679581782
transform 1 0 20064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679581782
transform 1 0 20736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679581782
transform 1 0 21408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_224
timestamp 1679581782
transform 1 0 22080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_231
timestamp 1679581782
transform 1 0 22752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_238
timestamp 1679581782
transform 1 0 23424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_245
timestamp 1679581782
transform 1 0 24096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_252
timestamp 1679581782
transform 1 0 24768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1679581782
transform 1 0 25440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_266
timestamp 1679581782
transform 1 0 26112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_273
timestamp 1679581782
transform 1 0 26784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_280
timestamp 1679581782
transform 1 0 27456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_287
timestamp 1679581782
transform 1 0 28128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_294
timestamp 1679581782
transform 1 0 28800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_301
timestamp 1679581782
transform 1 0 29472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_308
timestamp 1679581782
transform 1 0 30144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_315
timestamp 1679581782
transform 1 0 30816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_322
timestamp 1679581782
transform 1 0 31488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_329
timestamp 1679581782
transform 1 0 32160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_336
timestamp 1679581782
transform 1 0 32832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_343
timestamp 1679581782
transform 1 0 33504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_350
timestamp 1679581782
transform 1 0 34176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_357
timestamp 1679581782
transform 1 0 34848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_364
timestamp 1679581782
transform 1 0 35520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_371
timestamp 1679581782
transform 1 0 36192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_378
timestamp 1679581782
transform 1 0 36864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_385
timestamp 1679581782
transform 1 0 37536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679581782
transform 1 0 38208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_399
timestamp 1679581782
transform 1 0 38880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679581782
transform 1 0 39552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679581782
transform 1 0 40224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679581782
transform 1 0 40896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679581782
transform 1 0 41568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679581782
transform 1 0 42240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 42912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 43584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 44256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 44928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 45600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 46272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 46944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679581782
transform 1 0 47616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679581782
transform 1 0 48288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679581782
transform 1 0 48960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679581782
transform 1 0 49632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_518
timestamp 1679581782
transform 1 0 50304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_525
timestamp 1679581782
transform 1 0 50976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_532
timestamp 1679581782
transform 1 0 51648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_539
timestamp 1679581782
transform 1 0 52320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_546
timestamp 1679581782
transform 1 0 52992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_553
timestamp 1679581782
transform 1 0 53664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_560
timestamp 1679581782
transform 1 0 54336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_567
timestamp 1679581782
transform 1 0 55008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_574
timestamp 1679581782
transform 1 0 55680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_581
timestamp 1679581782
transform 1 0 56352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_588
timestamp 1679581782
transform 1 0 57024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_595
timestamp 1679581782
transform 1 0 57696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_602
timestamp 1679581782
transform 1 0 58368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_609
timestamp 1679581782
transform 1 0 59040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_616
timestamp 1679581782
transform 1 0 59712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_623
timestamp 1679581782
transform 1 0 60384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_630
timestamp 1679581782
transform 1 0 61056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_637
timestamp 1679581782
transform 1 0 61728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_644
timestamp 1679581782
transform 1 0 62400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_651
timestamp 1679581782
transform 1 0 63072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_658
timestamp 1679581782
transform 1 0 63744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_665
timestamp 1679581782
transform 1 0 64416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_672
timestamp 1679581782
transform 1 0 65088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_679
timestamp 1679581782
transform 1 0 65760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_686
timestamp 1679581782
transform 1 0 66432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_693
timestamp 1679581782
transform 1 0 67104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_700
timestamp 1679581782
transform 1 0 67776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_707
timestamp 1679581782
transform 1 0 68448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_714
timestamp 1679581782
transform 1 0 69120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_721
timestamp 1679581782
transform 1 0 69792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 70464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_735
timestamp 1679581782
transform 1 0 71136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_742
timestamp 1679581782
transform 1 0 71808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_749
timestamp 1679581782
transform 1 0 72480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_756
timestamp 1679581782
transform 1 0 73152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_763
timestamp 1679581782
transform 1 0 73824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_770
timestamp 1679581782
transform 1 0 74496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_777
timestamp 1679581782
transform 1 0 75168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_784
timestamp 1679581782
transform 1 0 75840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_791
timestamp 1679581782
transform 1 0 76512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_798
timestamp 1679581782
transform 1 0 77184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_805
timestamp 1679581782
transform 1 0 77856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_812
timestamp 1679581782
transform 1 0 78528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_819
timestamp 1679581782
transform 1 0 79200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_826
timestamp 1679581782
transform 1 0 79872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_833
timestamp 1679581782
transform 1 0 80544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_840
timestamp 1679581782
transform 1 0 81216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_847
timestamp 1679581782
transform 1 0 81888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_854
timestamp 1679581782
transform 1 0 82560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_861
timestamp 1679581782
transform 1 0 83232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_868
timestamp 1679581782
transform 1 0 83904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_875
timestamp 1679581782
transform 1 0 84576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_882
timestamp 1679581782
transform 1 0 85248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_889
timestamp 1679581782
transform 1 0 85920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_896
timestamp 1679581782
transform 1 0 86592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_903
timestamp 1679581782
transform 1 0 87264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_910
timestamp 1679581782
transform 1 0 87936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_917
timestamp 1679581782
transform 1 0 88608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_924
timestamp 1679581782
transform 1 0 89280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_931
timestamp 1679581782
transform 1 0 89952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_938
timestamp 1679581782
transform 1 0 90624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_945
timestamp 1679581782
transform 1 0 91296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_952
timestamp 1679581782
transform 1 0 91968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_959
timestamp 1679581782
transform 1 0 92640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_966
timestamp 1679581782
transform 1 0 93312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_973
timestamp 1679581782
transform 1 0 93984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_980
timestamp 1679581782
transform 1 0 94656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_987
timestamp 1679581782
transform 1 0 95328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_994
timestamp 1679581782
transform 1 0 96000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1001
timestamp 1679581782
transform 1 0 96672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1008
timestamp 1679581782
transform 1 0 97344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1015
timestamp 1679581782
transform 1 0 98016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1022
timestamp 1679581782
transform 1 0 98688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 1920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 2592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 3936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 4608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 5952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 6624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 7968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 8640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 9984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 10656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 12672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 14688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 16704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 18720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 20736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 21408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 22080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 22752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 23424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 24768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 25440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679581782
transform 1 0 26112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679581782
transform 1 0 26784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679581782
transform 1 0 27456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679581782
transform 1 0 28128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679581782
transform 1 0 28800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679581782
transform 1 0 29472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679581782
transform 1 0 30144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679581782
transform 1 0 30816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679581782
transform 1 0 31488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679581782
transform 1 0 32160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679581782
transform 1 0 32832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679581782
transform 1 0 33504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679581782
transform 1 0 34176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679581782
transform 1 0 34848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 35520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679581782
transform 1 0 36192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679581782
transform 1 0 36864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679581782
transform 1 0 37536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679581782
transform 1 0 38208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679581782
transform 1 0 38880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679581782
transform 1 0 39552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679581782
transform 1 0 40224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679581782
transform 1 0 40896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679581782
transform 1 0 41568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679581782
transform 1 0 42240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679581782
transform 1 0 42912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_448
timestamp 1679581782
transform 1 0 43584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_455
timestamp 1679581782
transform 1 0 44256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_462
timestamp 1679581782
transform 1 0 44928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_469
timestamp 1679581782
transform 1 0 45600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_476
timestamp 1679581782
transform 1 0 46272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_483
timestamp 1679581782
transform 1 0 46944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679581782
transform 1 0 47616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_497
timestamp 1679581782
transform 1 0 48288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_504
timestamp 1679581782
transform 1 0 48960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_511
timestamp 1679581782
transform 1 0 49632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_518
timestamp 1679581782
transform 1 0 50304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_525
timestamp 1679581782
transform 1 0 50976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_532
timestamp 1679581782
transform 1 0 51648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_539
timestamp 1679581782
transform 1 0 52320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_546
timestamp 1679581782
transform 1 0 52992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_553
timestamp 1679581782
transform 1 0 53664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_560
timestamp 1679581782
transform 1 0 54336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_567
timestamp 1679581782
transform 1 0 55008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_574
timestamp 1679581782
transform 1 0 55680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_581
timestamp 1679581782
transform 1 0 56352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_588
timestamp 1679581782
transform 1 0 57024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_595
timestamp 1679581782
transform 1 0 57696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_602
timestamp 1679581782
transform 1 0 58368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_609
timestamp 1679581782
transform 1 0 59040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_616
timestamp 1679581782
transform 1 0 59712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_623
timestamp 1679581782
transform 1 0 60384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_630
timestamp 1679581782
transform 1 0 61056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_637
timestamp 1679581782
transform 1 0 61728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_644
timestamp 1679581782
transform 1 0 62400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_651
timestamp 1679581782
transform 1 0 63072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_658
timestamp 1679581782
transform 1 0 63744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_665
timestamp 1679581782
transform 1 0 64416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_672
timestamp 1679581782
transform 1 0 65088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_679
timestamp 1679581782
transform 1 0 65760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_686
timestamp 1679581782
transform 1 0 66432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_693
timestamp 1679581782
transform 1 0 67104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_700
timestamp 1679581782
transform 1 0 67776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_707
timestamp 1679581782
transform 1 0 68448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_714
timestamp 1679581782
transform 1 0 69120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_721
timestamp 1679581782
transform 1 0 69792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_728
timestamp 1679581782
transform 1 0 70464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_735
timestamp 1679581782
transform 1 0 71136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679581782
transform 1 0 71808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679581782
transform 1 0 72480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_756
timestamp 1679581782
transform 1 0 73152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_763
timestamp 1679581782
transform 1 0 73824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_770
timestamp 1679581782
transform 1 0 74496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_777
timestamp 1679581782
transform 1 0 75168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_784
timestamp 1679581782
transform 1 0 75840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_791
timestamp 1679581782
transform 1 0 76512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_798
timestamp 1679581782
transform 1 0 77184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_805
timestamp 1679581782
transform 1 0 77856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_812
timestamp 1679581782
transform 1 0 78528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_819
timestamp 1679581782
transform 1 0 79200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_826
timestamp 1679581782
transform 1 0 79872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_833
timestamp 1679581782
transform 1 0 80544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_840
timestamp 1679581782
transform 1 0 81216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_847
timestamp 1679581782
transform 1 0 81888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_854
timestamp 1679581782
transform 1 0 82560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_861
timestamp 1679581782
transform 1 0 83232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_868
timestamp 1679581782
transform 1 0 83904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_875
timestamp 1679581782
transform 1 0 84576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_882
timestamp 1679581782
transform 1 0 85248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_889
timestamp 1679581782
transform 1 0 85920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_896
timestamp 1679581782
transform 1 0 86592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_903
timestamp 1679581782
transform 1 0 87264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_910
timestamp 1679581782
transform 1 0 87936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_917
timestamp 1679581782
transform 1 0 88608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_924
timestamp 1679581782
transform 1 0 89280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_931
timestamp 1679581782
transform 1 0 89952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_938
timestamp 1679581782
transform 1 0 90624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_945
timestamp 1679581782
transform 1 0 91296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_952
timestamp 1679581782
transform 1 0 91968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_959
timestamp 1679581782
transform 1 0 92640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_966
timestamp 1679581782
transform 1 0 93312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_973
timestamp 1679581782
transform 1 0 93984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_980
timestamp 1679581782
transform 1 0 94656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_987
timestamp 1679581782
transform 1 0 95328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_994
timestamp 1679581782
transform 1 0 96000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1001
timestamp 1679581782
transform 1 0 96672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1008
timestamp 1679581782
transform 1 0 97344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1015
timestamp 1679581782
transform 1 0 98016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1022
timestamp 1679581782
transform 1 0 98688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 1920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 2592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 3936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 4608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 5952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 6624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 7968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 8640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 9984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 10656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 11328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679581782
transform 1 0 12000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_126
timestamp 1679581782
transform 1 0 12672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_133
timestamp 1679581782
transform 1 0 13344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679581782
transform 1 0 14016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_147
timestamp 1679581782
transform 1 0 14688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679581782
transform 1 0 15360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_161
timestamp 1679581782
transform 1 0 16032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_168
timestamp 1679581782
transform 1 0 16704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_175
timestamp 1679581782
transform 1 0 17376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_182
timestamp 1679581782
transform 1 0 18048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679581782
transform 1 0 18720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_196
timestamp 1679581782
transform 1 0 19392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679581782
transform 1 0 20064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_210
timestamp 1679581782
transform 1 0 20736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_217
timestamp 1679581782
transform 1 0 21408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_224
timestamp 1679581782
transform 1 0 22080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_231
timestamp 1679581782
transform 1 0 22752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_238
timestamp 1679581782
transform 1 0 23424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_245
timestamp 1679581782
transform 1 0 24096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_252
timestamp 1679581782
transform 1 0 24768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_259
timestamp 1679581782
transform 1 0 25440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_266
timestamp 1679581782
transform 1 0 26112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679581782
transform 1 0 26784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679581782
transform 1 0 27456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_287
timestamp 1679581782
transform 1 0 28128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_294
timestamp 1679581782
transform 1 0 28800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_301
timestamp 1679581782
transform 1 0 29472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_308
timestamp 1679581782
transform 1 0 30144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_315
timestamp 1679581782
transform 1 0 30816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_322
timestamp 1679581782
transform 1 0 31488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_329
timestamp 1679581782
transform 1 0 32160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_336
timestamp 1679581782
transform 1 0 32832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_343
timestamp 1679581782
transform 1 0 33504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_350
timestamp 1679581782
transform 1 0 34176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_357
timestamp 1679581782
transform 1 0 34848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_364
timestamp 1679581782
transform 1 0 35520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_371
timestamp 1679581782
transform 1 0 36192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_378
timestamp 1679581782
transform 1 0 36864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_385
timestamp 1679581782
transform 1 0 37536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_392
timestamp 1679581782
transform 1 0 38208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_399
timestamp 1679581782
transform 1 0 38880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_406
timestamp 1679581782
transform 1 0 39552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_413
timestamp 1679581782
transform 1 0 40224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_420
timestamp 1679581782
transform 1 0 40896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_427
timestamp 1679581782
transform 1 0 41568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_434
timestamp 1679581782
transform 1 0 42240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_441
timestamp 1679581782
transform 1 0 42912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_448
timestamp 1679581782
transform 1 0 43584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_455
timestamp 1679581782
transform 1 0 44256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_462
timestamp 1679581782
transform 1 0 44928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_469
timestamp 1679581782
transform 1 0 45600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_476
timestamp 1679581782
transform 1 0 46272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_483
timestamp 1679581782
transform 1 0 46944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_490
timestamp 1679581782
transform 1 0 47616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_497
timestamp 1679581782
transform 1 0 48288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_504
timestamp 1679581782
transform 1 0 48960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_511
timestamp 1679581782
transform 1 0 49632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_518
timestamp 1679581782
transform 1 0 50304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_525
timestamp 1679581782
transform 1 0 50976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_532
timestamp 1679581782
transform 1 0 51648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_539
timestamp 1679581782
transform 1 0 52320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_546
timestamp 1679581782
transform 1 0 52992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_553
timestamp 1679581782
transform 1 0 53664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_560
timestamp 1679581782
transform 1 0 54336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_567
timestamp 1679581782
transform 1 0 55008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_574
timestamp 1679581782
transform 1 0 55680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_581
timestamp 1679581782
transform 1 0 56352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_588
timestamp 1679581782
transform 1 0 57024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_595
timestamp 1679581782
transform 1 0 57696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_602
timestamp 1679581782
transform 1 0 58368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_609
timestamp 1679581782
transform 1 0 59040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_616
timestamp 1679581782
transform 1 0 59712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_623
timestamp 1679581782
transform 1 0 60384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_630
timestamp 1679581782
transform 1 0 61056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_637
timestamp 1679581782
transform 1 0 61728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_644
timestamp 1679581782
transform 1 0 62400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_651
timestamp 1679581782
transform 1 0 63072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_658
timestamp 1679581782
transform 1 0 63744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_665
timestamp 1679581782
transform 1 0 64416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_672
timestamp 1679581782
transform 1 0 65088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_679
timestamp 1679581782
transform 1 0 65760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_686
timestamp 1679581782
transform 1 0 66432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_693
timestamp 1679581782
transform 1 0 67104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_700
timestamp 1679581782
transform 1 0 67776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_707
timestamp 1679581782
transform 1 0 68448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_714
timestamp 1679581782
transform 1 0 69120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_721
timestamp 1679581782
transform 1 0 69792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_728
timestamp 1679581782
transform 1 0 70464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_735
timestamp 1679581782
transform 1 0 71136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_742
timestamp 1679581782
transform 1 0 71808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_749
timestamp 1679581782
transform 1 0 72480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_756
timestamp 1679581782
transform 1 0 73152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_763
timestamp 1679581782
transform 1 0 73824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_770
timestamp 1679581782
transform 1 0 74496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_777
timestamp 1679581782
transform 1 0 75168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_784
timestamp 1679581782
transform 1 0 75840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_791
timestamp 1679581782
transform 1 0 76512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_798
timestamp 1679581782
transform 1 0 77184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_805
timestamp 1679581782
transform 1 0 77856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_812
timestamp 1679581782
transform 1 0 78528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_819
timestamp 1679581782
transform 1 0 79200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_826
timestamp 1679581782
transform 1 0 79872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_833
timestamp 1679581782
transform 1 0 80544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_840
timestamp 1679581782
transform 1 0 81216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_847
timestamp 1679581782
transform 1 0 81888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_854
timestamp 1679581782
transform 1 0 82560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_861
timestamp 1679581782
transform 1 0 83232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_868
timestamp 1679581782
transform 1 0 83904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_875
timestamp 1679581782
transform 1 0 84576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_882
timestamp 1679581782
transform 1 0 85248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_889
timestamp 1679581782
transform 1 0 85920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_896
timestamp 1679581782
transform 1 0 86592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_903
timestamp 1679581782
transform 1 0 87264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_910
timestamp 1679581782
transform 1 0 87936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_917
timestamp 1679581782
transform 1 0 88608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_924
timestamp 1679581782
transform 1 0 89280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_931
timestamp 1679581782
transform 1 0 89952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_938
timestamp 1679581782
transform 1 0 90624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_945
timestamp 1679581782
transform 1 0 91296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_952
timestamp 1679581782
transform 1 0 91968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_959
timestamp 1679581782
transform 1 0 92640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_966
timestamp 1679581782
transform 1 0 93312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_973
timestamp 1679581782
transform 1 0 93984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_980
timestamp 1679581782
transform 1 0 94656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_987
timestamp 1679581782
transform 1 0 95328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_994
timestamp 1679581782
transform 1 0 96000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1001
timestamp 1679581782
transform 1 0 96672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1008
timestamp 1679581782
transform 1 0 97344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1015
timestamp 1679581782
transform 1 0 98016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1022
timestamp 1679581782
transform 1 0 98688 0 1 8316
box -48 -56 720 834
<< labels >>
flabel metal6 s 4316 630 4756 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 9116 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 4496 99404 4936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 9198 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 3256 99404 3696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6200 9920 6280 10000 0 FreeSans 320 0 0 0 ena_i
port 2 nsew signal input
flabel metal2 s 17144 9920 17224 10000 0 FreeSans 320 0 0 0 input_ni[0]
port 3 nsew signal input
flabel metal2 s 28088 9920 28168 10000 0 FreeSans 320 0 0 0 input_ni[1]
port 4 nsew signal input
flabel metal2 s 39032 9920 39112 10000 0 FreeSans 320 0 0 0 input_ni[2]
port 5 nsew signal input
flabel metal2 s 49976 9920 50056 10000 0 FreeSans 320 0 0 0 input_ni[3]
port 6 nsew signal input
flabel metal2 s 60920 9920 61000 10000 0 FreeSans 320 0 0 0 input_ni[4]
port 7 nsew signal input
flabel metal2 s 71864 9920 71944 10000 0 FreeSans 320 0 0 0 input_ni[5]
port 8 nsew signal input
flabel metal2 s 82808 9920 82888 10000 0 FreeSans 320 0 0 0 input_ni[6]
port 9 nsew signal input
flabel metal2 s 93752 9920 93832 10000 0 FreeSans 320 0 0 0 input_ni[7]
port 10 nsew signal input
flabel metal2 s 824 0 904 80 0 FreeSans 320 0 0 0 output_no[0]
port 11 nsew signal output
flabel metal2 s 39224 0 39304 80 0 FreeSans 320 0 0 0 output_no[100]
port 12 nsew signal output
flabel metal2 s 39608 0 39688 80 0 FreeSans 320 0 0 0 output_no[101]
port 13 nsew signal output
flabel metal2 s 39992 0 40072 80 0 FreeSans 320 0 0 0 output_no[102]
port 14 nsew signal output
flabel metal2 s 40376 0 40456 80 0 FreeSans 320 0 0 0 output_no[103]
port 15 nsew signal output
flabel metal2 s 40760 0 40840 80 0 FreeSans 320 0 0 0 output_no[104]
port 16 nsew signal output
flabel metal2 s 41144 0 41224 80 0 FreeSans 320 0 0 0 output_no[105]
port 17 nsew signal output
flabel metal2 s 41528 0 41608 80 0 FreeSans 320 0 0 0 output_no[106]
port 18 nsew signal output
flabel metal2 s 41912 0 41992 80 0 FreeSans 320 0 0 0 output_no[107]
port 19 nsew signal output
flabel metal2 s 42296 0 42376 80 0 FreeSans 320 0 0 0 output_no[108]
port 20 nsew signal output
flabel metal2 s 42680 0 42760 80 0 FreeSans 320 0 0 0 output_no[109]
port 21 nsew signal output
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 output_no[10]
port 22 nsew signal output
flabel metal2 s 43064 0 43144 80 0 FreeSans 320 0 0 0 output_no[110]
port 23 nsew signal output
flabel metal2 s 43448 0 43528 80 0 FreeSans 320 0 0 0 output_no[111]
port 24 nsew signal output
flabel metal2 s 43832 0 43912 80 0 FreeSans 320 0 0 0 output_no[112]
port 25 nsew signal output
flabel metal2 s 44216 0 44296 80 0 FreeSans 320 0 0 0 output_no[113]
port 26 nsew signal output
flabel metal2 s 44600 0 44680 80 0 FreeSans 320 0 0 0 output_no[114]
port 27 nsew signal output
flabel metal2 s 44984 0 45064 80 0 FreeSans 320 0 0 0 output_no[115]
port 28 nsew signal output
flabel metal2 s 45368 0 45448 80 0 FreeSans 320 0 0 0 output_no[116]
port 29 nsew signal output
flabel metal2 s 45752 0 45832 80 0 FreeSans 320 0 0 0 output_no[117]
port 30 nsew signal output
flabel metal2 s 46136 0 46216 80 0 FreeSans 320 0 0 0 output_no[118]
port 31 nsew signal output
flabel metal2 s 46520 0 46600 80 0 FreeSans 320 0 0 0 output_no[119]
port 32 nsew signal output
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 output_no[11]
port 33 nsew signal output
flabel metal2 s 46904 0 46984 80 0 FreeSans 320 0 0 0 output_no[120]
port 34 nsew signal output
flabel metal2 s 47288 0 47368 80 0 FreeSans 320 0 0 0 output_no[121]
port 35 nsew signal output
flabel metal2 s 47672 0 47752 80 0 FreeSans 320 0 0 0 output_no[122]
port 36 nsew signal output
flabel metal2 s 48056 0 48136 80 0 FreeSans 320 0 0 0 output_no[123]
port 37 nsew signal output
flabel metal2 s 48440 0 48520 80 0 FreeSans 320 0 0 0 output_no[124]
port 38 nsew signal output
flabel metal2 s 48824 0 48904 80 0 FreeSans 320 0 0 0 output_no[125]
port 39 nsew signal output
flabel metal2 s 49208 0 49288 80 0 FreeSans 320 0 0 0 output_no[126]
port 40 nsew signal output
flabel metal2 s 49592 0 49672 80 0 FreeSans 320 0 0 0 output_no[127]
port 41 nsew signal output
flabel metal2 s 49976 0 50056 80 0 FreeSans 320 0 0 0 output_no[128]
port 42 nsew signal output
flabel metal2 s 50360 0 50440 80 0 FreeSans 320 0 0 0 output_no[129]
port 43 nsew signal output
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 output_no[12]
port 44 nsew signal output
flabel metal2 s 50744 0 50824 80 0 FreeSans 320 0 0 0 output_no[130]
port 45 nsew signal output
flabel metal2 s 51128 0 51208 80 0 FreeSans 320 0 0 0 output_no[131]
port 46 nsew signal output
flabel metal2 s 51512 0 51592 80 0 FreeSans 320 0 0 0 output_no[132]
port 47 nsew signal output
flabel metal2 s 51896 0 51976 80 0 FreeSans 320 0 0 0 output_no[133]
port 48 nsew signal output
flabel metal2 s 52280 0 52360 80 0 FreeSans 320 0 0 0 output_no[134]
port 49 nsew signal output
flabel metal2 s 52664 0 52744 80 0 FreeSans 320 0 0 0 output_no[135]
port 50 nsew signal output
flabel metal2 s 53048 0 53128 80 0 FreeSans 320 0 0 0 output_no[136]
port 51 nsew signal output
flabel metal2 s 53432 0 53512 80 0 FreeSans 320 0 0 0 output_no[137]
port 52 nsew signal output
flabel metal2 s 53816 0 53896 80 0 FreeSans 320 0 0 0 output_no[138]
port 53 nsew signal output
flabel metal2 s 54200 0 54280 80 0 FreeSans 320 0 0 0 output_no[139]
port 54 nsew signal output
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 output_no[13]
port 55 nsew signal output
flabel metal2 s 54584 0 54664 80 0 FreeSans 320 0 0 0 output_no[140]
port 56 nsew signal output
flabel metal2 s 54968 0 55048 80 0 FreeSans 320 0 0 0 output_no[141]
port 57 nsew signal output
flabel metal2 s 55352 0 55432 80 0 FreeSans 320 0 0 0 output_no[142]
port 58 nsew signal output
flabel metal2 s 55736 0 55816 80 0 FreeSans 320 0 0 0 output_no[143]
port 59 nsew signal output
flabel metal2 s 56120 0 56200 80 0 FreeSans 320 0 0 0 output_no[144]
port 60 nsew signal output
flabel metal2 s 56504 0 56584 80 0 FreeSans 320 0 0 0 output_no[145]
port 61 nsew signal output
flabel metal2 s 56888 0 56968 80 0 FreeSans 320 0 0 0 output_no[146]
port 62 nsew signal output
flabel metal2 s 57272 0 57352 80 0 FreeSans 320 0 0 0 output_no[147]
port 63 nsew signal output
flabel metal2 s 57656 0 57736 80 0 FreeSans 320 0 0 0 output_no[148]
port 64 nsew signal output
flabel metal2 s 58040 0 58120 80 0 FreeSans 320 0 0 0 output_no[149]
port 65 nsew signal output
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 output_no[14]
port 66 nsew signal output
flabel metal2 s 58424 0 58504 80 0 FreeSans 320 0 0 0 output_no[150]
port 67 nsew signal output
flabel metal2 s 58808 0 58888 80 0 FreeSans 320 0 0 0 output_no[151]
port 68 nsew signal output
flabel metal2 s 59192 0 59272 80 0 FreeSans 320 0 0 0 output_no[152]
port 69 nsew signal output
flabel metal2 s 59576 0 59656 80 0 FreeSans 320 0 0 0 output_no[153]
port 70 nsew signal output
flabel metal2 s 59960 0 60040 80 0 FreeSans 320 0 0 0 output_no[154]
port 71 nsew signal output
flabel metal2 s 60344 0 60424 80 0 FreeSans 320 0 0 0 output_no[155]
port 72 nsew signal output
flabel metal2 s 60728 0 60808 80 0 FreeSans 320 0 0 0 output_no[156]
port 73 nsew signal output
flabel metal2 s 61112 0 61192 80 0 FreeSans 320 0 0 0 output_no[157]
port 74 nsew signal output
flabel metal2 s 61496 0 61576 80 0 FreeSans 320 0 0 0 output_no[158]
port 75 nsew signal output
flabel metal2 s 61880 0 61960 80 0 FreeSans 320 0 0 0 output_no[159]
port 76 nsew signal output
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 output_no[15]
port 77 nsew signal output
flabel metal2 s 62264 0 62344 80 0 FreeSans 320 0 0 0 output_no[160]
port 78 nsew signal output
flabel metal2 s 62648 0 62728 80 0 FreeSans 320 0 0 0 output_no[161]
port 79 nsew signal output
flabel metal2 s 63032 0 63112 80 0 FreeSans 320 0 0 0 output_no[162]
port 80 nsew signal output
flabel metal2 s 63416 0 63496 80 0 FreeSans 320 0 0 0 output_no[163]
port 81 nsew signal output
flabel metal2 s 63800 0 63880 80 0 FreeSans 320 0 0 0 output_no[164]
port 82 nsew signal output
flabel metal2 s 64184 0 64264 80 0 FreeSans 320 0 0 0 output_no[165]
port 83 nsew signal output
flabel metal2 s 64568 0 64648 80 0 FreeSans 320 0 0 0 output_no[166]
port 84 nsew signal output
flabel metal2 s 64952 0 65032 80 0 FreeSans 320 0 0 0 output_no[167]
port 85 nsew signal output
flabel metal2 s 65336 0 65416 80 0 FreeSans 320 0 0 0 output_no[168]
port 86 nsew signal output
flabel metal2 s 65720 0 65800 80 0 FreeSans 320 0 0 0 output_no[169]
port 87 nsew signal output
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 output_no[16]
port 88 nsew signal output
flabel metal2 s 66104 0 66184 80 0 FreeSans 320 0 0 0 output_no[170]
port 89 nsew signal output
flabel metal2 s 66488 0 66568 80 0 FreeSans 320 0 0 0 output_no[171]
port 90 nsew signal output
flabel metal2 s 66872 0 66952 80 0 FreeSans 320 0 0 0 output_no[172]
port 91 nsew signal output
flabel metal2 s 67256 0 67336 80 0 FreeSans 320 0 0 0 output_no[173]
port 92 nsew signal output
flabel metal2 s 67640 0 67720 80 0 FreeSans 320 0 0 0 output_no[174]
port 93 nsew signal output
flabel metal2 s 68024 0 68104 80 0 FreeSans 320 0 0 0 output_no[175]
port 94 nsew signal output
flabel metal2 s 68408 0 68488 80 0 FreeSans 320 0 0 0 output_no[176]
port 95 nsew signal output
flabel metal2 s 68792 0 68872 80 0 FreeSans 320 0 0 0 output_no[177]
port 96 nsew signal output
flabel metal2 s 69176 0 69256 80 0 FreeSans 320 0 0 0 output_no[178]
port 97 nsew signal output
flabel metal2 s 69560 0 69640 80 0 FreeSans 320 0 0 0 output_no[179]
port 98 nsew signal output
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 output_no[17]
port 99 nsew signal output
flabel metal2 s 69944 0 70024 80 0 FreeSans 320 0 0 0 output_no[180]
port 100 nsew signal output
flabel metal2 s 70328 0 70408 80 0 FreeSans 320 0 0 0 output_no[181]
port 101 nsew signal output
flabel metal2 s 70712 0 70792 80 0 FreeSans 320 0 0 0 output_no[182]
port 102 nsew signal output
flabel metal2 s 71096 0 71176 80 0 FreeSans 320 0 0 0 output_no[183]
port 103 nsew signal output
flabel metal2 s 71480 0 71560 80 0 FreeSans 320 0 0 0 output_no[184]
port 104 nsew signal output
flabel metal2 s 71864 0 71944 80 0 FreeSans 320 0 0 0 output_no[185]
port 105 nsew signal output
flabel metal2 s 72248 0 72328 80 0 FreeSans 320 0 0 0 output_no[186]
port 106 nsew signal output
flabel metal2 s 72632 0 72712 80 0 FreeSans 320 0 0 0 output_no[187]
port 107 nsew signal output
flabel metal2 s 73016 0 73096 80 0 FreeSans 320 0 0 0 output_no[188]
port 108 nsew signal output
flabel metal2 s 73400 0 73480 80 0 FreeSans 320 0 0 0 output_no[189]
port 109 nsew signal output
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 output_no[18]
port 110 nsew signal output
flabel metal2 s 73784 0 73864 80 0 FreeSans 320 0 0 0 output_no[190]
port 111 nsew signal output
flabel metal2 s 74168 0 74248 80 0 FreeSans 320 0 0 0 output_no[191]
port 112 nsew signal output
flabel metal2 s 74552 0 74632 80 0 FreeSans 320 0 0 0 output_no[192]
port 113 nsew signal output
flabel metal2 s 74936 0 75016 80 0 FreeSans 320 0 0 0 output_no[193]
port 114 nsew signal output
flabel metal2 s 75320 0 75400 80 0 FreeSans 320 0 0 0 output_no[194]
port 115 nsew signal output
flabel metal2 s 75704 0 75784 80 0 FreeSans 320 0 0 0 output_no[195]
port 116 nsew signal output
flabel metal2 s 76088 0 76168 80 0 FreeSans 320 0 0 0 output_no[196]
port 117 nsew signal output
flabel metal2 s 76472 0 76552 80 0 FreeSans 320 0 0 0 output_no[197]
port 118 nsew signal output
flabel metal2 s 76856 0 76936 80 0 FreeSans 320 0 0 0 output_no[198]
port 119 nsew signal output
flabel metal2 s 77240 0 77320 80 0 FreeSans 320 0 0 0 output_no[199]
port 120 nsew signal output
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 output_no[19]
port 121 nsew signal output
flabel metal2 s 1208 0 1288 80 0 FreeSans 320 0 0 0 output_no[1]
port 122 nsew signal output
flabel metal2 s 77624 0 77704 80 0 FreeSans 320 0 0 0 output_no[200]
port 123 nsew signal output
flabel metal2 s 78008 0 78088 80 0 FreeSans 320 0 0 0 output_no[201]
port 124 nsew signal output
flabel metal2 s 78392 0 78472 80 0 FreeSans 320 0 0 0 output_no[202]
port 125 nsew signal output
flabel metal2 s 78776 0 78856 80 0 FreeSans 320 0 0 0 output_no[203]
port 126 nsew signal output
flabel metal2 s 79160 0 79240 80 0 FreeSans 320 0 0 0 output_no[204]
port 127 nsew signal output
flabel metal2 s 79544 0 79624 80 0 FreeSans 320 0 0 0 output_no[205]
port 128 nsew signal output
flabel metal2 s 79928 0 80008 80 0 FreeSans 320 0 0 0 output_no[206]
port 129 nsew signal output
flabel metal2 s 80312 0 80392 80 0 FreeSans 320 0 0 0 output_no[207]
port 130 nsew signal output
flabel metal2 s 80696 0 80776 80 0 FreeSans 320 0 0 0 output_no[208]
port 131 nsew signal output
flabel metal2 s 81080 0 81160 80 0 FreeSans 320 0 0 0 output_no[209]
port 132 nsew signal output
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 output_no[20]
port 133 nsew signal output
flabel metal2 s 81464 0 81544 80 0 FreeSans 320 0 0 0 output_no[210]
port 134 nsew signal output
flabel metal2 s 81848 0 81928 80 0 FreeSans 320 0 0 0 output_no[211]
port 135 nsew signal output
flabel metal2 s 82232 0 82312 80 0 FreeSans 320 0 0 0 output_no[212]
port 136 nsew signal output
flabel metal2 s 82616 0 82696 80 0 FreeSans 320 0 0 0 output_no[213]
port 137 nsew signal output
flabel metal2 s 83000 0 83080 80 0 FreeSans 320 0 0 0 output_no[214]
port 138 nsew signal output
flabel metal2 s 83384 0 83464 80 0 FreeSans 320 0 0 0 output_no[215]
port 139 nsew signal output
flabel metal2 s 83768 0 83848 80 0 FreeSans 320 0 0 0 output_no[216]
port 140 nsew signal output
flabel metal2 s 84152 0 84232 80 0 FreeSans 320 0 0 0 output_no[217]
port 141 nsew signal output
flabel metal2 s 84536 0 84616 80 0 FreeSans 320 0 0 0 output_no[218]
port 142 nsew signal output
flabel metal2 s 84920 0 85000 80 0 FreeSans 320 0 0 0 output_no[219]
port 143 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 output_no[21]
port 144 nsew signal output
flabel metal2 s 85304 0 85384 80 0 FreeSans 320 0 0 0 output_no[220]
port 145 nsew signal output
flabel metal2 s 85688 0 85768 80 0 FreeSans 320 0 0 0 output_no[221]
port 146 nsew signal output
flabel metal2 s 86072 0 86152 80 0 FreeSans 320 0 0 0 output_no[222]
port 147 nsew signal output
flabel metal2 s 86456 0 86536 80 0 FreeSans 320 0 0 0 output_no[223]
port 148 nsew signal output
flabel metal2 s 86840 0 86920 80 0 FreeSans 320 0 0 0 output_no[224]
port 149 nsew signal output
flabel metal2 s 87224 0 87304 80 0 FreeSans 320 0 0 0 output_no[225]
port 150 nsew signal output
flabel metal2 s 87608 0 87688 80 0 FreeSans 320 0 0 0 output_no[226]
port 151 nsew signal output
flabel metal2 s 87992 0 88072 80 0 FreeSans 320 0 0 0 output_no[227]
port 152 nsew signal output
flabel metal2 s 88376 0 88456 80 0 FreeSans 320 0 0 0 output_no[228]
port 153 nsew signal output
flabel metal2 s 88760 0 88840 80 0 FreeSans 320 0 0 0 output_no[229]
port 154 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 output_no[22]
port 155 nsew signal output
flabel metal2 s 89144 0 89224 80 0 FreeSans 320 0 0 0 output_no[230]
port 156 nsew signal output
flabel metal2 s 89528 0 89608 80 0 FreeSans 320 0 0 0 output_no[231]
port 157 nsew signal output
flabel metal2 s 89912 0 89992 80 0 FreeSans 320 0 0 0 output_no[232]
port 158 nsew signal output
flabel metal2 s 90296 0 90376 80 0 FreeSans 320 0 0 0 output_no[233]
port 159 nsew signal output
flabel metal2 s 90680 0 90760 80 0 FreeSans 320 0 0 0 output_no[234]
port 160 nsew signal output
flabel metal2 s 91064 0 91144 80 0 FreeSans 320 0 0 0 output_no[235]
port 161 nsew signal output
flabel metal2 s 91448 0 91528 80 0 FreeSans 320 0 0 0 output_no[236]
port 162 nsew signal output
flabel metal2 s 91832 0 91912 80 0 FreeSans 320 0 0 0 output_no[237]
port 163 nsew signal output
flabel metal2 s 92216 0 92296 80 0 FreeSans 320 0 0 0 output_no[238]
port 164 nsew signal output
flabel metal2 s 92600 0 92680 80 0 FreeSans 320 0 0 0 output_no[239]
port 165 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 output_no[23]
port 166 nsew signal output
flabel metal2 s 92984 0 93064 80 0 FreeSans 320 0 0 0 output_no[240]
port 167 nsew signal output
flabel metal2 s 93368 0 93448 80 0 FreeSans 320 0 0 0 output_no[241]
port 168 nsew signal output
flabel metal2 s 93752 0 93832 80 0 FreeSans 320 0 0 0 output_no[242]
port 169 nsew signal output
flabel metal2 s 94136 0 94216 80 0 FreeSans 320 0 0 0 output_no[243]
port 170 nsew signal output
flabel metal2 s 94520 0 94600 80 0 FreeSans 320 0 0 0 output_no[244]
port 171 nsew signal output
flabel metal2 s 94904 0 94984 80 0 FreeSans 320 0 0 0 output_no[245]
port 172 nsew signal output
flabel metal2 s 95288 0 95368 80 0 FreeSans 320 0 0 0 output_no[246]
port 173 nsew signal output
flabel metal2 s 95672 0 95752 80 0 FreeSans 320 0 0 0 output_no[247]
port 174 nsew signal output
flabel metal2 s 96056 0 96136 80 0 FreeSans 320 0 0 0 output_no[248]
port 175 nsew signal output
flabel metal2 s 96440 0 96520 80 0 FreeSans 320 0 0 0 output_no[249]
port 176 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 output_no[24]
port 177 nsew signal output
flabel metal2 s 96824 0 96904 80 0 FreeSans 320 0 0 0 output_no[250]
port 178 nsew signal output
flabel metal2 s 97208 0 97288 80 0 FreeSans 320 0 0 0 output_no[251]
port 179 nsew signal output
flabel metal2 s 97592 0 97672 80 0 FreeSans 320 0 0 0 output_no[252]
port 180 nsew signal output
flabel metal2 s 97976 0 98056 80 0 FreeSans 320 0 0 0 output_no[253]
port 181 nsew signal output
flabel metal2 s 98360 0 98440 80 0 FreeSans 320 0 0 0 output_no[254]
port 182 nsew signal output
flabel metal2 s 98744 0 98824 80 0 FreeSans 320 0 0 0 output_no[255]
port 183 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 output_no[25]
port 184 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 output_no[26]
port 185 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 output_no[27]
port 186 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 output_no[28]
port 187 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 output_no[29]
port 188 nsew signal output
flabel metal2 s 1592 0 1672 80 0 FreeSans 320 0 0 0 output_no[2]
port 189 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 output_no[30]
port 190 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 output_no[31]
port 191 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 output_no[32]
port 192 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 output_no[33]
port 193 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 output_no[34]
port 194 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 output_no[35]
port 195 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 output_no[36]
port 196 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 output_no[37]
port 197 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 output_no[38]
port 198 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 output_no[39]
port 199 nsew signal output
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 output_no[3]
port 200 nsew signal output
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 output_no[40]
port 201 nsew signal output
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 output_no[41]
port 202 nsew signal output
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 output_no[42]
port 203 nsew signal output
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 output_no[43]
port 204 nsew signal output
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 output_no[44]
port 205 nsew signal output
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 output_no[45]
port 206 nsew signal output
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 output_no[46]
port 207 nsew signal output
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 output_no[47]
port 208 nsew signal output
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 output_no[48]
port 209 nsew signal output
flabel metal2 s 19640 0 19720 80 0 FreeSans 320 0 0 0 output_no[49]
port 210 nsew signal output
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 output_no[4]
port 211 nsew signal output
flabel metal2 s 20024 0 20104 80 0 FreeSans 320 0 0 0 output_no[50]
port 212 nsew signal output
flabel metal2 s 20408 0 20488 80 0 FreeSans 320 0 0 0 output_no[51]
port 213 nsew signal output
flabel metal2 s 20792 0 20872 80 0 FreeSans 320 0 0 0 output_no[52]
port 214 nsew signal output
flabel metal2 s 21176 0 21256 80 0 FreeSans 320 0 0 0 output_no[53]
port 215 nsew signal output
flabel metal2 s 21560 0 21640 80 0 FreeSans 320 0 0 0 output_no[54]
port 216 nsew signal output
flabel metal2 s 21944 0 22024 80 0 FreeSans 320 0 0 0 output_no[55]
port 217 nsew signal output
flabel metal2 s 22328 0 22408 80 0 FreeSans 320 0 0 0 output_no[56]
port 218 nsew signal output
flabel metal2 s 22712 0 22792 80 0 FreeSans 320 0 0 0 output_no[57]
port 219 nsew signal output
flabel metal2 s 23096 0 23176 80 0 FreeSans 320 0 0 0 output_no[58]
port 220 nsew signal output
flabel metal2 s 23480 0 23560 80 0 FreeSans 320 0 0 0 output_no[59]
port 221 nsew signal output
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 output_no[5]
port 222 nsew signal output
flabel metal2 s 23864 0 23944 80 0 FreeSans 320 0 0 0 output_no[60]
port 223 nsew signal output
flabel metal2 s 24248 0 24328 80 0 FreeSans 320 0 0 0 output_no[61]
port 224 nsew signal output
flabel metal2 s 24632 0 24712 80 0 FreeSans 320 0 0 0 output_no[62]
port 225 nsew signal output
flabel metal2 s 25016 0 25096 80 0 FreeSans 320 0 0 0 output_no[63]
port 226 nsew signal output
flabel metal2 s 25400 0 25480 80 0 FreeSans 320 0 0 0 output_no[64]
port 227 nsew signal output
flabel metal2 s 25784 0 25864 80 0 FreeSans 320 0 0 0 output_no[65]
port 228 nsew signal output
flabel metal2 s 26168 0 26248 80 0 FreeSans 320 0 0 0 output_no[66]
port 229 nsew signal output
flabel metal2 s 26552 0 26632 80 0 FreeSans 320 0 0 0 output_no[67]
port 230 nsew signal output
flabel metal2 s 26936 0 27016 80 0 FreeSans 320 0 0 0 output_no[68]
port 231 nsew signal output
flabel metal2 s 27320 0 27400 80 0 FreeSans 320 0 0 0 output_no[69]
port 232 nsew signal output
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 output_no[6]
port 233 nsew signal output
flabel metal2 s 27704 0 27784 80 0 FreeSans 320 0 0 0 output_no[70]
port 234 nsew signal output
flabel metal2 s 28088 0 28168 80 0 FreeSans 320 0 0 0 output_no[71]
port 235 nsew signal output
flabel metal2 s 28472 0 28552 80 0 FreeSans 320 0 0 0 output_no[72]
port 236 nsew signal output
flabel metal2 s 28856 0 28936 80 0 FreeSans 320 0 0 0 output_no[73]
port 237 nsew signal output
flabel metal2 s 29240 0 29320 80 0 FreeSans 320 0 0 0 output_no[74]
port 238 nsew signal output
flabel metal2 s 29624 0 29704 80 0 FreeSans 320 0 0 0 output_no[75]
port 239 nsew signal output
flabel metal2 s 30008 0 30088 80 0 FreeSans 320 0 0 0 output_no[76]
port 240 nsew signal output
flabel metal2 s 30392 0 30472 80 0 FreeSans 320 0 0 0 output_no[77]
port 241 nsew signal output
flabel metal2 s 30776 0 30856 80 0 FreeSans 320 0 0 0 output_no[78]
port 242 nsew signal output
flabel metal2 s 31160 0 31240 80 0 FreeSans 320 0 0 0 output_no[79]
port 243 nsew signal output
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 output_no[7]
port 244 nsew signal output
flabel metal2 s 31544 0 31624 80 0 FreeSans 320 0 0 0 output_no[80]
port 245 nsew signal output
flabel metal2 s 31928 0 32008 80 0 FreeSans 320 0 0 0 output_no[81]
port 246 nsew signal output
flabel metal2 s 32312 0 32392 80 0 FreeSans 320 0 0 0 output_no[82]
port 247 nsew signal output
flabel metal2 s 32696 0 32776 80 0 FreeSans 320 0 0 0 output_no[83]
port 248 nsew signal output
flabel metal2 s 33080 0 33160 80 0 FreeSans 320 0 0 0 output_no[84]
port 249 nsew signal output
flabel metal2 s 33464 0 33544 80 0 FreeSans 320 0 0 0 output_no[85]
port 250 nsew signal output
flabel metal2 s 33848 0 33928 80 0 FreeSans 320 0 0 0 output_no[86]
port 251 nsew signal output
flabel metal2 s 34232 0 34312 80 0 FreeSans 320 0 0 0 output_no[87]
port 252 nsew signal output
flabel metal2 s 34616 0 34696 80 0 FreeSans 320 0 0 0 output_no[88]
port 253 nsew signal output
flabel metal2 s 35000 0 35080 80 0 FreeSans 320 0 0 0 output_no[89]
port 254 nsew signal output
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 output_no[8]
port 255 nsew signal output
flabel metal2 s 35384 0 35464 80 0 FreeSans 320 0 0 0 output_no[90]
port 256 nsew signal output
flabel metal2 s 35768 0 35848 80 0 FreeSans 320 0 0 0 output_no[91]
port 257 nsew signal output
flabel metal2 s 36152 0 36232 80 0 FreeSans 320 0 0 0 output_no[92]
port 258 nsew signal output
flabel metal2 s 36536 0 36616 80 0 FreeSans 320 0 0 0 output_no[93]
port 259 nsew signal output
flabel metal2 s 36920 0 37000 80 0 FreeSans 320 0 0 0 output_no[94]
port 260 nsew signal output
flabel metal2 s 37304 0 37384 80 0 FreeSans 320 0 0 0 output_no[95]
port 261 nsew signal output
flabel metal2 s 37688 0 37768 80 0 FreeSans 320 0 0 0 output_no[96]
port 262 nsew signal output
flabel metal2 s 38072 0 38152 80 0 FreeSans 320 0 0 0 output_no[97]
port 263 nsew signal output
flabel metal2 s 38456 0 38536 80 0 FreeSans 320 0 0 0 output_no[98]
port 264 nsew signal output
flabel metal2 s 38840 0 38920 80 0 FreeSans 320 0 0 0 output_no[99]
port 265 nsew signal output
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 output_no[9]
port 266 nsew signal output
flabel metal2 s 1016 0 1096 80 0 FreeSans 320 0 0 0 output_o[0]
port 267 nsew signal output
flabel metal2 s 39416 0 39496 80 0 FreeSans 320 0 0 0 output_o[100]
port 268 nsew signal output
flabel metal2 s 39800 0 39880 80 0 FreeSans 320 0 0 0 output_o[101]
port 269 nsew signal output
flabel metal2 s 40184 0 40264 80 0 FreeSans 320 0 0 0 output_o[102]
port 270 nsew signal output
flabel metal2 s 40568 0 40648 80 0 FreeSans 320 0 0 0 output_o[103]
port 271 nsew signal output
flabel metal2 s 40952 0 41032 80 0 FreeSans 320 0 0 0 output_o[104]
port 272 nsew signal output
flabel metal2 s 41336 0 41416 80 0 FreeSans 320 0 0 0 output_o[105]
port 273 nsew signal output
flabel metal2 s 41720 0 41800 80 0 FreeSans 320 0 0 0 output_o[106]
port 274 nsew signal output
flabel metal2 s 42104 0 42184 80 0 FreeSans 320 0 0 0 output_o[107]
port 275 nsew signal output
flabel metal2 s 42488 0 42568 80 0 FreeSans 320 0 0 0 output_o[108]
port 276 nsew signal output
flabel metal2 s 42872 0 42952 80 0 FreeSans 320 0 0 0 output_o[109]
port 277 nsew signal output
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 output_o[10]
port 278 nsew signal output
flabel metal2 s 43256 0 43336 80 0 FreeSans 320 0 0 0 output_o[110]
port 279 nsew signal output
flabel metal2 s 43640 0 43720 80 0 FreeSans 320 0 0 0 output_o[111]
port 280 nsew signal output
flabel metal2 s 44024 0 44104 80 0 FreeSans 320 0 0 0 output_o[112]
port 281 nsew signal output
flabel metal2 s 44408 0 44488 80 0 FreeSans 320 0 0 0 output_o[113]
port 282 nsew signal output
flabel metal2 s 44792 0 44872 80 0 FreeSans 320 0 0 0 output_o[114]
port 283 nsew signal output
flabel metal2 s 45176 0 45256 80 0 FreeSans 320 0 0 0 output_o[115]
port 284 nsew signal output
flabel metal2 s 45560 0 45640 80 0 FreeSans 320 0 0 0 output_o[116]
port 285 nsew signal output
flabel metal2 s 45944 0 46024 80 0 FreeSans 320 0 0 0 output_o[117]
port 286 nsew signal output
flabel metal2 s 46328 0 46408 80 0 FreeSans 320 0 0 0 output_o[118]
port 287 nsew signal output
flabel metal2 s 46712 0 46792 80 0 FreeSans 320 0 0 0 output_o[119]
port 288 nsew signal output
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 output_o[11]
port 289 nsew signal output
flabel metal2 s 47096 0 47176 80 0 FreeSans 320 0 0 0 output_o[120]
port 290 nsew signal output
flabel metal2 s 47480 0 47560 80 0 FreeSans 320 0 0 0 output_o[121]
port 291 nsew signal output
flabel metal2 s 47864 0 47944 80 0 FreeSans 320 0 0 0 output_o[122]
port 292 nsew signal output
flabel metal2 s 48248 0 48328 80 0 FreeSans 320 0 0 0 output_o[123]
port 293 nsew signal output
flabel metal2 s 48632 0 48712 80 0 FreeSans 320 0 0 0 output_o[124]
port 294 nsew signal output
flabel metal2 s 49016 0 49096 80 0 FreeSans 320 0 0 0 output_o[125]
port 295 nsew signal output
flabel metal2 s 49400 0 49480 80 0 FreeSans 320 0 0 0 output_o[126]
port 296 nsew signal output
flabel metal2 s 49784 0 49864 80 0 FreeSans 320 0 0 0 output_o[127]
port 297 nsew signal output
flabel metal2 s 50168 0 50248 80 0 FreeSans 320 0 0 0 output_o[128]
port 298 nsew signal output
flabel metal2 s 50552 0 50632 80 0 FreeSans 320 0 0 0 output_o[129]
port 299 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 output_o[12]
port 300 nsew signal output
flabel metal2 s 50936 0 51016 80 0 FreeSans 320 0 0 0 output_o[130]
port 301 nsew signal output
flabel metal2 s 51320 0 51400 80 0 FreeSans 320 0 0 0 output_o[131]
port 302 nsew signal output
flabel metal2 s 51704 0 51784 80 0 FreeSans 320 0 0 0 output_o[132]
port 303 nsew signal output
flabel metal2 s 52088 0 52168 80 0 FreeSans 320 0 0 0 output_o[133]
port 304 nsew signal output
flabel metal2 s 52472 0 52552 80 0 FreeSans 320 0 0 0 output_o[134]
port 305 nsew signal output
flabel metal2 s 52856 0 52936 80 0 FreeSans 320 0 0 0 output_o[135]
port 306 nsew signal output
flabel metal2 s 53240 0 53320 80 0 FreeSans 320 0 0 0 output_o[136]
port 307 nsew signal output
flabel metal2 s 53624 0 53704 80 0 FreeSans 320 0 0 0 output_o[137]
port 308 nsew signal output
flabel metal2 s 54008 0 54088 80 0 FreeSans 320 0 0 0 output_o[138]
port 309 nsew signal output
flabel metal2 s 54392 0 54472 80 0 FreeSans 320 0 0 0 output_o[139]
port 310 nsew signal output
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 output_o[13]
port 311 nsew signal output
flabel metal2 s 54776 0 54856 80 0 FreeSans 320 0 0 0 output_o[140]
port 312 nsew signal output
flabel metal2 s 55160 0 55240 80 0 FreeSans 320 0 0 0 output_o[141]
port 313 nsew signal output
flabel metal2 s 55544 0 55624 80 0 FreeSans 320 0 0 0 output_o[142]
port 314 nsew signal output
flabel metal2 s 55928 0 56008 80 0 FreeSans 320 0 0 0 output_o[143]
port 315 nsew signal output
flabel metal2 s 56312 0 56392 80 0 FreeSans 320 0 0 0 output_o[144]
port 316 nsew signal output
flabel metal2 s 56696 0 56776 80 0 FreeSans 320 0 0 0 output_o[145]
port 317 nsew signal output
flabel metal2 s 57080 0 57160 80 0 FreeSans 320 0 0 0 output_o[146]
port 318 nsew signal output
flabel metal2 s 57464 0 57544 80 0 FreeSans 320 0 0 0 output_o[147]
port 319 nsew signal output
flabel metal2 s 57848 0 57928 80 0 FreeSans 320 0 0 0 output_o[148]
port 320 nsew signal output
flabel metal2 s 58232 0 58312 80 0 FreeSans 320 0 0 0 output_o[149]
port 321 nsew signal output
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 output_o[14]
port 322 nsew signal output
flabel metal2 s 58616 0 58696 80 0 FreeSans 320 0 0 0 output_o[150]
port 323 nsew signal output
flabel metal2 s 59000 0 59080 80 0 FreeSans 320 0 0 0 output_o[151]
port 324 nsew signal output
flabel metal2 s 59384 0 59464 80 0 FreeSans 320 0 0 0 output_o[152]
port 325 nsew signal output
flabel metal2 s 59768 0 59848 80 0 FreeSans 320 0 0 0 output_o[153]
port 326 nsew signal output
flabel metal2 s 60152 0 60232 80 0 FreeSans 320 0 0 0 output_o[154]
port 327 nsew signal output
flabel metal2 s 60536 0 60616 80 0 FreeSans 320 0 0 0 output_o[155]
port 328 nsew signal output
flabel metal2 s 60920 0 61000 80 0 FreeSans 320 0 0 0 output_o[156]
port 329 nsew signal output
flabel metal2 s 61304 0 61384 80 0 FreeSans 320 0 0 0 output_o[157]
port 330 nsew signal output
flabel metal2 s 61688 0 61768 80 0 FreeSans 320 0 0 0 output_o[158]
port 331 nsew signal output
flabel metal2 s 62072 0 62152 80 0 FreeSans 320 0 0 0 output_o[159]
port 332 nsew signal output
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 output_o[15]
port 333 nsew signal output
flabel metal2 s 62456 0 62536 80 0 FreeSans 320 0 0 0 output_o[160]
port 334 nsew signal output
flabel metal2 s 62840 0 62920 80 0 FreeSans 320 0 0 0 output_o[161]
port 335 nsew signal output
flabel metal2 s 63224 0 63304 80 0 FreeSans 320 0 0 0 output_o[162]
port 336 nsew signal output
flabel metal2 s 63608 0 63688 80 0 FreeSans 320 0 0 0 output_o[163]
port 337 nsew signal output
flabel metal2 s 63992 0 64072 80 0 FreeSans 320 0 0 0 output_o[164]
port 338 nsew signal output
flabel metal2 s 64376 0 64456 80 0 FreeSans 320 0 0 0 output_o[165]
port 339 nsew signal output
flabel metal2 s 64760 0 64840 80 0 FreeSans 320 0 0 0 output_o[166]
port 340 nsew signal output
flabel metal2 s 65144 0 65224 80 0 FreeSans 320 0 0 0 output_o[167]
port 341 nsew signal output
flabel metal2 s 65528 0 65608 80 0 FreeSans 320 0 0 0 output_o[168]
port 342 nsew signal output
flabel metal2 s 65912 0 65992 80 0 FreeSans 320 0 0 0 output_o[169]
port 343 nsew signal output
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 output_o[16]
port 344 nsew signal output
flabel metal2 s 66296 0 66376 80 0 FreeSans 320 0 0 0 output_o[170]
port 345 nsew signal output
flabel metal2 s 66680 0 66760 80 0 FreeSans 320 0 0 0 output_o[171]
port 346 nsew signal output
flabel metal2 s 67064 0 67144 80 0 FreeSans 320 0 0 0 output_o[172]
port 347 nsew signal output
flabel metal2 s 67448 0 67528 80 0 FreeSans 320 0 0 0 output_o[173]
port 348 nsew signal output
flabel metal2 s 67832 0 67912 80 0 FreeSans 320 0 0 0 output_o[174]
port 349 nsew signal output
flabel metal2 s 68216 0 68296 80 0 FreeSans 320 0 0 0 output_o[175]
port 350 nsew signal output
flabel metal2 s 68600 0 68680 80 0 FreeSans 320 0 0 0 output_o[176]
port 351 nsew signal output
flabel metal2 s 68984 0 69064 80 0 FreeSans 320 0 0 0 output_o[177]
port 352 nsew signal output
flabel metal2 s 69368 0 69448 80 0 FreeSans 320 0 0 0 output_o[178]
port 353 nsew signal output
flabel metal2 s 69752 0 69832 80 0 FreeSans 320 0 0 0 output_o[179]
port 354 nsew signal output
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 output_o[17]
port 355 nsew signal output
flabel metal2 s 70136 0 70216 80 0 FreeSans 320 0 0 0 output_o[180]
port 356 nsew signal output
flabel metal2 s 70520 0 70600 80 0 FreeSans 320 0 0 0 output_o[181]
port 357 nsew signal output
flabel metal2 s 70904 0 70984 80 0 FreeSans 320 0 0 0 output_o[182]
port 358 nsew signal output
flabel metal2 s 71288 0 71368 80 0 FreeSans 320 0 0 0 output_o[183]
port 359 nsew signal output
flabel metal2 s 71672 0 71752 80 0 FreeSans 320 0 0 0 output_o[184]
port 360 nsew signal output
flabel metal2 s 72056 0 72136 80 0 FreeSans 320 0 0 0 output_o[185]
port 361 nsew signal output
flabel metal2 s 72440 0 72520 80 0 FreeSans 320 0 0 0 output_o[186]
port 362 nsew signal output
flabel metal2 s 72824 0 72904 80 0 FreeSans 320 0 0 0 output_o[187]
port 363 nsew signal output
flabel metal2 s 73208 0 73288 80 0 FreeSans 320 0 0 0 output_o[188]
port 364 nsew signal output
flabel metal2 s 73592 0 73672 80 0 FreeSans 320 0 0 0 output_o[189]
port 365 nsew signal output
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 output_o[18]
port 366 nsew signal output
flabel metal2 s 73976 0 74056 80 0 FreeSans 320 0 0 0 output_o[190]
port 367 nsew signal output
flabel metal2 s 74360 0 74440 80 0 FreeSans 320 0 0 0 output_o[191]
port 368 nsew signal output
flabel metal2 s 74744 0 74824 80 0 FreeSans 320 0 0 0 output_o[192]
port 369 nsew signal output
flabel metal2 s 75128 0 75208 80 0 FreeSans 320 0 0 0 output_o[193]
port 370 nsew signal output
flabel metal2 s 75512 0 75592 80 0 FreeSans 320 0 0 0 output_o[194]
port 371 nsew signal output
flabel metal2 s 75896 0 75976 80 0 FreeSans 320 0 0 0 output_o[195]
port 372 nsew signal output
flabel metal2 s 76280 0 76360 80 0 FreeSans 320 0 0 0 output_o[196]
port 373 nsew signal output
flabel metal2 s 76664 0 76744 80 0 FreeSans 320 0 0 0 output_o[197]
port 374 nsew signal output
flabel metal2 s 77048 0 77128 80 0 FreeSans 320 0 0 0 output_o[198]
port 375 nsew signal output
flabel metal2 s 77432 0 77512 80 0 FreeSans 320 0 0 0 output_o[199]
port 376 nsew signal output
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 output_o[19]
port 377 nsew signal output
flabel metal2 s 1400 0 1480 80 0 FreeSans 320 0 0 0 output_o[1]
port 378 nsew signal output
flabel metal2 s 77816 0 77896 80 0 FreeSans 320 0 0 0 output_o[200]
port 379 nsew signal output
flabel metal2 s 78200 0 78280 80 0 FreeSans 320 0 0 0 output_o[201]
port 380 nsew signal output
flabel metal2 s 78584 0 78664 80 0 FreeSans 320 0 0 0 output_o[202]
port 381 nsew signal output
flabel metal2 s 78968 0 79048 80 0 FreeSans 320 0 0 0 output_o[203]
port 382 nsew signal output
flabel metal2 s 79352 0 79432 80 0 FreeSans 320 0 0 0 output_o[204]
port 383 nsew signal output
flabel metal2 s 79736 0 79816 80 0 FreeSans 320 0 0 0 output_o[205]
port 384 nsew signal output
flabel metal2 s 80120 0 80200 80 0 FreeSans 320 0 0 0 output_o[206]
port 385 nsew signal output
flabel metal2 s 80504 0 80584 80 0 FreeSans 320 0 0 0 output_o[207]
port 386 nsew signal output
flabel metal2 s 80888 0 80968 80 0 FreeSans 320 0 0 0 output_o[208]
port 387 nsew signal output
flabel metal2 s 81272 0 81352 80 0 FreeSans 320 0 0 0 output_o[209]
port 388 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 output_o[20]
port 389 nsew signal output
flabel metal2 s 81656 0 81736 80 0 FreeSans 320 0 0 0 output_o[210]
port 390 nsew signal output
flabel metal2 s 82040 0 82120 80 0 FreeSans 320 0 0 0 output_o[211]
port 391 nsew signal output
flabel metal2 s 82424 0 82504 80 0 FreeSans 320 0 0 0 output_o[212]
port 392 nsew signal output
flabel metal2 s 82808 0 82888 80 0 FreeSans 320 0 0 0 output_o[213]
port 393 nsew signal output
flabel metal2 s 83192 0 83272 80 0 FreeSans 320 0 0 0 output_o[214]
port 394 nsew signal output
flabel metal2 s 83576 0 83656 80 0 FreeSans 320 0 0 0 output_o[215]
port 395 nsew signal output
flabel metal2 s 83960 0 84040 80 0 FreeSans 320 0 0 0 output_o[216]
port 396 nsew signal output
flabel metal2 s 84344 0 84424 80 0 FreeSans 320 0 0 0 output_o[217]
port 397 nsew signal output
flabel metal2 s 84728 0 84808 80 0 FreeSans 320 0 0 0 output_o[218]
port 398 nsew signal output
flabel metal2 s 85112 0 85192 80 0 FreeSans 320 0 0 0 output_o[219]
port 399 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 output_o[21]
port 400 nsew signal output
flabel metal2 s 85496 0 85576 80 0 FreeSans 320 0 0 0 output_o[220]
port 401 nsew signal output
flabel metal2 s 85880 0 85960 80 0 FreeSans 320 0 0 0 output_o[221]
port 402 nsew signal output
flabel metal2 s 86264 0 86344 80 0 FreeSans 320 0 0 0 output_o[222]
port 403 nsew signal output
flabel metal2 s 86648 0 86728 80 0 FreeSans 320 0 0 0 output_o[223]
port 404 nsew signal output
flabel metal2 s 87032 0 87112 80 0 FreeSans 320 0 0 0 output_o[224]
port 405 nsew signal output
flabel metal2 s 87416 0 87496 80 0 FreeSans 320 0 0 0 output_o[225]
port 406 nsew signal output
flabel metal2 s 87800 0 87880 80 0 FreeSans 320 0 0 0 output_o[226]
port 407 nsew signal output
flabel metal2 s 88184 0 88264 80 0 FreeSans 320 0 0 0 output_o[227]
port 408 nsew signal output
flabel metal2 s 88568 0 88648 80 0 FreeSans 320 0 0 0 output_o[228]
port 409 nsew signal output
flabel metal2 s 88952 0 89032 80 0 FreeSans 320 0 0 0 output_o[229]
port 410 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 output_o[22]
port 411 nsew signal output
flabel metal2 s 89336 0 89416 80 0 FreeSans 320 0 0 0 output_o[230]
port 412 nsew signal output
flabel metal2 s 89720 0 89800 80 0 FreeSans 320 0 0 0 output_o[231]
port 413 nsew signal output
flabel metal2 s 90104 0 90184 80 0 FreeSans 320 0 0 0 output_o[232]
port 414 nsew signal output
flabel metal2 s 90488 0 90568 80 0 FreeSans 320 0 0 0 output_o[233]
port 415 nsew signal output
flabel metal2 s 90872 0 90952 80 0 FreeSans 320 0 0 0 output_o[234]
port 416 nsew signal output
flabel metal2 s 91256 0 91336 80 0 FreeSans 320 0 0 0 output_o[235]
port 417 nsew signal output
flabel metal2 s 91640 0 91720 80 0 FreeSans 320 0 0 0 output_o[236]
port 418 nsew signal output
flabel metal2 s 92024 0 92104 80 0 FreeSans 320 0 0 0 output_o[237]
port 419 nsew signal output
flabel metal2 s 92408 0 92488 80 0 FreeSans 320 0 0 0 output_o[238]
port 420 nsew signal output
flabel metal2 s 92792 0 92872 80 0 FreeSans 320 0 0 0 output_o[239]
port 421 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 output_o[23]
port 422 nsew signal output
flabel metal2 s 93176 0 93256 80 0 FreeSans 320 0 0 0 output_o[240]
port 423 nsew signal output
flabel metal2 s 93560 0 93640 80 0 FreeSans 320 0 0 0 output_o[241]
port 424 nsew signal output
flabel metal2 s 93944 0 94024 80 0 FreeSans 320 0 0 0 output_o[242]
port 425 nsew signal output
flabel metal2 s 94328 0 94408 80 0 FreeSans 320 0 0 0 output_o[243]
port 426 nsew signal output
flabel metal2 s 94712 0 94792 80 0 FreeSans 320 0 0 0 output_o[244]
port 427 nsew signal output
flabel metal2 s 95096 0 95176 80 0 FreeSans 320 0 0 0 output_o[245]
port 428 nsew signal output
flabel metal2 s 95480 0 95560 80 0 FreeSans 320 0 0 0 output_o[246]
port 429 nsew signal output
flabel metal2 s 95864 0 95944 80 0 FreeSans 320 0 0 0 output_o[247]
port 430 nsew signal output
flabel metal2 s 96248 0 96328 80 0 FreeSans 320 0 0 0 output_o[248]
port 431 nsew signal output
flabel metal2 s 96632 0 96712 80 0 FreeSans 320 0 0 0 output_o[249]
port 432 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 output_o[24]
port 433 nsew signal output
flabel metal2 s 97016 0 97096 80 0 FreeSans 320 0 0 0 output_o[250]
port 434 nsew signal output
flabel metal2 s 97400 0 97480 80 0 FreeSans 320 0 0 0 output_o[251]
port 435 nsew signal output
flabel metal2 s 97784 0 97864 80 0 FreeSans 320 0 0 0 output_o[252]
port 436 nsew signal output
flabel metal2 s 98168 0 98248 80 0 FreeSans 320 0 0 0 output_o[253]
port 437 nsew signal output
flabel metal2 s 98552 0 98632 80 0 FreeSans 320 0 0 0 output_o[254]
port 438 nsew signal output
flabel metal2 s 98936 0 99016 80 0 FreeSans 320 0 0 0 output_o[255]
port 439 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 output_o[25]
port 440 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 output_o[26]
port 441 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 output_o[27]
port 442 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 output_o[28]
port 443 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 output_o[29]
port 444 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 output_o[2]
port 445 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 output_o[30]
port 446 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 output_o[31]
port 447 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 output_o[32]
port 448 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 output_o[33]
port 449 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 output_o[34]
port 450 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 output_o[35]
port 451 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 output_o[36]
port 452 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 output_o[37]
port 453 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 output_o[38]
port 454 nsew signal output
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 output_o[39]
port 455 nsew signal output
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 output_o[3]
port 456 nsew signal output
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 output_o[40]
port 457 nsew signal output
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 output_o[41]
port 458 nsew signal output
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 output_o[42]
port 459 nsew signal output
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 output_o[43]
port 460 nsew signal output
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 output_o[44]
port 461 nsew signal output
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 output_o[45]
port 462 nsew signal output
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 output_o[46]
port 463 nsew signal output
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 output_o[47]
port 464 nsew signal output
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 output_o[48]
port 465 nsew signal output
flabel metal2 s 19832 0 19912 80 0 FreeSans 320 0 0 0 output_o[49]
port 466 nsew signal output
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 output_o[4]
port 467 nsew signal output
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 output_o[50]
port 468 nsew signal output
flabel metal2 s 20600 0 20680 80 0 FreeSans 320 0 0 0 output_o[51]
port 469 nsew signal output
flabel metal2 s 20984 0 21064 80 0 FreeSans 320 0 0 0 output_o[52]
port 470 nsew signal output
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 output_o[53]
port 471 nsew signal output
flabel metal2 s 21752 0 21832 80 0 FreeSans 320 0 0 0 output_o[54]
port 472 nsew signal output
flabel metal2 s 22136 0 22216 80 0 FreeSans 320 0 0 0 output_o[55]
port 473 nsew signal output
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 output_o[56]
port 474 nsew signal output
flabel metal2 s 22904 0 22984 80 0 FreeSans 320 0 0 0 output_o[57]
port 475 nsew signal output
flabel metal2 s 23288 0 23368 80 0 FreeSans 320 0 0 0 output_o[58]
port 476 nsew signal output
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 output_o[59]
port 477 nsew signal output
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 output_o[5]
port 478 nsew signal output
flabel metal2 s 24056 0 24136 80 0 FreeSans 320 0 0 0 output_o[60]
port 479 nsew signal output
flabel metal2 s 24440 0 24520 80 0 FreeSans 320 0 0 0 output_o[61]
port 480 nsew signal output
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 output_o[62]
port 481 nsew signal output
flabel metal2 s 25208 0 25288 80 0 FreeSans 320 0 0 0 output_o[63]
port 482 nsew signal output
flabel metal2 s 25592 0 25672 80 0 FreeSans 320 0 0 0 output_o[64]
port 483 nsew signal output
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 output_o[65]
port 484 nsew signal output
flabel metal2 s 26360 0 26440 80 0 FreeSans 320 0 0 0 output_o[66]
port 485 nsew signal output
flabel metal2 s 26744 0 26824 80 0 FreeSans 320 0 0 0 output_o[67]
port 486 nsew signal output
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 output_o[68]
port 487 nsew signal output
flabel metal2 s 27512 0 27592 80 0 FreeSans 320 0 0 0 output_o[69]
port 488 nsew signal output
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 output_o[6]
port 489 nsew signal output
flabel metal2 s 27896 0 27976 80 0 FreeSans 320 0 0 0 output_o[70]
port 490 nsew signal output
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 output_o[71]
port 491 nsew signal output
flabel metal2 s 28664 0 28744 80 0 FreeSans 320 0 0 0 output_o[72]
port 492 nsew signal output
flabel metal2 s 29048 0 29128 80 0 FreeSans 320 0 0 0 output_o[73]
port 493 nsew signal output
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 output_o[74]
port 494 nsew signal output
flabel metal2 s 29816 0 29896 80 0 FreeSans 320 0 0 0 output_o[75]
port 495 nsew signal output
flabel metal2 s 30200 0 30280 80 0 FreeSans 320 0 0 0 output_o[76]
port 496 nsew signal output
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 output_o[77]
port 497 nsew signal output
flabel metal2 s 30968 0 31048 80 0 FreeSans 320 0 0 0 output_o[78]
port 498 nsew signal output
flabel metal2 s 31352 0 31432 80 0 FreeSans 320 0 0 0 output_o[79]
port 499 nsew signal output
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 output_o[7]
port 500 nsew signal output
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 output_o[80]
port 501 nsew signal output
flabel metal2 s 32120 0 32200 80 0 FreeSans 320 0 0 0 output_o[81]
port 502 nsew signal output
flabel metal2 s 32504 0 32584 80 0 FreeSans 320 0 0 0 output_o[82]
port 503 nsew signal output
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 output_o[83]
port 504 nsew signal output
flabel metal2 s 33272 0 33352 80 0 FreeSans 320 0 0 0 output_o[84]
port 505 nsew signal output
flabel metal2 s 33656 0 33736 80 0 FreeSans 320 0 0 0 output_o[85]
port 506 nsew signal output
flabel metal2 s 34040 0 34120 80 0 FreeSans 320 0 0 0 output_o[86]
port 507 nsew signal output
flabel metal2 s 34424 0 34504 80 0 FreeSans 320 0 0 0 output_o[87]
port 508 nsew signal output
flabel metal2 s 34808 0 34888 80 0 FreeSans 320 0 0 0 output_o[88]
port 509 nsew signal output
flabel metal2 s 35192 0 35272 80 0 FreeSans 320 0 0 0 output_o[89]
port 510 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 output_o[8]
port 511 nsew signal output
flabel metal2 s 35576 0 35656 80 0 FreeSans 320 0 0 0 output_o[90]
port 512 nsew signal output
flabel metal2 s 35960 0 36040 80 0 FreeSans 320 0 0 0 output_o[91]
port 513 nsew signal output
flabel metal2 s 36344 0 36424 80 0 FreeSans 320 0 0 0 output_o[92]
port 514 nsew signal output
flabel metal2 s 36728 0 36808 80 0 FreeSans 320 0 0 0 output_o[93]
port 515 nsew signal output
flabel metal2 s 37112 0 37192 80 0 FreeSans 320 0 0 0 output_o[94]
port 516 nsew signal output
flabel metal2 s 37496 0 37576 80 0 FreeSans 320 0 0 0 output_o[95]
port 517 nsew signal output
flabel metal2 s 37880 0 37960 80 0 FreeSans 320 0 0 0 output_o[96]
port 518 nsew signal output
flabel metal2 s 38264 0 38344 80 0 FreeSans 320 0 0 0 output_o[97]
port 519 nsew signal output
flabel metal2 s 38648 0 38728 80 0 FreeSans 320 0 0 0 output_o[98]
port 520 nsew signal output
flabel metal2 s 39032 0 39112 80 0 FreeSans 320 0 0 0 output_o[99]
port 521 nsew signal output
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 output_o[9]
port 522 nsew signal output
rlabel via1 49968 8316 49968 8316 0 VGND
rlabel metal1 49968 9072 49968 9072 0 VPWR
rlabel metal3 47232 3444 47232 3444 0 _000_
rlabel metal2 43776 1176 43776 1176 0 _001_
rlabel via2 5760 3024 5760 3024 0 _002_
rlabel metal2 6816 1974 6816 1974 0 _003_
rlabel metal3 35040 4116 35040 4116 0 _004_
rlabel metal2 49536 5292 49536 5292 0 _005_
rlabel metal2 53280 3486 53280 3486 0 _006_
rlabel metal2 56448 5880 56448 5880 0 _007_
rlabel metal2 68928 4032 68928 4032 0 _008_
rlabel metal3 59184 5628 59184 5628 0 _009_
rlabel metal2 55392 4788 55392 4788 0 _010_
rlabel metal2 48288 5586 48288 5586 0 _011_
rlabel metal2 46656 4578 46656 4578 0 _012_
rlabel metal2 50688 4830 50688 4830 0 _013_
rlabel metal2 32928 3990 32928 3990 0 _014_
rlabel metal3 61488 5040 61488 5040 0 _015_
rlabel metal2 62016 2646 62016 2646 0 _016_
rlabel metal2 48096 4662 48096 4662 0 _017_
rlabel metal2 50304 3402 50304 3402 0 _018_
rlabel metal3 50160 4116 50160 4116 0 _019_
rlabel metal3 50784 1260 50784 1260 0 _020_
rlabel metal2 57216 1890 57216 1890 0 _021_
rlabel metal2 47616 5922 47616 5922 0 _022_
rlabel metal2 57456 1764 57456 1764 0 _023_
rlabel metal2 52560 1092 52560 1092 0 _024_
rlabel metal2 58176 5334 58176 5334 0 _025_
rlabel metal2 52944 1764 52944 1764 0 _026_
rlabel metal2 48768 5166 48768 5166 0 _027_
rlabel metal2 53664 4200 53664 4200 0 _028_
rlabel metal2 59328 1008 59328 1008 0 _029_
rlabel metal2 55104 1344 55104 1344 0 _030_
rlabel via1 54624 1247 54624 1247 0 _031_
rlabel metal3 60672 4788 60672 4788 0 _032_
rlabel via2 55296 2759 55296 2759 0 _033_
rlabel metal2 61824 2688 61824 2688 0 _034_
rlabel metal2 37344 4242 37344 4242 0 _035_
rlabel metal3 67008 3444 67008 3444 0 _036_
rlabel metal2 67104 2352 67104 2352 0 _037_
rlabel metal2 68640 3486 68640 3486 0 _038_
rlabel metal4 54816 1470 54816 1470 0 _039_
rlabel metal2 1632 2856 1632 2856 0 _040_
rlabel metal4 1632 840 1632 840 0 _041_
rlabel metal3 2112 3486 2112 3486 0 _042_
rlabel metal2 13728 924 13728 924 0 _043_
rlabel metal5 3520 2646 3520 2646 0 _044_
rlabel metal3 49152 588 49152 588 0 _045_
rlabel metal2 2688 2940 2688 2940 0 _046_
rlabel metal4 50208 756 50208 756 0 _047_
rlabel metal2 3168 2688 3168 2688 0 _048_
rlabel metal2 14880 1134 14880 1134 0 _049_
rlabel metal3 3552 2646 3552 2646 0 _050_
rlabel metal2 15264 882 15264 882 0 _051_
rlabel metal2 33792 3024 33792 3024 0 _052_
rlabel metal2 15648 1050 15648 1050 0 _053_
rlabel metal2 4416 3528 4416 3528 0 _054_
rlabel metal2 46656 1050 46656 1050 0 _055_
rlabel metal2 4896 3318 4896 3318 0 _056_
rlabel metal2 51168 1596 51168 1596 0 _057_
rlabel metal3 5184 3402 5184 3402 0 _058_
rlabel metal2 16800 1182 16800 1182 0 _059_
rlabel metal2 35328 3234 35328 3234 0 _060_
rlabel metal3 47760 1092 47760 1092 0 _061_
rlabel metal2 35712 3612 35712 3612 0 _062_
rlabel metal2 48192 1134 48192 1134 0 _063_
rlabel metal2 36096 3234 36096 3234 0 _064_
rlabel metal2 53568 336 53568 336 0 _065_
rlabel metal2 92256 3192 92256 3192 0 _066_
rlabel metal4 48960 1050 48960 1050 0 _067_
rlabel metal4 36864 3066 36864 3066 0 _068_
rlabel metal2 49536 1176 49536 1176 0 _069_
rlabel metal2 37728 4158 37728 4158 0 _070_
rlabel metal2 68784 3444 68784 3444 0 _071_
rlabel metal2 68976 3612 68976 3612 0 _072_
rlabel metal3 91824 4116 91824 4116 0 _073_
rlabel metal2 75120 3444 75120 3444 0 _074_
rlabel metal2 74976 1260 74976 1260 0 _075_
rlabel metal2 85920 2646 85920 2646 0 _076_
rlabel metal2 82080 1134 82080 1134 0 _077_
rlabel metal2 87072 3528 87072 3528 0 _078_
rlabel metal2 87216 1092 87216 1092 0 _079_
rlabel metal2 93504 3528 93504 3528 0 _080_
rlabel metal2 93504 2772 93504 2772 0 _081_
rlabel metal2 11328 3528 11328 3528 0 _082_
rlabel metal2 12384 1134 12384 1134 0 _083_
rlabel metal2 18144 3738 18144 3738 0 _084_
rlabel metal3 19056 1092 19056 1092 0 _085_
rlabel metal3 19824 1932 19824 1932 0 _086_
rlabel metal2 25056 1596 25056 1596 0 _087_
rlabel metal2 7008 4200 7008 4200 0 _088_
rlabel metal3 30240 2604 30240 2604 0 _089_
rlabel metal2 29184 1134 29184 1134 0 _090_
rlabel metal3 33024 3444 33024 3444 0 _091_
rlabel metal2 35520 1134 35520 1134 0 _092_
rlabel metal2 37536 3738 37536 3738 0 _093_
rlabel metal2 37920 2142 37920 2142 0 _094_
rlabel metal2 6240 8456 6240 8456 0 ena_i
rlabel metal2 17184 8414 17184 8414 0 input_ni[0]
rlabel metal2 28128 8456 28128 8456 0 input_ni[1]
rlabel metal2 46752 6468 46752 6468 0 input_ni[2]
rlabel metal2 49440 8214 49440 8214 0 input_ni[3]
rlabel metal2 61056 5544 61056 5544 0 input_ni[4]
rlabel metal2 71904 7784 71904 7784 0 input_ni[5]
rlabel metal4 66816 4242 66816 4242 0 input_ni[6]
rlabel metal3 37248 3990 37248 3990 0 input_ni[7]
rlabel metal2 864 618 864 618 0 output_no[0]
rlabel metal2 39264 492 39264 492 0 output_no[100]
rlabel metal2 39648 492 39648 492 0 output_no[101]
rlabel metal2 40032 492 40032 492 0 output_no[102]
rlabel metal2 40224 1344 40224 1344 0 output_no[103]
rlabel metal2 40800 492 40800 492 0 output_no[104]
rlabel metal2 41184 492 41184 492 0 output_no[105]
rlabel metal2 41568 450 41568 450 0 output_no[106]
rlabel metal2 41952 324 41952 324 0 output_no[107]
rlabel metal2 42192 1344 42192 1344 0 output_no[108]
rlabel metal2 42720 492 42720 492 0 output_no[109]
rlabel metal2 4704 198 4704 198 0 output_no[10]
rlabel metal2 43104 492 43104 492 0 output_no[110]
rlabel metal3 43200 2016 43200 2016 0 output_no[111]
rlabel metal2 43872 870 43872 870 0 output_no[112]
rlabel metal2 44208 1260 44208 1260 0 output_no[113]
rlabel metal2 44640 1290 44640 1290 0 output_no[114]
rlabel metal2 44976 1260 44976 1260 0 output_no[115]
rlabel metal2 45408 660 45408 660 0 output_no[116]
rlabel metal2 45792 828 45792 828 0 output_no[117]
rlabel metal2 46176 1290 46176 1290 0 output_no[118]
rlabel metal2 46512 1260 46512 1260 0 output_no[119]
rlabel metal2 5088 114 5088 114 0 output_no[11]
rlabel metal2 46944 1626 46944 1626 0 output_no[120]
rlabel metal2 47328 1626 47328 1626 0 output_no[121]
rlabel metal2 47712 1626 47712 1626 0 output_no[122]
rlabel metal2 48096 660 48096 660 0 output_no[123]
rlabel metal2 48480 660 48480 660 0 output_no[124]
rlabel metal2 48864 660 48864 660 0 output_no[125]
rlabel metal2 49248 870 49248 870 0 output_no[126]
rlabel metal2 49632 912 49632 912 0 output_no[127]
rlabel metal2 50016 324 50016 324 0 output_no[128]
rlabel metal2 50400 492 50400 492 0 output_no[129]
rlabel metal2 5472 408 5472 408 0 output_no[12]
rlabel metal2 50784 492 50784 492 0 output_no[130]
rlabel metal2 51168 492 51168 492 0 output_no[131]
rlabel metal2 51552 870 51552 870 0 output_no[132]
rlabel metal2 51936 492 51936 492 0 output_no[133]
rlabel metal2 52320 912 52320 912 0 output_no[134]
rlabel metal2 52704 450 52704 450 0 output_no[135]
rlabel metal2 53088 786 53088 786 0 output_no[136]
rlabel metal2 53472 492 53472 492 0 output_no[137]
rlabel metal2 53856 282 53856 282 0 output_no[138]
rlabel metal2 54240 492 54240 492 0 output_no[139]
rlabel metal2 6240 1932 6240 1932 0 output_no[13]
rlabel metal2 54624 534 54624 534 0 output_no[140]
rlabel metal2 55008 1248 55008 1248 0 output_no[141]
rlabel metal2 55392 492 55392 492 0 output_no[142]
rlabel metal2 55776 702 55776 702 0 output_no[143]
rlabel metal2 56160 660 56160 660 0 output_no[144]
rlabel metal2 56544 1290 56544 1290 0 output_no[145]
rlabel metal2 56928 492 56928 492 0 output_no[146]
rlabel metal2 57312 492 57312 492 0 output_no[147]
rlabel metal2 57696 870 57696 870 0 output_no[148]
rlabel metal2 58080 492 58080 492 0 output_no[149]
rlabel metal2 6720 1890 6720 1890 0 output_no[14]
rlabel metal2 58464 1038 58464 1038 0 output_no[150]
rlabel metal2 58848 1248 58848 1248 0 output_no[151]
rlabel metal2 59232 2004 59232 2004 0 output_no[152]
rlabel metal2 59616 282 59616 282 0 output_no[153]
rlabel metal2 60000 492 60000 492 0 output_no[154]
rlabel metal2 60384 492 60384 492 0 output_no[155]
rlabel metal2 60720 4704 60720 4704 0 output_no[156]
rlabel metal2 61200 2436 61200 2436 0 output_no[157]
rlabel metal2 61584 2436 61584 2436 0 output_no[158]
rlabel metal2 61920 954 61920 954 0 output_no[159]
rlabel metal2 6624 114 6624 114 0 output_no[15]
rlabel metal2 62304 870 62304 870 0 output_no[160]
rlabel metal2 62784 1344 62784 1344 0 output_no[161]
rlabel metal2 63072 408 63072 408 0 output_no[162]
rlabel metal2 63408 1260 63408 1260 0 output_no[163]
rlabel metal2 63840 492 63840 492 0 output_no[164]
rlabel metal2 64320 2394 64320 2394 0 output_no[165]
rlabel metal2 64608 282 64608 282 0 output_no[166]
rlabel metal2 64992 324 64992 324 0 output_no[167]
rlabel metal2 65376 492 65376 492 0 output_no[168]
rlabel metal2 65712 3192 65712 3192 0 output_no[169]
rlabel metal2 7008 534 7008 534 0 output_no[16]
rlabel metal2 66096 3192 66096 3192 0 output_no[170]
rlabel metal2 66528 450 66528 450 0 output_no[171]
rlabel metal2 66912 2856 66912 2856 0 output_no[172]
rlabel metal2 67248 3192 67248 3192 0 output_no[173]
rlabel metal2 67488 1974 67488 1974 0 output_no[174]
rlabel metal2 68064 450 68064 450 0 output_no[175]
rlabel metal2 68544 3192 68544 3192 0 output_no[176]
rlabel metal2 68832 492 68832 492 0 output_no[177]
rlabel metal2 69504 2856 69504 2856 0 output_no[178]
rlabel metal2 69744 3192 69744 3192 0 output_no[179]
rlabel metal2 7440 3192 7440 3192 0 output_no[17]
rlabel metal2 70176 3192 70176 3192 0 output_no[180]
rlabel metal2 70368 450 70368 450 0 output_no[181]
rlabel metal2 71040 2856 71040 2856 0 output_no[182]
rlabel metal2 71328 3192 71328 3192 0 output_no[183]
rlabel metal2 71520 450 71520 450 0 output_no[184]
rlabel metal2 71904 408 71904 408 0 output_no[185]
rlabel metal2 72576 2856 72576 2856 0 output_no[186]
rlabel metal2 72864 3192 72864 3192 0 output_no[187]
rlabel metal2 73056 492 73056 492 0 output_no[188]
rlabel metal2 73392 1428 73392 1428 0 output_no[189]
rlabel metal2 7824 3192 7824 3192 0 output_no[18]
rlabel metal2 73776 1428 73776 1428 0 output_no[190]
rlabel metal2 74160 1428 74160 1428 0 output_no[191]
rlabel metal2 74688 1512 74688 1512 0 output_no[192]
rlabel metal2 74976 492 74976 492 0 output_no[193]
rlabel metal2 75360 492 75360 492 0 output_no[194]
rlabel metal2 75696 1344 75696 1344 0 output_no[195]
rlabel metal2 76128 492 76128 492 0 output_no[196]
rlabel metal2 76512 450 76512 450 0 output_no[197]
rlabel metal2 76896 450 76896 450 0 output_no[198]
rlabel metal2 77280 282 77280 282 0 output_no[199]
rlabel metal2 8160 1932 8160 1932 0 output_no[19]
rlabel metal2 1728 2310 1728 2310 0 output_no[1]
rlabel metal2 77664 492 77664 492 0 output_no[200]
rlabel metal2 78048 492 78048 492 0 output_no[201]
rlabel metal2 78432 492 78432 492 0 output_no[202]
rlabel metal2 78672 1680 78672 1680 0 output_no[203]
rlabel metal2 79200 282 79200 282 0 output_no[204]
rlabel metal2 79584 492 79584 492 0 output_no[205]
rlabel metal2 79968 324 79968 324 0 output_no[206]
rlabel metal2 80352 198 80352 198 0 output_no[207]
rlabel metal2 80736 870 80736 870 0 output_no[208]
rlabel metal2 81120 492 81120 492 0 output_no[209]
rlabel metal2 8592 3192 8592 3192 0 output_no[20]
rlabel metal2 81504 492 81504 492 0 output_no[210]
rlabel metal2 81984 1134 81984 1134 0 output_no[211]
rlabel metal2 82320 3192 82320 3192 0 output_no[212]
rlabel metal2 82704 3192 82704 3192 0 output_no[213]
rlabel metal2 83088 3192 83088 3192 0 output_no[214]
rlabel metal2 83328 1932 83328 1932 0 output_no[215]
rlabel metal2 83808 408 83808 408 0 output_no[216]
rlabel metal2 84096 2856 84096 2856 0 output_no[217]
rlabel metal2 84576 3192 84576 3192 0 output_no[218]
rlabel metal2 84864 1932 84864 1932 0 output_no[219]
rlabel metal2 8976 3192 8976 3192 0 output_no[21]
rlabel metal2 85344 450 85344 450 0 output_no[220]
rlabel metal2 85728 408 85728 408 0 output_no[221]
rlabel metal2 86016 1722 86016 1722 0 output_no[222]
rlabel metal2 86400 2394 86400 2394 0 output_no[223]
rlabel metal2 86928 3192 86928 3192 0 output_no[224]
rlabel metal2 87264 492 87264 492 0 output_no[225]
rlabel metal2 87648 492 87648 492 0 output_no[226]
rlabel metal2 88032 492 88032 492 0 output_no[227]
rlabel metal2 88416 492 88416 492 0 output_no[228]
rlabel metal2 88800 492 88800 492 0 output_no[229]
rlabel metal2 9360 3192 9360 3192 0 output_no[22]
rlabel metal2 89184 408 89184 408 0 output_no[230]
rlabel metal2 89568 492 89568 492 0 output_no[231]
rlabel metal2 89952 492 89952 492 0 output_no[232]
rlabel metal2 90336 492 90336 492 0 output_no[233]
rlabel metal2 90720 240 90720 240 0 output_no[234]
rlabel metal2 91104 492 91104 492 0 output_no[235]
rlabel metal2 91488 450 91488 450 0 output_no[236]
rlabel metal2 91872 492 91872 492 0 output_no[237]
rlabel metal2 92256 366 92256 366 0 output_no[238]
rlabel metal2 92640 492 92640 492 0 output_no[239]
rlabel metal2 9744 3192 9744 3192 0 output_no[23]
rlabel metal2 93024 450 93024 450 0 output_no[240]
rlabel metal2 93024 2478 93024 2478 0 output_no[241]
rlabel metal2 93360 3192 93360 3192 0 output_no[242]
rlabel metal2 93696 1890 93696 1890 0 output_no[243]
rlabel metal2 94224 3192 94224 3192 0 output_no[244]
rlabel metal2 94608 3192 94608 3192 0 output_no[245]
rlabel metal2 95328 324 95328 324 0 output_no[246]
rlabel metal2 95232 2478 95232 2478 0 output_no[247]
rlabel metal2 96096 492 96096 492 0 output_no[248]
rlabel metal2 96144 3192 96144 3192 0 output_no[249]
rlabel metal2 10080 2856 10080 2856 0 output_no[24]
rlabel metal2 96480 1974 96480 1974 0 output_no[250]
rlabel metal2 96864 2016 96864 2016 0 output_no[251]
rlabel metal2 97248 1932 97248 1932 0 output_no[252]
rlabel metal2 98016 492 98016 492 0 output_no[253]
rlabel metal2 98016 2184 98016 2184 0 output_no[254]
rlabel metal2 98784 450 98784 450 0 output_no[255]
rlabel metal2 10512 3192 10512 3192 0 output_no[25]
rlabel metal2 10896 3192 10896 3192 0 output_no[26]
rlabel metal2 11280 3192 11280 3192 0 output_no[27]
rlabel metal2 11616 534 11616 534 0 output_no[28]
rlabel metal2 12000 492 12000 492 0 output_no[29]
rlabel metal2 1968 3192 1968 3192 0 output_no[2]
rlabel metal2 12384 492 12384 492 0 output_no[30]
rlabel metal2 12768 1344 12768 1344 0 output_no[31]
rlabel metal2 13152 492 13152 492 0 output_no[32]
rlabel metal2 13536 492 13536 492 0 output_no[33]
rlabel metal2 13920 492 13920 492 0 output_no[34]
rlabel metal2 14304 408 14304 408 0 output_no[35]
rlabel metal2 14688 492 14688 492 0 output_no[36]
rlabel metal2 15072 492 15072 492 0 output_no[37]
rlabel metal2 15456 450 15456 450 0 output_no[38]
rlabel metal2 15840 492 15840 492 0 output_no[39]
rlabel metal2 2016 450 2016 450 0 output_no[3]
rlabel metal2 16224 492 16224 492 0 output_no[40]
rlabel metal2 16608 492 16608 492 0 output_no[41]
rlabel metal2 16992 492 16992 492 0 output_no[42]
rlabel metal2 17376 492 17376 492 0 output_no[43]
rlabel metal2 17760 408 17760 408 0 output_no[44]
rlabel metal2 18144 492 18144 492 0 output_no[45]
rlabel metal2 18528 450 18528 450 0 output_no[46]
rlabel metal2 18912 450 18912 450 0 output_no[47]
rlabel metal2 19296 72 19296 72 0 output_no[48]
rlabel metal2 19680 114 19680 114 0 output_no[49]
rlabel metal2 2400 282 2400 282 0 output_no[4]
rlabel via2 20064 72 20064 72 0 output_no[50]
rlabel metal2 20448 408 20448 408 0 output_no[51]
rlabel metal2 20832 492 20832 492 0 output_no[52]
rlabel metal2 21216 492 21216 492 0 output_no[53]
rlabel metal2 21600 492 21600 492 0 output_no[54]
rlabel metal2 22032 1344 22032 1344 0 output_no[55]
rlabel metal2 22368 408 22368 408 0 output_no[56]
rlabel metal2 22752 408 22752 408 0 output_no[57]
rlabel metal2 23136 408 23136 408 0 output_no[58]
rlabel metal2 23568 1344 23568 1344 0 output_no[59]
rlabel metal2 3072 2100 3072 2100 0 output_no[5]
rlabel metal2 23904 282 23904 282 0 output_no[60]
rlabel metal2 24288 408 24288 408 0 output_no[61]
rlabel metal2 24672 450 24672 450 0 output_no[62]
rlabel metal2 25056 450 25056 450 0 output_no[63]
rlabel metal2 25440 1626 25440 1626 0 output_no[64]
rlabel metal2 25824 1626 25824 1626 0 output_no[65]
rlabel metal2 26208 1626 26208 1626 0 output_no[66]
rlabel metal2 26544 2100 26544 2100 0 output_no[67]
rlabel metal2 26976 1290 26976 1290 0 output_no[68]
rlabel metal2 27360 1290 27360 1290 0 output_no[69]
rlabel metal2 3456 2100 3456 2100 0 output_no[6]
rlabel metal2 27744 1290 27744 1290 0 output_no[70]
rlabel metal2 28080 2100 28080 2100 0 output_no[71]
rlabel metal2 28512 1626 28512 1626 0 output_no[72]
rlabel metal2 28896 1626 28896 1626 0 output_no[73]
rlabel metal2 29280 1626 29280 1626 0 output_no[74]
rlabel metal2 29664 1290 29664 1290 0 output_no[75]
rlabel metal2 29904 3192 29904 3192 0 output_no[76]
rlabel metal2 30192 3192 30192 3192 0 output_no[77]
rlabel metal2 30576 3192 30576 3192 0 output_no[78]
rlabel metal2 30816 1932 30816 1932 0 output_no[79]
rlabel metal2 3840 2226 3840 2226 0 output_no[7]
rlabel metal2 31776 2142 31776 2142 0 output_no[80]
rlabel metal2 31344 3192 31344 3192 0 output_no[81]
rlabel metal2 32352 198 32352 198 0 output_no[82]
rlabel metal2 32304 3192 32304 3192 0 output_no[83]
rlabel metal2 33120 324 33120 324 0 output_no[84]
rlabel metal2 33504 366 33504 366 0 output_no[85]
rlabel metal2 33264 3192 33264 3192 0 output_no[86]
rlabel metal2 33792 3612 33792 3612 0 output_no[87]
rlabel metal2 34176 3192 34176 3192 0 output_no[88]
rlabel metal2 35040 240 35040 240 0 output_no[89]
rlabel metal2 4272 3192 4272 3192 0 output_no[8]
rlabel metal2 34848 2814 34848 2814 0 output_no[90]
rlabel metal2 35472 2856 35472 2856 0 output_no[91]
rlabel metal2 35760 3192 35760 3192 0 output_no[92]
rlabel metal2 36576 198 36576 198 0 output_no[93]
rlabel metal2 36960 156 36960 156 0 output_no[94]
rlabel metal2 37008 3192 37008 3192 0 output_no[95]
rlabel metal2 37728 1890 37728 1890 0 output_no[96]
rlabel metal2 38112 492 38112 492 0 output_no[97]
rlabel metal2 38352 1260 38352 1260 0 output_no[98]
rlabel metal2 38736 1344 38736 1344 0 output_no[99]
rlabel metal2 4320 324 4320 324 0 output_no[9]
rlabel metal2 1056 492 1056 492 0 output_o[0]
rlabel metal2 39456 492 39456 492 0 output_o[100]
rlabel metal2 39840 240 39840 240 0 output_o[101]
rlabel metal2 40224 492 40224 492 0 output_o[102]
rlabel metal2 40608 282 40608 282 0 output_o[103]
rlabel metal2 40992 492 40992 492 0 output_o[104]
rlabel metal2 41376 282 41376 282 0 output_o[105]
rlabel metal2 41760 492 41760 492 0 output_o[106]
rlabel metal2 42144 240 42144 240 0 output_o[107]
rlabel metal2 42528 492 42528 492 0 output_o[108]
rlabel metal2 42912 240 42912 240 0 output_o[109]
rlabel metal2 4896 492 4896 492 0 output_o[10]
rlabel metal2 43296 492 43296 492 0 output_o[110]
rlabel metal2 43680 198 43680 198 0 output_o[111]
rlabel metal2 44064 282 44064 282 0 output_o[112]
rlabel metal2 44448 366 44448 366 0 output_o[113]
rlabel metal2 44832 156 44832 156 0 output_o[114]
rlabel metal2 45216 366 45216 366 0 output_o[115]
rlabel metal2 45600 240 45600 240 0 output_o[116]
rlabel metal2 45984 366 45984 366 0 output_o[117]
rlabel metal2 46368 282 46368 282 0 output_o[118]
rlabel metal2 46752 366 46752 366 0 output_o[119]
rlabel metal2 5280 492 5280 492 0 output_o[11]
rlabel metal2 47136 282 47136 282 0 output_o[120]
rlabel metal2 47520 366 47520 366 0 output_o[121]
rlabel metal2 47904 282 47904 282 0 output_o[122]
rlabel metal2 48288 366 48288 366 0 output_o[123]
rlabel metal2 48672 282 48672 282 0 output_o[124]
rlabel metal2 49056 366 49056 366 0 output_o[125]
rlabel metal2 49440 114 49440 114 0 output_o[126]
rlabel metal2 49824 282 49824 282 0 output_o[127]
rlabel metal2 50208 240 50208 240 0 output_o[128]
rlabel metal2 50592 450 50592 450 0 output_o[129]
rlabel metal2 5664 492 5664 492 0 output_o[12]
rlabel metal2 50976 492 50976 492 0 output_o[130]
rlabel metal2 51360 576 51360 576 0 output_o[131]
rlabel metal2 51744 534 51744 534 0 output_o[132]
rlabel metal2 52128 492 52128 492 0 output_o[133]
rlabel metal2 52512 408 52512 408 0 output_o[134]
rlabel metal2 52896 660 52896 660 0 output_o[135]
rlabel metal2 53280 744 53280 744 0 output_o[136]
rlabel metal2 53664 492 53664 492 0 output_o[137]
rlabel metal2 54048 870 54048 870 0 output_o[138]
rlabel metal2 54432 198 54432 198 0 output_o[139]
rlabel metal2 6048 492 6048 492 0 output_o[13]
rlabel metal3 55008 4116 55008 4116 0 output_o[140]
rlabel metal2 55200 1416 55200 1416 0 output_o[141]
rlabel metal2 55584 408 55584 408 0 output_o[142]
rlabel metal2 55968 576 55968 576 0 output_o[143]
rlabel metal2 56352 282 56352 282 0 output_o[144]
rlabel metal2 56736 408 56736 408 0 output_o[145]
rlabel metal2 57120 408 57120 408 0 output_o[146]
rlabel metal2 57504 576 57504 576 0 output_o[147]
rlabel metal2 57888 870 57888 870 0 output_o[148]
rlabel metal2 58272 492 58272 492 0 output_o[149]
rlabel metal2 6432 492 6432 492 0 output_o[14]
rlabel metal2 58656 1206 58656 1206 0 output_o[150]
rlabel metal2 59040 870 59040 870 0 output_o[151]
rlabel metal2 59424 2004 59424 2004 0 output_o[152]
rlabel metal2 59808 282 59808 282 0 output_o[153]
rlabel metal2 60192 450 60192 450 0 output_o[154]
rlabel metal2 60576 492 60576 492 0 output_o[155]
rlabel metal2 60960 492 60960 492 0 output_o[156]
rlabel metal2 61344 1248 61344 1248 0 output_o[157]
rlabel metal2 61728 1248 61728 1248 0 output_o[158]
rlabel metal2 62112 2004 62112 2004 0 output_o[159]
rlabel metal2 6816 198 6816 198 0 output_o[15]
rlabel metal2 62496 492 62496 492 0 output_o[160]
rlabel metal2 62880 282 62880 282 0 output_o[161]
rlabel metal2 63264 492 63264 492 0 output_o[162]
rlabel metal2 63648 282 63648 282 0 output_o[163]
rlabel metal2 64032 282 64032 282 0 output_o[164]
rlabel metal2 64416 408 64416 408 0 output_o[165]
rlabel metal2 64800 282 64800 282 0 output_o[166]
rlabel metal2 65184 240 65184 240 0 output_o[167]
rlabel metal2 65568 492 65568 492 0 output_o[168]
rlabel metal2 65952 282 65952 282 0 output_o[169]
rlabel metal2 7200 282 7200 282 0 output_o[16]
rlabel metal2 66336 240 66336 240 0 output_o[170]
rlabel metal2 66720 492 66720 492 0 output_o[171]
rlabel metal2 67104 492 67104 492 0 output_o[172]
rlabel metal2 67488 366 67488 366 0 output_o[173]
rlabel metal2 67872 282 67872 282 0 output_o[174]
rlabel metal2 68256 492 68256 492 0 output_o[175]
rlabel metal2 68640 366 68640 366 0 output_o[176]
rlabel metal2 69024 282 69024 282 0 output_o[177]
rlabel metal2 69408 492 69408 492 0 output_o[178]
rlabel metal2 69792 282 69792 282 0 output_o[179]
rlabel metal2 7584 492 7584 492 0 output_o[17]
rlabel metal2 70176 492 70176 492 0 output_o[180]
rlabel metal2 70560 114 70560 114 0 output_o[181]
rlabel metal2 70944 282 70944 282 0 output_o[182]
rlabel metal2 71328 282 71328 282 0 output_o[183]
rlabel metal2 71712 492 71712 492 0 output_o[184]
rlabel metal2 72096 492 72096 492 0 output_o[185]
rlabel metal2 72480 282 72480 282 0 output_o[186]
rlabel metal2 72864 492 72864 492 0 output_o[187]
rlabel metal2 73248 156 73248 156 0 output_o[188]
rlabel metal2 73632 492 73632 492 0 output_o[189]
rlabel metal2 7968 282 7968 282 0 output_o[18]
rlabel metal2 74016 156 74016 156 0 output_o[190]
rlabel metal2 74400 282 74400 282 0 output_o[191]
rlabel metal2 74784 492 74784 492 0 output_o[192]
rlabel metal2 75168 282 75168 282 0 output_o[193]
rlabel metal2 75552 492 75552 492 0 output_o[194]
rlabel metal2 75936 282 75936 282 0 output_o[195]
rlabel metal2 76320 492 76320 492 0 output_o[196]
rlabel metal2 76704 282 76704 282 0 output_o[197]
rlabel metal2 77088 492 77088 492 0 output_o[198]
rlabel metal2 77472 282 77472 282 0 output_o[199]
rlabel metal2 8352 492 8352 492 0 output_o[19]
rlabel metal2 1440 492 1440 492 0 output_o[1]
rlabel metal2 77856 240 77856 240 0 output_o[200]
rlabel metal2 78240 240 78240 240 0 output_o[201]
rlabel metal2 78624 282 78624 282 0 output_o[202]
rlabel metal2 79008 492 79008 492 0 output_o[203]
rlabel metal2 79392 198 79392 198 0 output_o[204]
rlabel metal2 79776 492 79776 492 0 output_o[205]
rlabel metal2 80160 282 80160 282 0 output_o[206]
rlabel metal2 80544 492 80544 492 0 output_o[207]
rlabel metal2 80928 492 80928 492 0 output_o[208]
rlabel metal2 81312 492 81312 492 0 output_o[209]
rlabel metal2 8736 282 8736 282 0 output_o[20]
rlabel metal2 81696 282 81696 282 0 output_o[210]
rlabel metal2 82080 492 82080 492 0 output_o[211]
rlabel metal2 82464 492 82464 492 0 output_o[212]
rlabel metal2 82848 408 82848 408 0 output_o[213]
rlabel metal2 83232 492 83232 492 0 output_o[214]
rlabel metal2 83616 492 83616 492 0 output_o[215]
rlabel metal2 84000 492 84000 492 0 output_o[216]
rlabel metal2 84384 492 84384 492 0 output_o[217]
rlabel metal2 84768 492 84768 492 0 output_o[218]
rlabel metal2 85152 492 85152 492 0 output_o[219]
rlabel metal2 9120 492 9120 492 0 output_o[21]
rlabel metal2 85536 492 85536 492 0 output_o[220]
rlabel metal2 85920 492 85920 492 0 output_o[221]
rlabel metal2 86304 492 86304 492 0 output_o[222]
rlabel metal2 86688 492 86688 492 0 output_o[223]
rlabel metal2 87072 492 87072 492 0 output_o[224]
rlabel metal2 87456 492 87456 492 0 output_o[225]
rlabel metal2 87840 492 87840 492 0 output_o[226]
rlabel metal2 88224 492 88224 492 0 output_o[227]
rlabel metal2 88608 492 88608 492 0 output_o[228]
rlabel metal2 88992 492 88992 492 0 output_o[229]
rlabel metal2 9504 282 9504 282 0 output_o[22]
rlabel metal2 89376 492 89376 492 0 output_o[230]
rlabel metal2 89760 492 89760 492 0 output_o[231]
rlabel metal2 90144 492 90144 492 0 output_o[232]
rlabel metal2 90528 492 90528 492 0 output_o[233]
rlabel metal2 90912 492 90912 492 0 output_o[234]
rlabel metal2 91296 492 91296 492 0 output_o[235]
rlabel metal2 91680 282 91680 282 0 output_o[236]
rlabel metal2 92064 492 92064 492 0 output_o[237]
rlabel metal2 92448 492 92448 492 0 output_o[238]
rlabel metal2 92832 492 92832 492 0 output_o[239]
rlabel metal2 9888 492 9888 492 0 output_o[23]
rlabel metal2 93216 492 93216 492 0 output_o[240]
rlabel metal2 93600 492 93600 492 0 output_o[241]
rlabel metal2 93984 492 93984 492 0 output_o[242]
rlabel metal2 94368 492 94368 492 0 output_o[243]
rlabel metal2 94752 492 94752 492 0 output_o[244]
rlabel via2 95136 72 95136 72 0 output_o[245]
rlabel metal2 95520 492 95520 492 0 output_o[246]
rlabel metal2 95904 492 95904 492 0 output_o[247]
rlabel metal2 96288 492 96288 492 0 output_o[248]
rlabel metal2 96672 492 96672 492 0 output_o[249]
rlabel metal2 10272 282 10272 282 0 output_o[24]
rlabel metal2 97056 492 97056 492 0 output_o[250]
rlabel metal2 97440 282 97440 282 0 output_o[251]
rlabel metal2 97824 408 97824 408 0 output_o[252]
rlabel metal2 98208 450 98208 450 0 output_o[253]
rlabel metal2 98592 492 98592 492 0 output_o[254]
rlabel metal2 98976 492 98976 492 0 output_o[255]
rlabel metal2 10656 492 10656 492 0 output_o[25]
rlabel metal2 11040 156 11040 156 0 output_o[26]
rlabel metal2 11424 492 11424 492 0 output_o[27]
rlabel metal2 11808 114 11808 114 0 output_o[28]
rlabel metal2 12192 282 12192 282 0 output_o[29]
rlabel metal2 1824 492 1824 492 0 output_o[2]
rlabel metal2 12576 492 12576 492 0 output_o[30]
rlabel metal2 12960 282 12960 282 0 output_o[31]
rlabel metal2 13344 492 13344 492 0 output_o[32]
rlabel metal2 13728 282 13728 282 0 output_o[33]
rlabel metal2 14112 492 14112 492 0 output_o[34]
rlabel metal2 14496 366 14496 366 0 output_o[35]
rlabel metal2 14880 492 14880 492 0 output_o[36]
rlabel metal2 15264 156 15264 156 0 output_o[37]
rlabel metal2 15648 156 15648 156 0 output_o[38]
rlabel metal2 16032 492 16032 492 0 output_o[39]
rlabel metal2 2208 492 2208 492 0 output_o[3]
rlabel metal2 16416 156 16416 156 0 output_o[40]
rlabel metal2 16800 534 16800 534 0 output_o[41]
rlabel metal2 17184 492 17184 492 0 output_o[42]
rlabel metal2 17568 282 17568 282 0 output_o[43]
rlabel metal2 17952 450 17952 450 0 output_o[44]
rlabel metal2 18336 492 18336 492 0 output_o[45]
rlabel metal2 18720 282 18720 282 0 output_o[46]
rlabel metal2 19104 492 19104 492 0 output_o[47]
rlabel metal2 19488 198 19488 198 0 output_o[48]
rlabel via2 19872 72 19872 72 0 output_o[49]
rlabel metal2 2592 492 2592 492 0 output_o[4]
rlabel metal2 20256 492 20256 492 0 output_o[50]
rlabel metal2 20640 282 20640 282 0 output_o[51]
rlabel metal2 21024 492 21024 492 0 output_o[52]
rlabel metal2 21408 282 21408 282 0 output_o[53]
rlabel metal2 21792 198 21792 198 0 output_o[54]
rlabel metal2 22176 156 22176 156 0 output_o[55]
rlabel metal2 22560 492 22560 492 0 output_o[56]
rlabel metal2 22944 282 22944 282 0 output_o[57]
rlabel metal2 23328 492 23328 492 0 output_o[58]
rlabel metal2 23712 156 23712 156 0 output_o[59]
rlabel metal2 2976 492 2976 492 0 output_o[5]
rlabel metal2 24096 492 24096 492 0 output_o[60]
rlabel metal2 24480 492 24480 492 0 output_o[61]
rlabel metal2 24864 282 24864 282 0 output_o[62]
rlabel metal2 25248 492 25248 492 0 output_o[63]
rlabel metal2 25632 198 25632 198 0 output_o[64]
rlabel metal2 26016 282 26016 282 0 output_o[65]
rlabel metal2 26400 366 26400 366 0 output_o[66]
rlabel metal2 26784 282 26784 282 0 output_o[67]
rlabel metal2 27168 366 27168 366 0 output_o[68]
rlabel metal2 27552 282 27552 282 0 output_o[69]
rlabel metal2 3360 492 3360 492 0 output_o[6]
rlabel metal2 27936 366 27936 366 0 output_o[70]
rlabel metal2 28320 282 28320 282 0 output_o[71]
rlabel metal2 28704 366 28704 366 0 output_o[72]
rlabel metal2 29088 198 29088 198 0 output_o[73]
rlabel metal2 29472 282 29472 282 0 output_o[74]
rlabel metal2 29856 366 29856 366 0 output_o[75]
rlabel metal2 30240 282 30240 282 0 output_o[76]
rlabel metal2 30624 366 30624 366 0 output_o[77]
rlabel metal2 31008 324 31008 324 0 output_o[78]
rlabel metal2 31392 492 31392 492 0 output_o[79]
rlabel metal2 3744 492 3744 492 0 output_o[7]
rlabel metal2 31776 870 31776 870 0 output_o[80]
rlabel metal2 32160 660 32160 660 0 output_o[81]
rlabel metal2 32544 240 32544 240 0 output_o[82]
rlabel metal2 32928 282 32928 282 0 output_o[83]
rlabel metal2 33312 492 33312 492 0 output_o[84]
rlabel metal2 33696 282 33696 282 0 output_o[85]
rlabel metal2 34080 240 34080 240 0 output_o[86]
rlabel metal2 34464 282 34464 282 0 output_o[87]
rlabel metal2 34848 240 34848 240 0 output_o[88]
rlabel metal2 35232 492 35232 492 0 output_o[89]
rlabel metal2 4128 492 4128 492 0 output_o[8]
rlabel metal2 35616 114 35616 114 0 output_o[90]
rlabel metal2 36000 492 36000 492 0 output_o[91]
rlabel metal2 36384 282 36384 282 0 output_o[92]
rlabel metal2 36768 282 36768 282 0 output_o[93]
rlabel metal2 37152 282 37152 282 0 output_o[94]
rlabel metal2 37536 240 37536 240 0 output_o[95]
rlabel metal2 37920 492 37920 492 0 output_o[96]
rlabel metal2 38304 282 38304 282 0 output_o[97]
rlabel metal2 38688 492 38688 492 0 output_o[98]
rlabel metal2 39072 282 39072 282 0 output_o[99]
rlabel metal2 4512 282 4512 282 0 output_o[9]
<< properties >>
string FIXED_BBOX 0 0 100000 10000
<< end >>
