module decoder (ena_i,
    input_ni,
    output_no,
    output_o);
 input ena_i;
 input [7:0] input_ni;
 output [255:0] output_no;
 output [255:0] output_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;

 sg13g2_inv_1 _095_ (.Y(_004_),
    .A(input_ni[6]));
 sg13g2_nor2_1 _096_ (.A(input_ni[3]),
    .B(input_ni[2]),
    .Y(_005_));
 sg13g2_nor2_1 _097_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .Y(_006_));
 sg13g2_nor4_1 _098_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .C(input_ni[3]),
    .D(input_ni[2]),
    .Y(_007_));
 sg13g2_nor2b_1 _099_ (.A(input_ni[7]),
    .B_N(input_ni[6]),
    .Y(_008_));
 sg13g2_and4_1 _100_ (.A(input_ni[4]),
    .B(input_ni[5]),
    .C(ena_i),
    .D(_008_),
    .X(_009_));
 sg13g2_nand4_1 _101_ (.B(input_ni[5]),
    .C(ena_i),
    .A(input_ni[4]),
    .Y(_010_),
    .D(_008_));
 sg13g2_and2_1 _102_ (.A(_007_),
    .B(_009_),
    .X(output_o[143]));
 sg13g2_nand2_1 _103_ (.Y(output_no[143]),
    .A(_007_),
    .B(_009_));
 sg13g2_and2_1 _104_ (.A(input_ni[3]),
    .B(input_ni[2]),
    .X(_011_));
 sg13g2_and2_1 _105_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .X(_012_));
 sg13g2_nand2_1 _106_ (.Y(_013_),
    .A(_011_),
    .B(_012_));
 sg13g2_nor2b_1 _107_ (.A(input_ni[4]),
    .B_N(input_ni[5]),
    .Y(_014_));
 sg13g2_and3_1 _108_ (.X(_015_),
    .A(ena_i),
    .B(_008_),
    .C(_014_));
 sg13g2_nand3_1 _109_ (.B(_008_),
    .C(_014_),
    .A(ena_i),
    .Y(_016_));
 sg13g2_nor2_1 _110_ (.A(_013_),
    .B(_016_),
    .Y(output_o[144]));
 sg13g2_nand2b_1 _111_ (.Y(output_no[144]),
    .B(_015_),
    .A_N(_013_));
 sg13g2_nor2b_1 _112_ (.A(input_ni[0]),
    .B_N(input_ni[1]),
    .Y(_017_));
 sg13g2_nand2_1 _113_ (.Y(_018_),
    .A(_011_),
    .B(_017_));
 sg13g2_nor2_1 _114_ (.A(_016_),
    .B(_018_),
    .Y(output_o[145]));
 sg13g2_or2_1 _115_ (.X(output_no[145]),
    .B(_018_),
    .A(_016_));
 sg13g2_nor2b_1 _116_ (.A(input_ni[1]),
    .B_N(input_ni[0]),
    .Y(_019_));
 sg13g2_nand2_1 _117_ (.Y(_020_),
    .A(_011_),
    .B(_019_));
 sg13g2_nor2_1 _118_ (.A(_016_),
    .B(_020_),
    .Y(output_o[146]));
 sg13g2_or2_1 _119_ (.X(output_no[146]),
    .B(_020_),
    .A(_016_));
 sg13g2_nand2_1 _120_ (.Y(_021_),
    .A(_006_),
    .B(_011_));
 sg13g2_nor2_1 _121_ (.A(_016_),
    .B(_021_),
    .Y(output_o[147]));
 sg13g2_or2_1 _122_ (.X(output_no[147]),
    .B(_021_),
    .A(_016_));
 sg13g2_nor2b_1 _123_ (.A(input_ni[2]),
    .B_N(input_ni[3]),
    .Y(_022_));
 sg13g2_nand2_1 _124_ (.Y(_023_),
    .A(_012_),
    .B(_022_));
 sg13g2_nor2_1 _125_ (.A(_016_),
    .B(_023_),
    .Y(output_o[148]));
 sg13g2_or2_1 _126_ (.X(output_no[148]),
    .B(_023_),
    .A(_016_));
 sg13g2_nand2_1 _127_ (.Y(_024_),
    .A(_017_),
    .B(_022_));
 sg13g2_nor2_1 _128_ (.A(_016_),
    .B(_024_),
    .Y(output_o[149]));
 sg13g2_or2_1 _129_ (.X(output_no[149]),
    .B(_024_),
    .A(_016_));
 sg13g2_nand2_1 _130_ (.Y(_025_),
    .A(_019_),
    .B(_022_));
 sg13g2_nor2_1 _131_ (.A(_016_),
    .B(_025_),
    .Y(output_o[150]));
 sg13g2_or2_1 _132_ (.X(output_no[150]),
    .B(_025_),
    .A(_016_));
 sg13g2_nand2_1 _133_ (.Y(_026_),
    .A(_006_),
    .B(_022_));
 sg13g2_nor2_1 _134_ (.A(_016_),
    .B(_026_),
    .Y(output_o[151]));
 sg13g2_or2_1 _135_ (.X(output_no[151]),
    .B(_026_),
    .A(_016_));
 sg13g2_nor2b_1 _136_ (.A(input_ni[3]),
    .B_N(input_ni[2]),
    .Y(_027_));
 sg13g2_nand2_1 _137_ (.Y(_028_),
    .A(_012_),
    .B(_027_));
 sg13g2_nor2_1 _138_ (.A(_016_),
    .B(_028_),
    .Y(output_o[152]));
 sg13g2_or2_1 _139_ (.X(output_no[152]),
    .B(_028_),
    .A(_016_));
 sg13g2_nand2_1 _140_ (.Y(_029_),
    .A(_017_),
    .B(_027_));
 sg13g2_nor2_1 _141_ (.A(_016_),
    .B(_029_),
    .Y(output_o[153]));
 sg13g2_or2_1 _142_ (.X(output_no[153]),
    .B(_029_),
    .A(_016_));
 sg13g2_nand2_1 _143_ (.Y(_030_),
    .A(_019_),
    .B(_027_));
 sg13g2_nor2_1 _144_ (.A(_016_),
    .B(_030_),
    .Y(output_o[154]));
 sg13g2_or2_1 _145_ (.X(output_no[154]),
    .B(_030_),
    .A(_016_));
 sg13g2_nand2_1 _146_ (.Y(_031_),
    .A(_006_),
    .B(_027_));
 sg13g2_nor2_1 _147_ (.A(_016_),
    .B(_031_),
    .Y(output_o[155]));
 sg13g2_or2_1 _148_ (.X(output_no[155]),
    .B(_031_),
    .A(_016_));
 sg13g2_nand2_1 _149_ (.Y(_032_),
    .A(_005_),
    .B(_012_));
 sg13g2_nor2_1 _150_ (.A(_016_),
    .B(_032_),
    .Y(output_o[156]));
 sg13g2_or2_1 _151_ (.X(output_no[156]),
    .B(_032_),
    .A(_016_));
 sg13g2_nand2_1 _152_ (.Y(_033_),
    .A(_005_),
    .B(_017_));
 sg13g2_nor2_1 _153_ (.A(_016_),
    .B(_033_),
    .Y(output_o[157]));
 sg13g2_or2_1 _154_ (.X(output_no[157]),
    .B(_033_),
    .A(_016_));
 sg13g2_nand2_1 _155_ (.Y(_034_),
    .A(_005_),
    .B(_019_));
 sg13g2_nor2_1 _156_ (.A(_016_),
    .B(_034_),
    .Y(output_o[158]));
 sg13g2_or2_1 _157_ (.X(output_no[158]),
    .B(_034_),
    .A(_016_));
 sg13g2_and2_1 _158_ (.A(_007_),
    .B(_015_),
    .X(output_o[159]));
 sg13g2_nand2_1 _159_ (.Y(output_no[159]),
    .A(_007_),
    .B(_015_));
 sg13g2_nor2b_1 _160_ (.A(input_ni[5]),
    .B_N(input_ni[4]),
    .Y(_035_));
 sg13g2_and2_1 _161_ (.A(_008_),
    .B(_035_),
    .X(_036_));
 sg13g2_nand2_1 _162_ (.Y(_037_),
    .A(_008_),
    .B(_035_));
 sg13g2_and3_1 _163_ (.X(_038_),
    .A(ena_i),
    .B(_011_),
    .C(_012_));
 sg13g2_nand3_1 _164_ (.B(_011_),
    .C(_012_),
    .A(ena_i),
    .Y(_039_));
 sg13g2_nor2_1 _165_ (.A(_037_),
    .B(_039_),
    .Y(output_o[160]));
 sg13g2_nand2_1 _166_ (.Y(output_no[160]),
    .A(_036_),
    .B(_038_));
 sg13g2_and3_1 _167_ (.X(_040_),
    .A(ena_i),
    .B(_011_),
    .C(_017_));
 sg13g2_nand3_1 _168_ (.B(_011_),
    .C(_017_),
    .A(ena_i),
    .Y(_041_));
 sg13g2_nor2_1 _169_ (.A(_037_),
    .B(_041_),
    .Y(output_o[161]));
 sg13g2_nand2_1 _170_ (.Y(output_no[161]),
    .A(_036_),
    .B(_040_));
 sg13g2_and3_1 _171_ (.X(_042_),
    .A(ena_i),
    .B(_011_),
    .C(_019_));
 sg13g2_nand3_1 _172_ (.B(_011_),
    .C(_019_),
    .A(ena_i),
    .Y(_043_));
 sg13g2_nor2_1 _173_ (.A(_037_),
    .B(_043_),
    .Y(output_o[162]));
 sg13g2_nand2_1 _174_ (.Y(output_no[162]),
    .A(_036_),
    .B(_042_));
 sg13g2_and3_1 _175_ (.X(_044_),
    .A(ena_i),
    .B(_006_),
    .C(_011_));
 sg13g2_nand3_1 _176_ (.B(_006_),
    .C(_011_),
    .A(ena_i),
    .Y(_045_));
 sg13g2_nor2_1 _177_ (.A(_037_),
    .B(_045_),
    .Y(output_o[163]));
 sg13g2_nand2_1 _178_ (.Y(output_no[163]),
    .A(_036_),
    .B(_044_));
 sg13g2_and3_1 _179_ (.X(_046_),
    .A(ena_i),
    .B(_012_),
    .C(_022_));
 sg13g2_nand3_1 _180_ (.B(_012_),
    .C(_022_),
    .A(ena_i),
    .Y(_047_));
 sg13g2_nor2_1 _181_ (.A(_037_),
    .B(_047_),
    .Y(output_o[164]));
 sg13g2_nand2_1 _182_ (.Y(output_no[164]),
    .A(_036_),
    .B(_046_));
 sg13g2_and3_1 _183_ (.X(_048_),
    .A(ena_i),
    .B(_017_),
    .C(_022_));
 sg13g2_nand3_1 _184_ (.B(_017_),
    .C(_022_),
    .A(ena_i),
    .Y(_049_));
 sg13g2_nor2_1 _185_ (.A(_037_),
    .B(_049_),
    .Y(output_o[165]));
 sg13g2_nand2_1 _186_ (.Y(output_no[165]),
    .A(_036_),
    .B(_048_));
 sg13g2_and3_1 _187_ (.X(_050_),
    .A(ena_i),
    .B(_019_),
    .C(_022_));
 sg13g2_nand3_1 _188_ (.B(_019_),
    .C(_022_),
    .A(ena_i),
    .Y(_051_));
 sg13g2_nor2_1 _189_ (.A(_037_),
    .B(_051_),
    .Y(output_o[166]));
 sg13g2_nand2_1 _190_ (.Y(output_no[166]),
    .A(_036_),
    .B(_050_));
 sg13g2_and3_1 _191_ (.X(_052_),
    .A(ena_i),
    .B(_006_),
    .C(_022_));
 sg13g2_nand3_1 _192_ (.B(_006_),
    .C(_022_),
    .A(ena_i),
    .Y(_053_));
 sg13g2_nor2_1 _193_ (.A(_037_),
    .B(_053_),
    .Y(output_o[167]));
 sg13g2_nand2_1 _194_ (.Y(output_no[167]),
    .A(_036_),
    .B(_052_));
 sg13g2_and3_1 _195_ (.X(_054_),
    .A(ena_i),
    .B(_012_),
    .C(_027_));
 sg13g2_nand3_1 _196_ (.B(_012_),
    .C(_027_),
    .A(ena_i),
    .Y(_055_));
 sg13g2_nor2_1 _197_ (.A(_037_),
    .B(_055_),
    .Y(output_o[168]));
 sg13g2_nand2_1 _198_ (.Y(output_no[168]),
    .A(_036_),
    .B(_054_));
 sg13g2_and3_1 _199_ (.X(_056_),
    .A(ena_i),
    .B(_017_),
    .C(_027_));
 sg13g2_nand3_1 _200_ (.B(_017_),
    .C(_027_),
    .A(ena_i),
    .Y(_057_));
 sg13g2_nor2_1 _201_ (.A(_037_),
    .B(_057_),
    .Y(output_o[169]));
 sg13g2_nand2_1 _202_ (.Y(output_no[169]),
    .A(_036_),
    .B(_056_));
 sg13g2_and3_1 _203_ (.X(_058_),
    .A(ena_i),
    .B(_019_),
    .C(_027_));
 sg13g2_nand3_1 _204_ (.B(_019_),
    .C(_027_),
    .A(ena_i),
    .Y(_059_));
 sg13g2_nor2_1 _205_ (.A(_037_),
    .B(_059_),
    .Y(output_o[170]));
 sg13g2_nand2_1 _206_ (.Y(output_no[170]),
    .A(_036_),
    .B(_058_));
 sg13g2_and3_1 _207_ (.X(_060_),
    .A(ena_i),
    .B(_006_),
    .C(_027_));
 sg13g2_nand3_1 _208_ (.B(_006_),
    .C(_027_),
    .A(ena_i),
    .Y(_061_));
 sg13g2_nor2_1 _209_ (.A(_037_),
    .B(_061_),
    .Y(output_o[171]));
 sg13g2_nand2_1 _210_ (.Y(output_no[171]),
    .A(_036_),
    .B(_060_));
 sg13g2_and3_1 _211_ (.X(_062_),
    .A(ena_i),
    .B(_005_),
    .C(_012_));
 sg13g2_nand3_1 _212_ (.B(_005_),
    .C(_012_),
    .A(ena_i),
    .Y(_063_));
 sg13g2_nor2_1 _213_ (.A(_037_),
    .B(_063_),
    .Y(output_o[172]));
 sg13g2_nand2_1 _214_ (.Y(output_no[172]),
    .A(_036_),
    .B(_062_));
 sg13g2_and3_1 _215_ (.X(_064_),
    .A(ena_i),
    .B(_005_),
    .C(_017_));
 sg13g2_nand3_1 _216_ (.B(_005_),
    .C(_017_),
    .A(ena_i),
    .Y(_065_));
 sg13g2_nor2_1 _217_ (.A(_037_),
    .B(_065_),
    .Y(output_o[173]));
 sg13g2_nand2_1 _218_ (.Y(output_no[173]),
    .A(_036_),
    .B(_064_));
 sg13g2_and3_1 _219_ (.X(_066_),
    .A(ena_i),
    .B(_005_),
    .C(_019_));
 sg13g2_nand3_1 _220_ (.B(_005_),
    .C(_019_),
    .A(ena_i),
    .Y(_067_));
 sg13g2_nor2_1 _221_ (.A(_037_),
    .B(_067_),
    .Y(output_o[174]));
 sg13g2_nand2_1 _222_ (.Y(output_no[174]),
    .A(_036_),
    .B(_066_));
 sg13g2_and2_1 _223_ (.A(ena_i),
    .B(_007_),
    .X(_068_));
 sg13g2_nand2_1 _224_ (.Y(_069_),
    .A(ena_i),
    .B(_007_));
 sg13g2_nor2_1 _225_ (.A(_037_),
    .B(_069_),
    .Y(output_o[175]));
 sg13g2_nand2_1 _226_ (.Y(output_no[175]),
    .A(_036_),
    .B(_068_));
 sg13g2_nor2_1 _227_ (.A(input_ni[4]),
    .B(input_ni[5]),
    .Y(_070_));
 sg13g2_and2_1 _228_ (.A(_008_),
    .B(_070_),
    .X(_071_));
 sg13g2_nand2_1 _229_ (.Y(_072_),
    .A(_008_),
    .B(_070_));
 sg13g2_nor2_1 _230_ (.A(_039_),
    .B(_072_),
    .Y(output_o[176]));
 sg13g2_nand2_1 _231_ (.Y(output_no[176]),
    .A(_038_),
    .B(_071_));
 sg13g2_nor2_1 _232_ (.A(_041_),
    .B(_072_),
    .Y(output_o[177]));
 sg13g2_nand2_1 _233_ (.Y(output_no[177]),
    .A(_040_),
    .B(_071_));
 sg13g2_nor2_1 _234_ (.A(_043_),
    .B(_072_),
    .Y(output_o[178]));
 sg13g2_nand2_1 _235_ (.Y(output_no[178]),
    .A(_042_),
    .B(_071_));
 sg13g2_nor2_1 _236_ (.A(_045_),
    .B(_072_),
    .Y(output_o[179]));
 sg13g2_nand2_1 _237_ (.Y(output_no[179]),
    .A(_044_),
    .B(_071_));
 sg13g2_nor2_1 _238_ (.A(_047_),
    .B(_072_),
    .Y(output_o[180]));
 sg13g2_nand2_1 _239_ (.Y(output_no[180]),
    .A(_046_),
    .B(_071_));
 sg13g2_nor2_1 _240_ (.A(_049_),
    .B(_072_),
    .Y(output_o[181]));
 sg13g2_nand2_1 _241_ (.Y(output_no[181]),
    .A(_048_),
    .B(_071_));
 sg13g2_nor2_1 _242_ (.A(_051_),
    .B(_072_),
    .Y(output_o[182]));
 sg13g2_nand2_1 _243_ (.Y(output_no[182]),
    .A(_050_),
    .B(_071_));
 sg13g2_nor2_1 _244_ (.A(_053_),
    .B(_072_),
    .Y(output_o[183]));
 sg13g2_nand2_1 _245_ (.Y(output_no[183]),
    .A(_052_),
    .B(_071_));
 sg13g2_nor2_1 _246_ (.A(_055_),
    .B(_072_),
    .Y(output_o[184]));
 sg13g2_nand2_1 _247_ (.Y(output_no[184]),
    .A(_054_),
    .B(_071_));
 sg13g2_nor2_1 _248_ (.A(_057_),
    .B(_072_),
    .Y(output_o[185]));
 sg13g2_nand2_1 _249_ (.Y(output_no[185]),
    .A(_056_),
    .B(_071_));
 sg13g2_nor2_1 _250_ (.A(_059_),
    .B(_072_),
    .Y(output_o[186]));
 sg13g2_nand2_1 _251_ (.Y(output_no[186]),
    .A(_058_),
    .B(_071_));
 sg13g2_nor2_1 _252_ (.A(_061_),
    .B(_072_),
    .Y(output_o[187]));
 sg13g2_nand2_1 _253_ (.Y(output_no[187]),
    .A(_060_),
    .B(_071_));
 sg13g2_nor2_1 _254_ (.A(_063_),
    .B(_072_),
    .Y(output_o[188]));
 sg13g2_nand2_1 _255_ (.Y(output_no[188]),
    .A(_062_),
    .B(_071_));
 sg13g2_nor2_1 _256_ (.A(_065_),
    .B(_072_),
    .Y(output_o[189]));
 sg13g2_nand2_1 _257_ (.Y(output_no[189]),
    .A(_064_),
    .B(_071_));
 sg13g2_nor2_1 _258_ (.A(_067_),
    .B(_072_),
    .Y(output_o[190]));
 sg13g2_nand2_1 _259_ (.Y(output_no[190]),
    .A(_066_),
    .B(_071_));
 sg13g2_nor2_1 _260_ (.A(_069_),
    .B(_072_),
    .Y(output_o[191]));
 sg13g2_nand2_1 _261_ (.Y(output_no[191]),
    .A(_068_),
    .B(_071_));
 sg13g2_nor2_1 _262_ (.A(input_ni[7]),
    .B(input_ni[6]),
    .Y(_073_));
 sg13g2_and3_1 _263_ (.X(_074_),
    .A(input_ni[4]),
    .B(input_ni[5]),
    .C(_073_));
 sg13g2_nand3_1 _264_ (.B(input_ni[5]),
    .C(_073_),
    .A(input_ni[4]),
    .Y(_075_));
 sg13g2_nor2_1 _265_ (.A(_039_),
    .B(_075_),
    .Y(output_o[192]));
 sg13g2_nand2_1 _266_ (.Y(output_no[192]),
    .A(_038_),
    .B(_074_));
 sg13g2_nor2_1 _267_ (.A(_041_),
    .B(_075_),
    .Y(output_o[193]));
 sg13g2_nand2_1 _268_ (.Y(output_no[193]),
    .A(_040_),
    .B(_074_));
 sg13g2_nor2_1 _269_ (.A(_043_),
    .B(_075_),
    .Y(output_o[194]));
 sg13g2_nand2_1 _270_ (.Y(output_no[194]),
    .A(_042_),
    .B(_074_));
 sg13g2_nor2_1 _271_ (.A(_045_),
    .B(_075_),
    .Y(output_o[195]));
 sg13g2_nand2_1 _272_ (.Y(output_no[195]),
    .A(_044_),
    .B(_074_));
 sg13g2_nor2_1 _273_ (.A(_047_),
    .B(_075_),
    .Y(output_o[196]));
 sg13g2_nand2_1 _274_ (.Y(output_no[196]),
    .A(_046_),
    .B(_074_));
 sg13g2_nor2_1 _275_ (.A(_049_),
    .B(_075_),
    .Y(output_o[197]));
 sg13g2_nand2_1 _276_ (.Y(output_no[197]),
    .A(_048_),
    .B(_074_));
 sg13g2_nor2_1 _277_ (.A(_051_),
    .B(_075_),
    .Y(output_o[198]));
 sg13g2_nand2_1 _278_ (.Y(output_no[198]),
    .A(_050_),
    .B(_074_));
 sg13g2_nor2_1 _279_ (.A(_053_),
    .B(_075_),
    .Y(output_o[199]));
 sg13g2_nand2_1 _280_ (.Y(output_no[199]),
    .A(_052_),
    .B(_074_));
 sg13g2_nor2_1 _281_ (.A(_055_),
    .B(_075_),
    .Y(output_o[200]));
 sg13g2_nand2_1 _282_ (.Y(output_no[200]),
    .A(_054_),
    .B(_074_));
 sg13g2_nor2_1 _283_ (.A(_057_),
    .B(_075_),
    .Y(output_o[201]));
 sg13g2_nand2_1 _284_ (.Y(output_no[201]),
    .A(_056_),
    .B(_074_));
 sg13g2_nor2_1 _285_ (.A(_059_),
    .B(_075_),
    .Y(output_o[202]));
 sg13g2_nand2_1 _286_ (.Y(output_no[202]),
    .A(_058_),
    .B(_074_));
 sg13g2_nor2_1 _287_ (.A(_061_),
    .B(_075_),
    .Y(output_o[203]));
 sg13g2_nand2_1 _288_ (.Y(output_no[203]),
    .A(_060_),
    .B(_074_));
 sg13g2_nor2_1 _289_ (.A(_063_),
    .B(_075_),
    .Y(output_o[204]));
 sg13g2_nand2_1 _290_ (.Y(output_no[204]),
    .A(_062_),
    .B(_074_));
 sg13g2_nor2_1 _291_ (.A(_065_),
    .B(_075_),
    .Y(output_o[205]));
 sg13g2_nand2_1 _292_ (.Y(output_no[205]),
    .A(_064_),
    .B(_074_));
 sg13g2_nor2_1 _293_ (.A(_067_),
    .B(_075_),
    .Y(output_o[206]));
 sg13g2_nand2_1 _294_ (.Y(output_no[206]),
    .A(_066_),
    .B(_074_));
 sg13g2_nor2_1 _295_ (.A(_069_),
    .B(_075_),
    .Y(output_o[207]));
 sg13g2_nand2_1 _296_ (.Y(output_no[207]),
    .A(_068_),
    .B(_074_));
 sg13g2_and2_1 _297_ (.A(_014_),
    .B(_073_),
    .X(_076_));
 sg13g2_nand2_1 _298_ (.Y(_077_),
    .A(_014_),
    .B(_073_));
 sg13g2_nor2_1 _299_ (.A(_039_),
    .B(_077_),
    .Y(output_o[208]));
 sg13g2_nand2_1 _300_ (.Y(output_no[208]),
    .A(_038_),
    .B(_076_));
 sg13g2_nor2_1 _301_ (.A(_041_),
    .B(_077_),
    .Y(output_o[209]));
 sg13g2_nand2_1 _302_ (.Y(output_no[209]),
    .A(_040_),
    .B(_076_));
 sg13g2_nor2_1 _303_ (.A(_043_),
    .B(_077_),
    .Y(output_o[210]));
 sg13g2_nand2_1 _304_ (.Y(output_no[210]),
    .A(_042_),
    .B(_076_));
 sg13g2_nor2_1 _305_ (.A(_045_),
    .B(_077_),
    .Y(output_o[211]));
 sg13g2_nand2_1 _306_ (.Y(output_no[211]),
    .A(_044_),
    .B(_076_));
 sg13g2_nor2_1 _307_ (.A(_047_),
    .B(_077_),
    .Y(output_o[212]));
 sg13g2_nand2_1 _308_ (.Y(output_no[212]),
    .A(_046_),
    .B(_076_));
 sg13g2_nor2_1 _309_ (.A(_049_),
    .B(_077_),
    .Y(output_o[213]));
 sg13g2_nand2_1 _310_ (.Y(output_no[213]),
    .A(_048_),
    .B(_076_));
 sg13g2_nor2_1 _311_ (.A(_051_),
    .B(_077_),
    .Y(output_o[214]));
 sg13g2_nand2_1 _312_ (.Y(output_no[214]),
    .A(_050_),
    .B(_076_));
 sg13g2_nor2_1 _313_ (.A(_053_),
    .B(_077_),
    .Y(output_o[215]));
 sg13g2_nand2_1 _314_ (.Y(output_no[215]),
    .A(_052_),
    .B(_076_));
 sg13g2_nor2_1 _315_ (.A(_055_),
    .B(_077_),
    .Y(output_o[216]));
 sg13g2_nand2_1 _316_ (.Y(output_no[216]),
    .A(_054_),
    .B(_076_));
 sg13g2_nor2_1 _317_ (.A(_057_),
    .B(_077_),
    .Y(output_o[217]));
 sg13g2_nand2_1 _318_ (.Y(output_no[217]),
    .A(_056_),
    .B(_076_));
 sg13g2_nor2_1 _319_ (.A(_059_),
    .B(_077_),
    .Y(output_o[218]));
 sg13g2_nand2_1 _320_ (.Y(output_no[218]),
    .A(_058_),
    .B(_076_));
 sg13g2_nor2_1 _321_ (.A(_061_),
    .B(_077_),
    .Y(output_o[219]));
 sg13g2_nand2_1 _322_ (.Y(output_no[219]),
    .A(_060_),
    .B(_076_));
 sg13g2_nor2_1 _323_ (.A(_063_),
    .B(_077_),
    .Y(output_o[220]));
 sg13g2_nand2_1 _324_ (.Y(output_no[220]),
    .A(_062_),
    .B(_076_));
 sg13g2_nor2_1 _325_ (.A(_065_),
    .B(_077_),
    .Y(output_o[221]));
 sg13g2_nand2_1 _326_ (.Y(output_no[221]),
    .A(_064_),
    .B(_076_));
 sg13g2_nor2_1 _327_ (.A(_067_),
    .B(_077_),
    .Y(output_o[222]));
 sg13g2_nand2_1 _328_ (.Y(output_no[222]),
    .A(_066_),
    .B(_076_));
 sg13g2_nor2_1 _329_ (.A(_069_),
    .B(_077_),
    .Y(output_o[223]));
 sg13g2_nand2_1 _330_ (.Y(output_no[223]),
    .A(_068_),
    .B(_076_));
 sg13g2_and2_1 _331_ (.A(_035_),
    .B(_073_),
    .X(_078_));
 sg13g2_nand2_1 _332_ (.Y(_079_),
    .A(_035_),
    .B(_073_));
 sg13g2_nor2_1 _333_ (.A(_039_),
    .B(_079_),
    .Y(output_o[224]));
 sg13g2_nand2_1 _334_ (.Y(output_no[224]),
    .A(_038_),
    .B(_078_));
 sg13g2_nor2_1 _335_ (.A(_041_),
    .B(_079_),
    .Y(output_o[225]));
 sg13g2_nand2_1 _336_ (.Y(output_no[225]),
    .A(_040_),
    .B(_078_));
 sg13g2_nor2_1 _337_ (.A(_043_),
    .B(_079_),
    .Y(output_o[226]));
 sg13g2_nand2_1 _338_ (.Y(output_no[226]),
    .A(_042_),
    .B(_078_));
 sg13g2_nor2_1 _339_ (.A(_045_),
    .B(_079_),
    .Y(output_o[227]));
 sg13g2_nand2_1 _340_ (.Y(output_no[227]),
    .A(_044_),
    .B(_078_));
 sg13g2_nor2_1 _341_ (.A(_047_),
    .B(_079_),
    .Y(output_o[228]));
 sg13g2_nand2_1 _342_ (.Y(output_no[228]),
    .A(_046_),
    .B(_078_));
 sg13g2_nor2_1 _343_ (.A(_049_),
    .B(_079_),
    .Y(output_o[229]));
 sg13g2_nand2_1 _344_ (.Y(output_no[229]),
    .A(_048_),
    .B(_078_));
 sg13g2_nor2_1 _345_ (.A(_051_),
    .B(_079_),
    .Y(output_o[230]));
 sg13g2_nand2_1 _346_ (.Y(output_no[230]),
    .A(_050_),
    .B(_078_));
 sg13g2_nor2_1 _347_ (.A(_053_),
    .B(_079_),
    .Y(output_o[231]));
 sg13g2_nand2_1 _348_ (.Y(output_no[231]),
    .A(_052_),
    .B(_078_));
 sg13g2_nor2_1 _349_ (.A(_055_),
    .B(_079_),
    .Y(output_o[232]));
 sg13g2_nand2_1 _350_ (.Y(output_no[232]),
    .A(_054_),
    .B(_078_));
 sg13g2_nor2_1 _351_ (.A(_057_),
    .B(_079_),
    .Y(output_o[233]));
 sg13g2_nand2_1 _352_ (.Y(output_no[233]),
    .A(_056_),
    .B(_078_));
 sg13g2_nor2_1 _353_ (.A(_059_),
    .B(_079_),
    .Y(output_o[234]));
 sg13g2_nand2_1 _354_ (.Y(output_no[234]),
    .A(_058_),
    .B(_078_));
 sg13g2_nor2_1 _355_ (.A(_061_),
    .B(_079_),
    .Y(output_o[235]));
 sg13g2_nand2_1 _356_ (.Y(output_no[235]),
    .A(_060_),
    .B(_078_));
 sg13g2_nor2_1 _357_ (.A(_063_),
    .B(_079_),
    .Y(output_o[236]));
 sg13g2_nand2_1 _358_ (.Y(output_no[236]),
    .A(_062_),
    .B(_078_));
 sg13g2_nor2_1 _359_ (.A(_065_),
    .B(_079_),
    .Y(output_o[237]));
 sg13g2_nand2_1 _360_ (.Y(output_no[237]),
    .A(_064_),
    .B(_078_));
 sg13g2_nor2_1 _361_ (.A(_067_),
    .B(_079_),
    .Y(output_o[238]));
 sg13g2_nand2_1 _362_ (.Y(output_no[238]),
    .A(_066_),
    .B(_078_));
 sg13g2_nor2_1 _363_ (.A(_069_),
    .B(_079_),
    .Y(output_o[239]));
 sg13g2_nand2_1 _364_ (.Y(output_no[239]),
    .A(_068_),
    .B(_078_));
 sg13g2_and2_1 _365_ (.A(_070_),
    .B(_073_),
    .X(_080_));
 sg13g2_nand2_1 _366_ (.Y(_081_),
    .A(_070_),
    .B(_073_));
 sg13g2_nor2_1 _367_ (.A(_039_),
    .B(_081_),
    .Y(output_o[240]));
 sg13g2_nand2_1 _368_ (.Y(output_no[240]),
    .A(_038_),
    .B(_080_));
 sg13g2_nor2_1 _369_ (.A(_041_),
    .B(_081_),
    .Y(output_o[241]));
 sg13g2_nand2_1 _370_ (.Y(output_no[241]),
    .A(_040_),
    .B(_080_));
 sg13g2_nor2_1 _371_ (.A(_043_),
    .B(_081_),
    .Y(output_o[242]));
 sg13g2_nand2_1 _372_ (.Y(output_no[242]),
    .A(_042_),
    .B(_080_));
 sg13g2_nor2_1 _373_ (.A(_045_),
    .B(_081_),
    .Y(output_o[243]));
 sg13g2_nand2_1 _374_ (.Y(output_no[243]),
    .A(_044_),
    .B(_080_));
 sg13g2_nor2_1 _375_ (.A(_047_),
    .B(_081_),
    .Y(output_o[244]));
 sg13g2_nand2_1 _376_ (.Y(output_no[244]),
    .A(_046_),
    .B(_080_));
 sg13g2_nor2_1 _377_ (.A(_049_),
    .B(_081_),
    .Y(output_o[245]));
 sg13g2_nand2_1 _378_ (.Y(output_no[245]),
    .A(_048_),
    .B(_080_));
 sg13g2_nor2_1 _379_ (.A(_051_),
    .B(_081_),
    .Y(output_o[246]));
 sg13g2_nand2_1 _380_ (.Y(output_no[246]),
    .A(_050_),
    .B(_080_));
 sg13g2_nor2_1 _381_ (.A(_053_),
    .B(_081_),
    .Y(output_o[247]));
 sg13g2_nand2_1 _382_ (.Y(output_no[247]),
    .A(_052_),
    .B(_080_));
 sg13g2_nor2_1 _383_ (.A(_055_),
    .B(_081_),
    .Y(output_o[248]));
 sg13g2_nand2_1 _384_ (.Y(output_no[248]),
    .A(_054_),
    .B(_080_));
 sg13g2_nor2_1 _385_ (.A(_057_),
    .B(_081_),
    .Y(output_o[249]));
 sg13g2_nand2_1 _386_ (.Y(output_no[249]),
    .A(_056_),
    .B(_080_));
 sg13g2_nor2_1 _387_ (.A(_059_),
    .B(_081_),
    .Y(output_o[250]));
 sg13g2_nand2_1 _388_ (.Y(output_no[250]),
    .A(_058_),
    .B(_080_));
 sg13g2_nor2_1 _389_ (.A(_061_),
    .B(_081_),
    .Y(output_o[251]));
 sg13g2_nand2_1 _390_ (.Y(output_no[251]),
    .A(_060_),
    .B(_080_));
 sg13g2_nor2_1 _391_ (.A(_063_),
    .B(_081_),
    .Y(output_o[252]));
 sg13g2_nand2_1 _392_ (.Y(output_no[252]),
    .A(_062_),
    .B(_080_));
 sg13g2_nor2_1 _393_ (.A(_065_),
    .B(_081_),
    .Y(output_o[253]));
 sg13g2_nand2_1 _394_ (.Y(output_no[253]),
    .A(_064_),
    .B(_080_));
 sg13g2_nor2_1 _395_ (.A(_067_),
    .B(_081_),
    .Y(output_o[254]));
 sg13g2_nand2_1 _396_ (.Y(output_no[254]),
    .A(_066_),
    .B(_080_));
 sg13g2_nor2_1 _397_ (.A(_069_),
    .B(_081_),
    .Y(output_o[255]));
 sg13g2_nand2_1 _398_ (.Y(output_no[255]),
    .A(_068_),
    .B(_080_));
 sg13g2_and3_1 _399_ (.X(_082_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_014_));
 sg13g2_nand3_1 _400_ (.B(input_ni[6]),
    .C(_014_),
    .A(input_ni[7]),
    .Y(_083_));
 sg13g2_nor2_1 _401_ (.A(_039_),
    .B(_083_),
    .Y(output_o[16]));
 sg13g2_nand2_1 _402_ (.Y(output_no[16]),
    .A(_038_),
    .B(_082_));
 sg13g2_nor2_1 _403_ (.A(_041_),
    .B(_083_),
    .Y(output_o[17]));
 sg13g2_nand2_1 _404_ (.Y(output_no[17]),
    .A(_040_),
    .B(_082_));
 sg13g2_nor2_1 _405_ (.A(_043_),
    .B(_083_),
    .Y(output_o[18]));
 sg13g2_nand2_1 _406_ (.Y(output_no[18]),
    .A(_042_),
    .B(_082_));
 sg13g2_nor2_1 _407_ (.A(_045_),
    .B(_083_),
    .Y(output_o[19]));
 sg13g2_nand2_1 _408_ (.Y(output_no[19]),
    .A(_044_),
    .B(_082_));
 sg13g2_nor2_1 _409_ (.A(_047_),
    .B(_083_),
    .Y(output_o[20]));
 sg13g2_nand2_1 _410_ (.Y(output_no[20]),
    .A(_046_),
    .B(_082_));
 sg13g2_nor2_1 _411_ (.A(_049_),
    .B(_083_),
    .Y(output_o[21]));
 sg13g2_nand2_1 _412_ (.Y(output_no[21]),
    .A(_048_),
    .B(_082_));
 sg13g2_nor2_1 _413_ (.A(_051_),
    .B(_083_),
    .Y(output_o[22]));
 sg13g2_nand2_1 _414_ (.Y(output_no[22]),
    .A(_050_),
    .B(_082_));
 sg13g2_nor2_1 _415_ (.A(_053_),
    .B(_083_),
    .Y(output_o[23]));
 sg13g2_nand2_1 _416_ (.Y(output_no[23]),
    .A(_052_),
    .B(_082_));
 sg13g2_nor2_1 _417_ (.A(_055_),
    .B(_083_),
    .Y(output_o[24]));
 sg13g2_nand2_1 _418_ (.Y(output_no[24]),
    .A(_054_),
    .B(_082_));
 sg13g2_nor2_1 _419_ (.A(_057_),
    .B(_083_),
    .Y(output_o[25]));
 sg13g2_nand2_1 _420_ (.Y(output_no[25]),
    .A(_056_),
    .B(_082_));
 sg13g2_nor2_1 _421_ (.A(_059_),
    .B(_083_),
    .Y(output_o[26]));
 sg13g2_nand2_1 _422_ (.Y(output_no[26]),
    .A(_058_),
    .B(_082_));
 sg13g2_nor2_1 _423_ (.A(_061_),
    .B(_083_),
    .Y(output_o[27]));
 sg13g2_nand2_1 _424_ (.Y(output_no[27]),
    .A(_060_),
    .B(_082_));
 sg13g2_nor2_1 _425_ (.A(_063_),
    .B(_083_),
    .Y(output_o[28]));
 sg13g2_nand2_1 _426_ (.Y(output_no[28]),
    .A(_062_),
    .B(_082_));
 sg13g2_nor2_1 _427_ (.A(_065_),
    .B(_083_),
    .Y(output_o[29]));
 sg13g2_nand2_1 _428_ (.Y(output_no[29]),
    .A(_064_),
    .B(_082_));
 sg13g2_nor2_1 _429_ (.A(_067_),
    .B(_083_),
    .Y(output_o[30]));
 sg13g2_nand2_1 _430_ (.Y(output_no[30]),
    .A(_066_),
    .B(_082_));
 sg13g2_nor2_1 _431_ (.A(_069_),
    .B(_083_),
    .Y(output_o[31]));
 sg13g2_nand2_1 _432_ (.Y(output_no[31]),
    .A(_068_),
    .B(_082_));
 sg13g2_and3_1 _433_ (.X(_084_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_035_));
 sg13g2_nand3_1 _434_ (.B(input_ni[6]),
    .C(_035_),
    .A(input_ni[7]),
    .Y(_085_));
 sg13g2_nor2_1 _435_ (.A(_039_),
    .B(_085_),
    .Y(output_o[32]));
 sg13g2_nand2_1 _436_ (.Y(output_no[32]),
    .A(_038_),
    .B(_084_));
 sg13g2_nor2_1 _437_ (.A(_041_),
    .B(_085_),
    .Y(output_o[33]));
 sg13g2_nand2_1 _438_ (.Y(output_no[33]),
    .A(_040_),
    .B(_084_));
 sg13g2_nor2_1 _439_ (.A(_043_),
    .B(_085_),
    .Y(output_o[34]));
 sg13g2_nand2_1 _440_ (.Y(output_no[34]),
    .A(_042_),
    .B(_084_));
 sg13g2_nor2_1 _441_ (.A(_045_),
    .B(_085_),
    .Y(output_o[35]));
 sg13g2_nand2_1 _442_ (.Y(output_no[35]),
    .A(_044_),
    .B(_084_));
 sg13g2_nor2_1 _443_ (.A(_047_),
    .B(_085_),
    .Y(output_o[36]));
 sg13g2_nand2_1 _444_ (.Y(output_no[36]),
    .A(_046_),
    .B(_084_));
 sg13g2_nor2_1 _445_ (.A(_049_),
    .B(_085_),
    .Y(output_o[37]));
 sg13g2_nand2_1 _446_ (.Y(output_no[37]),
    .A(_048_),
    .B(_084_));
 sg13g2_nor2_1 _447_ (.A(_051_),
    .B(_085_),
    .Y(output_o[38]));
 sg13g2_nand2_1 _448_ (.Y(output_no[38]),
    .A(_050_),
    .B(_084_));
 sg13g2_nor2_1 _449_ (.A(_053_),
    .B(_085_),
    .Y(output_o[39]));
 sg13g2_nand2_1 _450_ (.Y(output_no[39]),
    .A(_052_),
    .B(_084_));
 sg13g2_nor2_1 _451_ (.A(_055_),
    .B(_085_),
    .Y(output_o[40]));
 sg13g2_nand2_1 _452_ (.Y(output_no[40]),
    .A(_054_),
    .B(_084_));
 sg13g2_nor2_1 _453_ (.A(_057_),
    .B(_085_),
    .Y(output_o[41]));
 sg13g2_nand2_1 _454_ (.Y(output_no[41]),
    .A(_056_),
    .B(_084_));
 sg13g2_nor2_1 _455_ (.A(_059_),
    .B(_085_),
    .Y(output_o[42]));
 sg13g2_nand2_1 _456_ (.Y(output_no[42]),
    .A(_058_),
    .B(_084_));
 sg13g2_nor2_1 _457_ (.A(_061_),
    .B(_085_),
    .Y(output_o[43]));
 sg13g2_nand2_1 _458_ (.Y(output_no[43]),
    .A(_060_),
    .B(_084_));
 sg13g2_nor2_1 _459_ (.A(_063_),
    .B(_085_),
    .Y(output_o[44]));
 sg13g2_nand2_1 _460_ (.Y(output_no[44]),
    .A(_062_),
    .B(_084_));
 sg13g2_nor2_1 _461_ (.A(_065_),
    .B(_085_),
    .Y(output_o[45]));
 sg13g2_nand2_1 _462_ (.Y(output_no[45]),
    .A(_064_),
    .B(_084_));
 sg13g2_nor2_1 _463_ (.A(_067_),
    .B(_085_),
    .Y(output_o[46]));
 sg13g2_nand2_1 _464_ (.Y(output_no[46]),
    .A(_066_),
    .B(_084_));
 sg13g2_nor2_1 _465_ (.A(_069_),
    .B(_085_),
    .Y(output_o[47]));
 sg13g2_nand2_1 _466_ (.Y(output_no[47]),
    .A(_068_),
    .B(_084_));
 sg13g2_and3_1 _467_ (.X(_086_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_070_));
 sg13g2_nand3_1 _468_ (.B(input_ni[6]),
    .C(_070_),
    .A(input_ni[7]),
    .Y(_087_));
 sg13g2_nor2_1 _469_ (.A(_039_),
    .B(_087_),
    .Y(output_o[48]));
 sg13g2_nand2_1 _470_ (.Y(output_no[48]),
    .A(_038_),
    .B(_086_));
 sg13g2_nor2_1 _471_ (.A(_041_),
    .B(_087_),
    .Y(output_o[49]));
 sg13g2_nand2_1 _472_ (.Y(output_no[49]),
    .A(_040_),
    .B(_086_));
 sg13g2_nor2_1 _473_ (.A(_043_),
    .B(_087_),
    .Y(output_o[50]));
 sg13g2_nand2_1 _474_ (.Y(output_no[50]),
    .A(_042_),
    .B(_086_));
 sg13g2_nor2_1 _475_ (.A(_045_),
    .B(_087_),
    .Y(output_o[51]));
 sg13g2_nand2_1 _476_ (.Y(output_no[51]),
    .A(_044_),
    .B(_086_));
 sg13g2_nor2_1 _477_ (.A(_047_),
    .B(_087_),
    .Y(output_o[52]));
 sg13g2_nand2_1 _478_ (.Y(output_no[52]),
    .A(_046_),
    .B(_086_));
 sg13g2_nor2_1 _479_ (.A(_049_),
    .B(_087_),
    .Y(output_o[53]));
 sg13g2_nand2_1 _480_ (.Y(output_no[53]),
    .A(_048_),
    .B(_086_));
 sg13g2_nor2_1 _481_ (.A(_051_),
    .B(_087_),
    .Y(output_o[54]));
 sg13g2_nand2_1 _482_ (.Y(output_no[54]),
    .A(_050_),
    .B(_086_));
 sg13g2_nor2_1 _483_ (.A(_053_),
    .B(_087_),
    .Y(output_o[55]));
 sg13g2_nand2_1 _484_ (.Y(output_no[55]),
    .A(_052_),
    .B(_086_));
 sg13g2_nor2_1 _485_ (.A(_055_),
    .B(_087_),
    .Y(output_o[56]));
 sg13g2_nand2_1 _486_ (.Y(output_no[56]),
    .A(_054_),
    .B(_086_));
 sg13g2_nor2_1 _487_ (.A(_057_),
    .B(_087_),
    .Y(output_o[57]));
 sg13g2_nand2_1 _488_ (.Y(output_no[57]),
    .A(_056_),
    .B(_086_));
 sg13g2_nor2_1 _489_ (.A(_059_),
    .B(_087_),
    .Y(output_o[58]));
 sg13g2_nand2_1 _490_ (.Y(output_no[58]),
    .A(_058_),
    .B(_086_));
 sg13g2_nor2_1 _491_ (.A(_061_),
    .B(_087_),
    .Y(output_o[59]));
 sg13g2_nand2_1 _492_ (.Y(output_no[59]),
    .A(_060_),
    .B(_086_));
 sg13g2_nor2_1 _493_ (.A(_063_),
    .B(_087_),
    .Y(output_o[60]));
 sg13g2_nand2_1 _494_ (.Y(output_no[60]),
    .A(_062_),
    .B(_086_));
 sg13g2_nor2_1 _495_ (.A(_065_),
    .B(_087_),
    .Y(output_o[61]));
 sg13g2_nand2_1 _496_ (.Y(output_no[61]),
    .A(_064_),
    .B(_086_));
 sg13g2_nor2_1 _497_ (.A(_067_),
    .B(_087_),
    .Y(output_o[62]));
 sg13g2_nand2_1 _498_ (.Y(output_no[62]),
    .A(_066_),
    .B(_086_));
 sg13g2_nor2_1 _499_ (.A(_069_),
    .B(_087_),
    .Y(output_o[63]));
 sg13g2_nand2_1 _500_ (.Y(output_no[63]),
    .A(_068_),
    .B(_086_));
 sg13g2_nand3_1 _501_ (.B(input_ni[5]),
    .C(input_ni[7]),
    .A(input_ni[4]),
    .Y(_088_));
 sg13g2_nor2_1 _502_ (.A(input_ni[6]),
    .B(_088_),
    .Y(_089_));
 sg13g2_nand2b_1 _503_ (.Y(_090_),
    .B(_004_),
    .A_N(_088_));
 sg13g2_nor2_1 _504_ (.A(_039_),
    .B(_090_),
    .Y(output_o[64]));
 sg13g2_nand2_1 _505_ (.Y(output_no[64]),
    .A(_038_),
    .B(_089_));
 sg13g2_nor2_1 _506_ (.A(_041_),
    .B(_090_),
    .Y(output_o[65]));
 sg13g2_nand2_1 _507_ (.Y(output_no[65]),
    .A(_040_),
    .B(_089_));
 sg13g2_nor2_1 _508_ (.A(_043_),
    .B(_090_),
    .Y(output_o[66]));
 sg13g2_nand2_1 _509_ (.Y(output_no[66]),
    .A(_042_),
    .B(_089_));
 sg13g2_nor2_1 _510_ (.A(_045_),
    .B(_090_),
    .Y(output_o[67]));
 sg13g2_nand2_1 _511_ (.Y(output_no[67]),
    .A(_044_),
    .B(_089_));
 sg13g2_nor2_1 _512_ (.A(_047_),
    .B(_090_),
    .Y(output_o[68]));
 sg13g2_nand2_1 _513_ (.Y(output_no[68]),
    .A(_046_),
    .B(_089_));
 sg13g2_nor2_1 _514_ (.A(_049_),
    .B(_090_),
    .Y(output_o[69]));
 sg13g2_nand2_1 _515_ (.Y(output_no[69]),
    .A(_048_),
    .B(_089_));
 sg13g2_nor2_1 _516_ (.A(_051_),
    .B(_090_),
    .Y(output_o[70]));
 sg13g2_nand2_1 _517_ (.Y(output_no[70]),
    .A(_050_),
    .B(_089_));
 sg13g2_nor2_1 _518_ (.A(_053_),
    .B(_090_),
    .Y(output_o[71]));
 sg13g2_nand2_1 _519_ (.Y(output_no[71]),
    .A(_052_),
    .B(_089_));
 sg13g2_nor2_1 _520_ (.A(_055_),
    .B(_090_),
    .Y(output_o[72]));
 sg13g2_nand2_1 _521_ (.Y(output_no[72]),
    .A(_054_),
    .B(_089_));
 sg13g2_nor2_1 _522_ (.A(_057_),
    .B(_090_),
    .Y(output_o[73]));
 sg13g2_nand2_1 _523_ (.Y(output_no[73]),
    .A(_056_),
    .B(_089_));
 sg13g2_nor2_1 _524_ (.A(_059_),
    .B(_090_),
    .Y(output_o[74]));
 sg13g2_nand2_1 _525_ (.Y(output_no[74]),
    .A(_058_),
    .B(_089_));
 sg13g2_nor2_1 _526_ (.A(_061_),
    .B(_090_),
    .Y(output_o[75]));
 sg13g2_nand2_1 _527_ (.Y(output_no[75]),
    .A(_060_),
    .B(_089_));
 sg13g2_nor2_1 _528_ (.A(_063_),
    .B(_090_),
    .Y(output_o[76]));
 sg13g2_nand2_1 _529_ (.Y(output_no[76]),
    .A(_062_),
    .B(_089_));
 sg13g2_nor2_1 _530_ (.A(_065_),
    .B(_090_),
    .Y(output_o[77]));
 sg13g2_nand2_1 _531_ (.Y(output_no[77]),
    .A(_064_),
    .B(_089_));
 sg13g2_nor2_1 _532_ (.A(_067_),
    .B(_090_),
    .Y(output_o[78]));
 sg13g2_nand2_1 _533_ (.Y(output_no[78]),
    .A(_066_),
    .B(_089_));
 sg13g2_nor2_1 _534_ (.A(_069_),
    .B(_090_),
    .Y(output_o[79]));
 sg13g2_nand2_1 _535_ (.Y(output_no[79]),
    .A(_068_),
    .B(_089_));
 sg13g2_and3_1 _536_ (.X(_091_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_014_));
 sg13g2_nand3_1 _537_ (.B(_004_),
    .C(_014_),
    .A(input_ni[7]),
    .Y(_092_));
 sg13g2_nor2_1 _538_ (.A(_039_),
    .B(_092_),
    .Y(output_o[80]));
 sg13g2_nand2_1 _539_ (.Y(output_no[80]),
    .A(_038_),
    .B(_091_));
 sg13g2_nor2_1 _540_ (.A(_041_),
    .B(_092_),
    .Y(output_o[81]));
 sg13g2_nand2_1 _541_ (.Y(output_no[81]),
    .A(_040_),
    .B(_091_));
 sg13g2_nor2_1 _542_ (.A(_043_),
    .B(_092_),
    .Y(output_o[82]));
 sg13g2_nand2_1 _543_ (.Y(output_no[82]),
    .A(_042_),
    .B(_091_));
 sg13g2_nor2_1 _544_ (.A(_045_),
    .B(_092_),
    .Y(output_o[83]));
 sg13g2_nand2_1 _545_ (.Y(output_no[83]),
    .A(_044_),
    .B(_091_));
 sg13g2_nor2_1 _546_ (.A(_047_),
    .B(_092_),
    .Y(output_o[84]));
 sg13g2_nand2_1 _547_ (.Y(output_no[84]),
    .A(_046_),
    .B(_091_));
 sg13g2_nor2_1 _548_ (.A(_049_),
    .B(_092_),
    .Y(output_o[85]));
 sg13g2_nand2_1 _549_ (.Y(output_no[85]),
    .A(_048_),
    .B(_091_));
 sg13g2_nor2_1 _550_ (.A(_051_),
    .B(_092_),
    .Y(output_o[86]));
 sg13g2_nand2_1 _551_ (.Y(output_no[86]),
    .A(_050_),
    .B(_091_));
 sg13g2_nor2_1 _552_ (.A(_053_),
    .B(_092_),
    .Y(output_o[87]));
 sg13g2_nand2_1 _553_ (.Y(output_no[87]),
    .A(_052_),
    .B(_091_));
 sg13g2_nor2_1 _554_ (.A(_055_),
    .B(_092_),
    .Y(output_o[88]));
 sg13g2_nand2_1 _555_ (.Y(output_no[88]),
    .A(_054_),
    .B(_091_));
 sg13g2_nor2_1 _556_ (.A(_057_),
    .B(_092_),
    .Y(output_o[89]));
 sg13g2_nand2_1 _557_ (.Y(output_no[89]),
    .A(_056_),
    .B(_091_));
 sg13g2_nor2_1 _558_ (.A(_059_),
    .B(_092_),
    .Y(output_o[90]));
 sg13g2_nand2_1 _559_ (.Y(output_no[90]),
    .A(_058_),
    .B(_091_));
 sg13g2_nor2_1 _560_ (.A(_061_),
    .B(_092_),
    .Y(output_o[91]));
 sg13g2_nand2_1 _561_ (.Y(output_no[91]),
    .A(_060_),
    .B(_091_));
 sg13g2_nor2_1 _562_ (.A(_063_),
    .B(_092_),
    .Y(output_o[92]));
 sg13g2_nand2_1 _563_ (.Y(output_no[92]),
    .A(_062_),
    .B(_091_));
 sg13g2_nor2_1 _564_ (.A(_065_),
    .B(_092_),
    .Y(output_o[93]));
 sg13g2_nand2_1 _565_ (.Y(output_no[93]),
    .A(_064_),
    .B(_091_));
 sg13g2_nor2_1 _566_ (.A(_067_),
    .B(_092_),
    .Y(output_o[94]));
 sg13g2_nand2_1 _567_ (.Y(output_no[94]),
    .A(_066_),
    .B(_091_));
 sg13g2_nor2_1 _568_ (.A(_069_),
    .B(_092_),
    .Y(output_o[95]));
 sg13g2_nand2_1 _569_ (.Y(output_no[95]),
    .A(_068_),
    .B(_091_));
 sg13g2_and3_1 _570_ (.X(_093_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_035_));
 sg13g2_nand3_1 _571_ (.B(_004_),
    .C(_035_),
    .A(input_ni[7]),
    .Y(_094_));
 sg13g2_nor2_1 _572_ (.A(_039_),
    .B(_094_),
    .Y(output_o[96]));
 sg13g2_nand2_1 _573_ (.Y(output_no[96]),
    .A(_038_),
    .B(_093_));
 sg13g2_nor2_1 _574_ (.A(_041_),
    .B(_094_),
    .Y(output_o[97]));
 sg13g2_nand2_1 _575_ (.Y(output_no[97]),
    .A(_040_),
    .B(_093_));
 sg13g2_nor2_1 _576_ (.A(_043_),
    .B(_094_),
    .Y(output_o[98]));
 sg13g2_nand2_1 _577_ (.Y(output_no[98]),
    .A(_042_),
    .B(_093_));
 sg13g2_nor2_1 _578_ (.A(_045_),
    .B(_094_),
    .Y(output_o[99]));
 sg13g2_nand2_1 _579_ (.Y(output_no[99]),
    .A(_044_),
    .B(_093_));
 sg13g2_nor2_1 _580_ (.A(_047_),
    .B(_094_),
    .Y(output_o[100]));
 sg13g2_nand2_1 _581_ (.Y(output_no[100]),
    .A(_046_),
    .B(_093_));
 sg13g2_nor2_1 _582_ (.A(_049_),
    .B(_094_),
    .Y(output_o[101]));
 sg13g2_nand2_1 _583_ (.Y(output_no[101]),
    .A(_048_),
    .B(_093_));
 sg13g2_nor2_1 _584_ (.A(_051_),
    .B(_094_),
    .Y(output_o[102]));
 sg13g2_nand2_1 _585_ (.Y(output_no[102]),
    .A(_050_),
    .B(_093_));
 sg13g2_nor2_1 _586_ (.A(_053_),
    .B(_094_),
    .Y(output_o[103]));
 sg13g2_nand2_1 _587_ (.Y(output_no[103]),
    .A(_052_),
    .B(_093_));
 sg13g2_nor2_1 _588_ (.A(_055_),
    .B(_094_),
    .Y(output_o[104]));
 sg13g2_nand2_1 _589_ (.Y(output_no[104]),
    .A(_054_),
    .B(_093_));
 sg13g2_nor2_1 _590_ (.A(_057_),
    .B(_094_),
    .Y(output_o[105]));
 sg13g2_nand2_1 _591_ (.Y(output_no[105]),
    .A(_056_),
    .B(_093_));
 sg13g2_nor2_1 _592_ (.A(_059_),
    .B(_094_),
    .Y(output_o[106]));
 sg13g2_nand2_1 _593_ (.Y(output_no[106]),
    .A(_058_),
    .B(_093_));
 sg13g2_nor2_1 _594_ (.A(_061_),
    .B(_094_),
    .Y(output_o[107]));
 sg13g2_nand2_1 _595_ (.Y(output_no[107]),
    .A(_060_),
    .B(_093_));
 sg13g2_nor2_1 _596_ (.A(_063_),
    .B(_094_),
    .Y(output_o[108]));
 sg13g2_nand2_1 _597_ (.Y(output_no[108]),
    .A(_062_),
    .B(_093_));
 sg13g2_nor2_1 _598_ (.A(_065_),
    .B(_094_),
    .Y(output_o[109]));
 sg13g2_nand2_1 _599_ (.Y(output_no[109]),
    .A(_064_),
    .B(_093_));
 sg13g2_nor2_1 _600_ (.A(_067_),
    .B(_094_),
    .Y(output_o[110]));
 sg13g2_nand2_1 _601_ (.Y(output_no[110]),
    .A(_066_),
    .B(_093_));
 sg13g2_nor2_1 _602_ (.A(_069_),
    .B(_094_),
    .Y(output_o[111]));
 sg13g2_nand2_1 _603_ (.Y(output_no[111]),
    .A(_068_),
    .B(_093_));
 sg13g2_and3_1 _604_ (.X(_000_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_070_));
 sg13g2_nand3_1 _605_ (.B(_004_),
    .C(_070_),
    .A(input_ni[7]),
    .Y(_001_));
 sg13g2_nor2_1 _606_ (.A(_039_),
    .B(_001_),
    .Y(output_o[112]));
 sg13g2_nand2_1 _607_ (.Y(output_no[112]),
    .A(_038_),
    .B(_000_));
 sg13g2_nor2_1 _608_ (.A(_041_),
    .B(_001_),
    .Y(output_o[113]));
 sg13g2_nand2_1 _609_ (.Y(output_no[113]),
    .A(_040_),
    .B(_000_));
 sg13g2_nor2_1 _610_ (.A(_043_),
    .B(_001_),
    .Y(output_o[114]));
 sg13g2_nand2_1 _611_ (.Y(output_no[114]),
    .A(_042_),
    .B(_000_));
 sg13g2_nor2_1 _612_ (.A(_045_),
    .B(_001_),
    .Y(output_o[115]));
 sg13g2_nand2_1 _613_ (.Y(output_no[115]),
    .A(_044_),
    .B(_000_));
 sg13g2_nor2_1 _614_ (.A(_047_),
    .B(_001_),
    .Y(output_o[116]));
 sg13g2_nand2_1 _615_ (.Y(output_no[116]),
    .A(_046_),
    .B(_000_));
 sg13g2_nor2_1 _616_ (.A(_049_),
    .B(_001_),
    .Y(output_o[117]));
 sg13g2_nand2_1 _617_ (.Y(output_no[117]),
    .A(_048_),
    .B(_000_));
 sg13g2_nor2_1 _618_ (.A(_051_),
    .B(_001_),
    .Y(output_o[118]));
 sg13g2_nand2_1 _619_ (.Y(output_no[118]),
    .A(_050_),
    .B(_000_));
 sg13g2_nor2_1 _620_ (.A(_053_),
    .B(_001_),
    .Y(output_o[119]));
 sg13g2_nand2_1 _621_ (.Y(output_no[119]),
    .A(_052_),
    .B(_000_));
 sg13g2_nor2_1 _622_ (.A(_055_),
    .B(_001_),
    .Y(output_o[120]));
 sg13g2_nand2_1 _623_ (.Y(output_no[120]),
    .A(_054_),
    .B(_000_));
 sg13g2_nor2_1 _624_ (.A(_057_),
    .B(_001_),
    .Y(output_o[121]));
 sg13g2_nand2_1 _625_ (.Y(output_no[121]),
    .A(_056_),
    .B(_000_));
 sg13g2_nor2_1 _626_ (.A(_059_),
    .B(_001_),
    .Y(output_o[122]));
 sg13g2_nand2_1 _627_ (.Y(output_no[122]),
    .A(_058_),
    .B(_000_));
 sg13g2_nor2_1 _628_ (.A(_061_),
    .B(_001_),
    .Y(output_o[123]));
 sg13g2_nand2_1 _629_ (.Y(output_no[123]),
    .A(_060_),
    .B(_000_));
 sg13g2_nor2_1 _630_ (.A(_063_),
    .B(_001_),
    .Y(output_o[124]));
 sg13g2_nand2_1 _631_ (.Y(output_no[124]),
    .A(_062_),
    .B(_000_));
 sg13g2_nor2_1 _632_ (.A(_065_),
    .B(_001_),
    .Y(output_o[125]));
 sg13g2_nand2_1 _633_ (.Y(output_no[125]),
    .A(_064_),
    .B(_000_));
 sg13g2_nor2_1 _634_ (.A(_067_),
    .B(_001_),
    .Y(output_o[126]));
 sg13g2_nand2_1 _635_ (.Y(output_no[126]),
    .A(_066_),
    .B(_000_));
 sg13g2_nor2_1 _636_ (.A(_069_),
    .B(_001_),
    .Y(output_o[127]));
 sg13g2_nand2_1 _637_ (.Y(output_no[127]),
    .A(_068_),
    .B(_000_));
 sg13g2_nor2_1 _638_ (.A(_010_),
    .B(_013_),
    .Y(output_o[128]));
 sg13g2_or2_1 _639_ (.X(output_no[128]),
    .B(_013_),
    .A(_010_));
 sg13g2_nor2_1 _640_ (.A(_010_),
    .B(_018_),
    .Y(output_o[129]));
 sg13g2_or2_1 _641_ (.X(output_no[129]),
    .B(_018_),
    .A(_010_));
 sg13g2_nor2_1 _642_ (.A(_010_),
    .B(_020_),
    .Y(output_o[130]));
 sg13g2_or2_1 _643_ (.X(output_no[130]),
    .B(_020_),
    .A(_010_));
 sg13g2_nor2_1 _644_ (.A(_010_),
    .B(_021_),
    .Y(output_o[131]));
 sg13g2_or2_1 _645_ (.X(output_no[131]),
    .B(_021_),
    .A(_010_));
 sg13g2_nor2_1 _646_ (.A(_010_),
    .B(_023_),
    .Y(output_o[132]));
 sg13g2_or2_1 _647_ (.X(output_no[132]),
    .B(_023_),
    .A(_010_));
 sg13g2_nor2_1 _648_ (.A(_010_),
    .B(_024_),
    .Y(output_o[133]));
 sg13g2_or2_1 _649_ (.X(output_no[133]),
    .B(_024_),
    .A(_010_));
 sg13g2_nor2_1 _650_ (.A(_010_),
    .B(_025_),
    .Y(output_o[134]));
 sg13g2_or2_1 _651_ (.X(output_no[134]),
    .B(_025_),
    .A(_010_));
 sg13g2_nor2_1 _652_ (.A(_010_),
    .B(_026_),
    .Y(output_o[135]));
 sg13g2_or2_1 _653_ (.X(output_no[135]),
    .B(_026_),
    .A(_010_));
 sg13g2_nor2_1 _654_ (.A(_010_),
    .B(_028_),
    .Y(output_o[136]));
 sg13g2_or2_1 _655_ (.X(output_no[136]),
    .B(_028_),
    .A(_010_));
 sg13g2_nor2_1 _656_ (.A(_010_),
    .B(_029_),
    .Y(output_o[137]));
 sg13g2_or2_1 _657_ (.X(output_no[137]),
    .B(_029_),
    .A(_010_));
 sg13g2_nor2_1 _658_ (.A(_010_),
    .B(_030_),
    .Y(output_o[138]));
 sg13g2_or2_1 _659_ (.X(output_no[138]),
    .B(_030_),
    .A(_010_));
 sg13g2_nor2_1 _660_ (.A(_010_),
    .B(_031_),
    .Y(output_o[139]));
 sg13g2_or2_1 _661_ (.X(output_no[139]),
    .B(_031_),
    .A(_010_));
 sg13g2_nor2_1 _662_ (.A(_010_),
    .B(_032_),
    .Y(output_o[140]));
 sg13g2_or2_1 _663_ (.X(output_no[140]),
    .B(_032_),
    .A(_010_));
 sg13g2_nor2_1 _664_ (.A(_010_),
    .B(_033_),
    .Y(output_o[141]));
 sg13g2_or2_1 _665_ (.X(output_no[141]),
    .B(_033_),
    .A(_010_));
 sg13g2_nor2_1 _666_ (.A(_010_),
    .B(_034_),
    .Y(output_o[142]));
 sg13g2_or2_1 _667_ (.X(output_no[142]),
    .B(_034_),
    .A(_010_));
 sg13g2_nor2_1 _668_ (.A(_004_),
    .B(_088_),
    .Y(_002_));
 sg13g2_or2_1 _669_ (.X(_003_),
    .B(_088_),
    .A(_004_));
 sg13g2_nor2_1 _670_ (.A(_039_),
    .B(_003_),
    .Y(output_o[0]));
 sg13g2_nand2_1 _671_ (.Y(output_no[0]),
    .A(_038_),
    .B(_002_));
 sg13g2_nor2_1 _672_ (.A(_041_),
    .B(_003_),
    .Y(output_o[1]));
 sg13g2_nand2_1 _673_ (.Y(output_no[1]),
    .A(_040_),
    .B(_002_));
 sg13g2_nor2_1 _674_ (.A(_043_),
    .B(_003_),
    .Y(output_o[2]));
 sg13g2_nand2_1 _675_ (.Y(output_no[2]),
    .A(_042_),
    .B(_002_));
 sg13g2_nor2_1 _676_ (.A(_045_),
    .B(_003_),
    .Y(output_o[3]));
 sg13g2_nand2_1 _677_ (.Y(output_no[3]),
    .A(_044_),
    .B(_002_));
 sg13g2_nor2_1 _678_ (.A(_047_),
    .B(_003_),
    .Y(output_o[4]));
 sg13g2_nand2_1 _679_ (.Y(output_no[4]),
    .A(_046_),
    .B(_002_));
 sg13g2_nor2_1 _680_ (.A(_049_),
    .B(_003_),
    .Y(output_o[5]));
 sg13g2_nand2_1 _681_ (.Y(output_no[5]),
    .A(_048_),
    .B(_002_));
 sg13g2_nor2_1 _682_ (.A(_051_),
    .B(_003_),
    .Y(output_o[6]));
 sg13g2_nand2_1 _683_ (.Y(output_no[6]),
    .A(_050_),
    .B(_002_));
 sg13g2_nor2_1 _684_ (.A(_053_),
    .B(_003_),
    .Y(output_o[7]));
 sg13g2_nand2_1 _685_ (.Y(output_no[7]),
    .A(_052_),
    .B(_002_));
 sg13g2_nor2_1 _686_ (.A(_055_),
    .B(_003_),
    .Y(output_o[8]));
 sg13g2_nand2_1 _687_ (.Y(output_no[8]),
    .A(_054_),
    .B(_002_));
 sg13g2_nor2_1 _688_ (.A(_057_),
    .B(_003_),
    .Y(output_o[9]));
 sg13g2_nand2_1 _689_ (.Y(output_no[9]),
    .A(_056_),
    .B(_002_));
 sg13g2_nor2_1 _690_ (.A(_059_),
    .B(_003_),
    .Y(output_o[10]));
 sg13g2_nand2_1 _691_ (.Y(output_no[10]),
    .A(_058_),
    .B(_002_));
 sg13g2_nor2_1 _692_ (.A(_061_),
    .B(_003_),
    .Y(output_o[11]));
 sg13g2_nand2_1 _693_ (.Y(output_no[11]),
    .A(_060_),
    .B(_002_));
 sg13g2_nor2_1 _694_ (.A(_063_),
    .B(_003_),
    .Y(output_o[12]));
 sg13g2_nand2_1 _695_ (.Y(output_no[12]),
    .A(_062_),
    .B(_002_));
 sg13g2_nor2_1 _696_ (.A(_065_),
    .B(_003_),
    .Y(output_o[13]));
 sg13g2_nand2_1 _697_ (.Y(output_no[13]),
    .A(_064_),
    .B(_002_));
 sg13g2_nor2_1 _698_ (.A(_067_),
    .B(_003_),
    .Y(output_o[14]));
 sg13g2_nand2_1 _699_ (.Y(output_no[14]),
    .A(_066_),
    .B(_002_));
 sg13g2_nor2_1 _700_ (.A(_069_),
    .B(_003_),
    .Y(output_o[15]));
 sg13g2_nand2_1 _701_ (.Y(output_no[15]),
    .A(_068_),
    .B(_002_));
 sg13g2_decap_4 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_256 ();
 sg13g2_fill_1 FILLER_0_258 ();
 sg13g2_fill_2 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_381 ();
 sg13g2_fill_1 FILLER_0_446 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_fill_2 FILLER_0_532 ();
 sg13g2_fill_1 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_4 FILLER_0_574 ();
 sg13g2_fill_1 FILLER_0_578 ();
 sg13g2_fill_1 FILLER_0_593 ();
 sg13g2_decap_4 FILLER_0_603 ();
 sg13g2_fill_2 FILLER_0_607 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_639 ();
 sg13g2_fill_2 FILLER_0_834 ();
 sg13g2_fill_1 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_13 ();
 sg13g2_decap_8 FILLER_1_20 ();
 sg13g2_decap_8 FILLER_1_27 ();
 sg13g2_decap_8 FILLER_1_34 ();
 sg13g2_decap_8 FILLER_1_41 ();
 sg13g2_fill_1 FILLER_1_48 ();
 sg13g2_decap_8 FILLER_1_53 ();
 sg13g2_decap_4 FILLER_1_60 ();
 sg13g2_decap_8 FILLER_1_68 ();
 sg13g2_decap_8 FILLER_1_75 ();
 sg13g2_decap_8 FILLER_1_82 ();
 sg13g2_decap_8 FILLER_1_89 ();
 sg13g2_decap_8 FILLER_1_96 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_8 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_decap_8 FILLER_1_124 ();
 sg13g2_decap_8 FILLER_1_131 ();
 sg13g2_decap_8 FILLER_1_138 ();
 sg13g2_decap_8 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_decap_8 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_fill_1 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_206 ();
 sg13g2_decap_8 FILLER_1_213 ();
 sg13g2_decap_8 FILLER_1_220 ();
 sg13g2_decap_8 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_241 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_288 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_fill_2 FILLER_1_323 ();
 sg13g2_fill_1 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_decap_8 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_4 FILLER_1_442 ();
 sg13g2_fill_2 FILLER_1_446 ();
 sg13g2_decap_8 FILLER_1_452 ();
 sg13g2_decap_8 FILLER_1_459 ();
 sg13g2_decap_8 FILLER_1_466 ();
 sg13g2_decap_8 FILLER_1_473 ();
 sg13g2_decap_8 FILLER_1_480 ();
 sg13g2_decap_8 FILLER_1_487 ();
 sg13g2_decap_8 FILLER_1_494 ();
 sg13g2_decap_8 FILLER_1_501 ();
 sg13g2_decap_8 FILLER_1_508 ();
 sg13g2_decap_8 FILLER_1_515 ();
 sg13g2_decap_4 FILLER_1_522 ();
 sg13g2_fill_1 FILLER_1_526 ();
 sg13g2_fill_2 FILLER_1_540 ();
 sg13g2_decap_8 FILLER_1_551 ();
 sg13g2_fill_1 FILLER_1_558 ();
 sg13g2_decap_8 FILLER_1_563 ();
 sg13g2_decap_8 FILLER_1_570 ();
 sg13g2_decap_8 FILLER_1_577 ();
 sg13g2_fill_2 FILLER_1_584 ();
 sg13g2_fill_1 FILLER_1_586 ();
 sg13g2_decap_4 FILLER_1_600 ();
 sg13g2_fill_1 FILLER_1_604 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_fill_2 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_622 ();
 sg13g2_decap_8 FILLER_1_629 ();
 sg13g2_decap_8 FILLER_1_636 ();
 sg13g2_fill_2 FILLER_1_643 ();
 sg13g2_decap_8 FILLER_1_649 ();
 sg13g2_decap_8 FILLER_1_656 ();
 sg13g2_decap_4 FILLER_1_663 ();
 sg13g2_fill_2 FILLER_1_667 ();
 sg13g2_decap_8 FILLER_1_673 ();
 sg13g2_decap_4 FILLER_1_680 ();
 sg13g2_fill_1 FILLER_1_684 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_fill_2 FILLER_1_696 ();
 sg13g2_decap_8 FILLER_1_702 ();
 sg13g2_decap_8 FILLER_1_709 ();
 sg13g2_decap_8 FILLER_1_716 ();
 sg13g2_decap_8 FILLER_1_723 ();
 sg13g2_decap_8 FILLER_1_730 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_decap_8 FILLER_1_751 ();
 sg13g2_decap_8 FILLER_1_758 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_decap_8 FILLER_1_772 ();
 sg13g2_decap_8 FILLER_1_779 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_4 FILLER_1_821 ();
 sg13g2_fill_1 FILLER_1_825 ();
 sg13g2_decap_4 FILLER_1_830 ();
 sg13g2_fill_1 FILLER_1_834 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_decap_8 FILLER_1_930 ();
 sg13g2_decap_8 FILLER_1_937 ();
 sg13g2_decap_8 FILLER_1_944 ();
 sg13g2_decap_4 FILLER_1_951 ();
 sg13g2_fill_2 FILLER_1_955 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_decap_8 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_989 ();
 sg13g2_decap_8 FILLER_1_996 ();
 sg13g2_decap_8 FILLER_1_1003 ();
 sg13g2_fill_2 FILLER_1_1010 ();
 sg13g2_fill_1 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1017 ();
 sg13g2_decap_4 FILLER_1_1024 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_9 ();
 sg13g2_fill_1 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_23 ();
 sg13g2_decap_8 FILLER_2_36 ();
 sg13g2_decap_8 FILLER_2_43 ();
 sg13g2_decap_8 FILLER_2_50 ();
 sg13g2_fill_1 FILLER_2_61 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_4 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_4 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_197 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_decap_8 FILLER_2_208 ();
 sg13g2_decap_4 FILLER_2_215 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_225 ();
 sg13g2_decap_4 FILLER_2_232 ();
 sg13g2_fill_1 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_241 ();
 sg13g2_decap_8 FILLER_2_248 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_decap_4 FILLER_2_262 ();
 sg13g2_fill_2 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_4 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_288 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_fill_1 FILLER_2_312 ();
 sg13g2_decap_4 FILLER_2_317 ();
 sg13g2_fill_2 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_fill_2 FILLER_2_383 ();
 sg13g2_fill_2 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_4 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_414 ();
 sg13g2_decap_4 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_425 ();
 sg13g2_decap_4 FILLER_2_435 ();
 sg13g2_decap_8 FILLER_2_443 ();
 sg13g2_fill_2 FILLER_2_450 ();
 sg13g2_decap_4 FILLER_2_456 ();
 sg13g2_decap_8 FILLER_2_464 ();
 sg13g2_decap_4 FILLER_2_471 ();
 sg13g2_fill_1 FILLER_2_475 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_4 FILLER_2_487 ();
 sg13g2_fill_1 FILLER_2_491 ();
 sg13g2_fill_1 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_509 ();
 sg13g2_decap_8 FILLER_2_516 ();
 sg13g2_decap_8 FILLER_2_523 ();
 sg13g2_decap_8 FILLER_2_530 ();
 sg13g2_decap_8 FILLER_2_537 ();
 sg13g2_decap_8 FILLER_2_544 ();
 sg13g2_decap_8 FILLER_2_551 ();
 sg13g2_decap_4 FILLER_2_558 ();
 sg13g2_fill_1 FILLER_2_562 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_fill_1 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_608 ();
 sg13g2_decap_8 FILLER_2_615 ();
 sg13g2_fill_1 FILLER_2_622 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_fill_1 FILLER_2_652 ();
 sg13g2_decap_8 FILLER_2_657 ();
 sg13g2_decap_8 FILLER_2_664 ();
 sg13g2_decap_8 FILLER_2_671 ();
 sg13g2_decap_8 FILLER_2_678 ();
 sg13g2_decap_8 FILLER_2_685 ();
 sg13g2_fill_2 FILLER_2_692 ();
 sg13g2_fill_1 FILLER_2_694 ();
 sg13g2_decap_8 FILLER_2_699 ();
 sg13g2_decap_8 FILLER_2_706 ();
 sg13g2_decap_8 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_720 ();
 sg13g2_decap_8 FILLER_2_727 ();
 sg13g2_decap_8 FILLER_2_734 ();
 sg13g2_decap_8 FILLER_2_741 ();
 sg13g2_decap_4 FILLER_2_748 ();
 sg13g2_fill_1 FILLER_2_752 ();
 sg13g2_fill_2 FILLER_2_769 ();
 sg13g2_fill_1 FILLER_2_771 ();
 sg13g2_decap_4 FILLER_2_776 ();
 sg13g2_fill_1 FILLER_2_780 ();
 sg13g2_decap_8 FILLER_2_785 ();
 sg13g2_decap_4 FILLER_2_792 ();
 sg13g2_decap_8 FILLER_2_800 ();
 sg13g2_decap_4 FILLER_2_807 ();
 sg13g2_fill_1 FILLER_2_811 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_848 ();
 sg13g2_decap_4 FILLER_2_855 ();
 sg13g2_fill_1 FILLER_2_859 ();
 sg13g2_decap_8 FILLER_2_864 ();
 sg13g2_decap_4 FILLER_2_871 ();
 sg13g2_fill_1 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_fill_2 FILLER_2_959 ();
 sg13g2_fill_2 FILLER_2_965 ();
 sg13g2_fill_1 FILLER_2_967 ();
 sg13g2_decap_8 FILLER_2_972 ();
 sg13g2_decap_4 FILLER_2_979 ();
 sg13g2_fill_1 FILLER_2_983 ();
 sg13g2_decap_8 FILLER_2_988 ();
 sg13g2_fill_2 FILLER_2_995 ();
 sg13g2_decap_8 FILLER_2_1017 ();
 sg13g2_decap_4 FILLER_2_1024 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_17 ();
 sg13g2_decap_8 FILLER_3_24 ();
 sg13g2_decap_4 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_57 ();
 sg13g2_fill_1 FILLER_3_64 ();
 sg13g2_decap_4 FILLER_3_77 ();
 sg13g2_decap_4 FILLER_3_125 ();
 sg13g2_fill_1 FILLER_3_141 ();
 sg13g2_decap_4 FILLER_3_195 ();
 sg13g2_fill_2 FILLER_3_199 ();
 sg13g2_decap_4 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_223 ();
 sg13g2_fill_2 FILLER_3_236 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_decap_4 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_2 FILLER_3_269 ();
 sg13g2_fill_1 FILLER_3_271 ();
 sg13g2_fill_1 FILLER_3_280 ();
 sg13g2_decap_4 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_301 ();
 sg13g2_decap_4 FILLER_3_314 ();
 sg13g2_fill_1 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_fill_1 FILLER_3_386 ();
 sg13g2_fill_2 FILLER_3_396 ();
 sg13g2_fill_2 FILLER_3_410 ();
 sg13g2_fill_1 FILLER_3_412 ();
 sg13g2_fill_1 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_3_443 ();
 sg13g2_decap_4 FILLER_3_450 ();
 sg13g2_fill_2 FILLER_3_454 ();
 sg13g2_decap_4 FILLER_3_460 ();
 sg13g2_decap_4 FILLER_3_476 ();
 sg13g2_fill_1 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_493 ();
 sg13g2_fill_2 FILLER_3_500 ();
 sg13g2_fill_1 FILLER_3_502 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_fill_1 FILLER_3_514 ();
 sg13g2_decap_8 FILLER_3_528 ();
 sg13g2_decap_4 FILLER_3_535 ();
 sg13g2_fill_2 FILLER_3_539 ();
 sg13g2_fill_2 FILLER_3_545 ();
 sg13g2_fill_1 FILLER_3_547 ();
 sg13g2_decap_8 FILLER_3_552 ();
 sg13g2_decap_4 FILLER_3_559 ();
 sg13g2_fill_2 FILLER_3_563 ();
 sg13g2_decap_8 FILLER_3_573 ();
 sg13g2_fill_1 FILLER_3_580 ();
 sg13g2_decap_8 FILLER_3_590 ();
 sg13g2_fill_2 FILLER_3_597 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_fill_1 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_639 ();
 sg13g2_decap_4 FILLER_3_646 ();
 sg13g2_fill_1 FILLER_3_650 ();
 sg13g2_fill_2 FILLER_3_655 ();
 sg13g2_fill_1 FILLER_3_657 ();
 sg13g2_fill_2 FILLER_3_670 ();
 sg13g2_fill_1 FILLER_3_672 ();
 sg13g2_decap_4 FILLER_3_685 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_4 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_4 FILLER_3_770 ();
 sg13g2_fill_2 FILLER_3_782 ();
 sg13g2_fill_1 FILLER_3_784 ();
 sg13g2_fill_2 FILLER_3_797 ();
 sg13g2_fill_1 FILLER_3_799 ();
 sg13g2_fill_1 FILLER_3_804 ();
 sg13g2_fill_2 FILLER_3_813 ();
 sg13g2_fill_1 FILLER_3_815 ();
 sg13g2_decap_4 FILLER_3_832 ();
 sg13g2_fill_2 FILLER_3_836 ();
 sg13g2_fill_2 FILLER_3_846 ();
 sg13g2_fill_1 FILLER_3_848 ();
 sg13g2_fill_2 FILLER_3_861 ();
 sg13g2_fill_1 FILLER_3_863 ();
 sg13g2_decap_8 FILLER_3_876 ();
 sg13g2_decap_8 FILLER_3_883 ();
 sg13g2_decap_8 FILLER_3_890 ();
 sg13g2_fill_1 FILLER_3_897 ();
 sg13g2_fill_2 FILLER_3_962 ();
 sg13g2_fill_1 FILLER_3_964 ();
 sg13g2_decap_4 FILLER_3_969 ();
 sg13g2_fill_2 FILLER_3_985 ();
 sg13g2_fill_1 FILLER_3_987 ();
 sg13g2_fill_1 FILLER_3_992 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_decap_8 FILLER_4_75 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_decap_8 FILLER_4_89 ();
 sg13g2_decap_8 FILLER_4_96 ();
 sg13g2_decap_8 FILLER_4_103 ();
 sg13g2_decap_8 FILLER_4_110 ();
 sg13g2_decap_8 FILLER_4_117 ();
 sg13g2_decap_8 FILLER_4_124 ();
 sg13g2_decap_8 FILLER_4_131 ();
 sg13g2_decap_8 FILLER_4_138 ();
 sg13g2_decap_8 FILLER_4_145 ();
 sg13g2_decap_8 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_159 ();
 sg13g2_decap_8 FILLER_4_166 ();
 sg13g2_decap_8 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_180 ();
 sg13g2_decap_8 FILLER_4_201 ();
 sg13g2_decap_8 FILLER_4_208 ();
 sg13g2_decap_8 FILLER_4_215 ();
 sg13g2_decap_8 FILLER_4_222 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_fill_2 FILLER_4_243 ();
 sg13g2_decap_4 FILLER_4_257 ();
 sg13g2_fill_2 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_4 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_4 FILLER_4_373 ();
 sg13g2_fill_2 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_4 FILLER_4_419 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_fill_2 FILLER_4_452 ();
 sg13g2_fill_1 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_472 ();
 sg13g2_decap_8 FILLER_4_478 ();
 sg13g2_decap_8 FILLER_4_485 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_fill_1 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_505 ();
 sg13g2_decap_4 FILLER_4_512 ();
 sg13g2_fill_2 FILLER_4_524 ();
 sg13g2_fill_1 FILLER_4_526 ();
 sg13g2_decap_4 FILLER_4_532 ();
 sg13g2_fill_1 FILLER_4_536 ();
 sg13g2_fill_2 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_556 ();
 sg13g2_decap_4 FILLER_4_563 ();
 sg13g2_decap_8 FILLER_4_572 ();
 sg13g2_decap_8 FILLER_4_579 ();
 sg13g2_decap_8 FILLER_4_586 ();
 sg13g2_decap_4 FILLER_4_593 ();
 sg13g2_fill_1 FILLER_4_597 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_fill_2 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_646 ();
 sg13g2_decap_8 FILLER_4_653 ();
 sg13g2_decap_8 FILLER_4_660 ();
 sg13g2_decap_8 FILLER_4_667 ();
 sg13g2_decap_8 FILLER_4_674 ();
 sg13g2_fill_2 FILLER_4_681 ();
 sg13g2_fill_1 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_4 FILLER_4_700 ();
 sg13g2_fill_2 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_715 ();
 sg13g2_decap_8 FILLER_4_722 ();
 sg13g2_decap_8 FILLER_4_729 ();
 sg13g2_decap_8 FILLER_4_736 ();
 sg13g2_decap_8 FILLER_4_743 ();
 sg13g2_decap_8 FILLER_4_750 ();
 sg13g2_decap_8 FILLER_4_757 ();
 sg13g2_fill_1 FILLER_4_764 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_4 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_904 ();
 sg13g2_decap_8 FILLER_4_911 ();
 sg13g2_decap_8 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_925 ();
 sg13g2_decap_8 FILLER_4_932 ();
 sg13g2_decap_8 FILLER_4_939 ();
 sg13g2_fill_1 FILLER_4_946 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1026 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_8 FILLER_5_404 ();
 sg13g2_decap_8 FILLER_5_411 ();
 sg13g2_decap_4 FILLER_5_418 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_decap_8 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_457 ();
 sg13g2_decap_4 FILLER_5_464 ();
 sg13g2_fill_1 FILLER_5_468 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_fill_2 FILLER_5_490 ();
 sg13g2_fill_1 FILLER_5_506 ();
 sg13g2_decap_4 FILLER_5_512 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_4 FILLER_5_532 ();
 sg13g2_fill_1 FILLER_5_536 ();
 sg13g2_decap_4 FILLER_5_546 ();
 sg13g2_fill_1 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_555 ();
 sg13g2_fill_1 FILLER_5_562 ();
 sg13g2_decap_4 FILLER_5_572 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_fill_2 FILLER_5_592 ();
 sg13g2_fill_1 FILLER_5_594 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_4 FILLER_5_616 ();
 sg13g2_fill_2 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_4 FILLER_5_751 ();
 sg13g2_fill_2 FILLER_5_755 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_decap_8 FILLER_5_778 ();
 sg13g2_decap_8 FILLER_5_785 ();
 sg13g2_decap_8 FILLER_5_792 ();
 sg13g2_decap_8 FILLER_5_799 ();
 sg13g2_decap_8 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_813 ();
 sg13g2_decap_8 FILLER_5_820 ();
 sg13g2_decap_8 FILLER_5_827 ();
 sg13g2_decap_8 FILLER_5_834 ();
 sg13g2_decap_8 FILLER_5_841 ();
 sg13g2_fill_1 FILLER_5_848 ();
 sg13g2_decap_8 FILLER_5_853 ();
 sg13g2_decap_8 FILLER_5_860 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_881 ();
 sg13g2_decap_8 FILLER_5_888 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_916 ();
 sg13g2_decap_8 FILLER_5_923 ();
 sg13g2_decap_8 FILLER_5_930 ();
 sg13g2_decap_8 FILLER_5_937 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_fill_1 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_433 ();
 sg13g2_decap_8 FILLER_6_440 ();
 sg13g2_decap_4 FILLER_6_447 ();
 sg13g2_fill_1 FILLER_6_451 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_478 ();
 sg13g2_decap_8 FILLER_6_485 ();
 sg13g2_decap_8 FILLER_6_492 ();
 sg13g2_decap_8 FILLER_6_499 ();
 sg13g2_decap_8 FILLER_6_506 ();
 sg13g2_decap_4 FILLER_6_513 ();
 sg13g2_fill_2 FILLER_6_517 ();
 sg13g2_decap_8 FILLER_6_523 ();
 sg13g2_decap_4 FILLER_6_530 ();
 sg13g2_decap_4 FILLER_6_545 ();
 sg13g2_fill_1 FILLER_6_549 ();
 sg13g2_fill_2 FILLER_6_557 ();
 sg13g2_decap_4 FILLER_6_563 ();
 sg13g2_fill_2 FILLER_6_567 ();
 sg13g2_fill_2 FILLER_6_576 ();
 sg13g2_decap_8 FILLER_6_587 ();
 sg13g2_decap_4 FILLER_6_594 ();
 sg13g2_fill_1 FILLER_6_598 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_decap_8 FILLER_6_610 ();
 sg13g2_decap_8 FILLER_6_617 ();
 sg13g2_decap_4 FILLER_6_624 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_8 FILLER_6_663 ();
 sg13g2_decap_8 FILLER_6_670 ();
 sg13g2_decap_8 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_698 ();
 sg13g2_decap_8 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_8 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_866 ();
 sg13g2_decap_8 FILLER_6_873 ();
 sg13g2_decap_8 FILLER_6_880 ();
 sg13g2_decap_8 FILLER_6_887 ();
 sg13g2_decap_8 FILLER_6_894 ();
 sg13g2_decap_8 FILLER_6_901 ();
 sg13g2_decap_8 FILLER_6_908 ();
 sg13g2_decap_8 FILLER_6_915 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_943 ();
 sg13g2_decap_8 FILLER_6_950 ();
 sg13g2_decap_8 FILLER_6_957 ();
 sg13g2_decap_8 FILLER_6_964 ();
 sg13g2_decap_8 FILLER_6_971 ();
 sg13g2_decap_8 FILLER_6_978 ();
 sg13g2_decap_8 FILLER_6_985 ();
 sg13g2_decap_8 FILLER_6_992 ();
 sg13g2_decap_8 FILLER_6_999 ();
 sg13g2_decap_8 FILLER_6_1006 ();
 sg13g2_decap_8 FILLER_6_1013 ();
 sg13g2_decap_8 FILLER_6_1020 ();
 sg13g2_fill_2 FILLER_6_1027 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_1 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_433 ();
 sg13g2_decap_8 FILLER_7_440 ();
 sg13g2_decap_8 FILLER_7_447 ();
 sg13g2_fill_2 FILLER_7_454 ();
 sg13g2_fill_1 FILLER_7_456 ();
 sg13g2_decap_8 FILLER_7_461 ();
 sg13g2_fill_2 FILLER_7_468 ();
 sg13g2_fill_2 FILLER_7_475 ();
 sg13g2_decap_4 FILLER_7_483 ();
 sg13g2_fill_2 FILLER_7_487 ();
 sg13g2_fill_2 FILLER_7_494 ();
 sg13g2_decap_8 FILLER_7_510 ();
 sg13g2_decap_8 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_524 ();
 sg13g2_decap_8 FILLER_7_531 ();
 sg13g2_decap_8 FILLER_7_538 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_decap_8 FILLER_7_559 ();
 sg13g2_decap_8 FILLER_7_566 ();
 sg13g2_decap_8 FILLER_7_573 ();
 sg13g2_decap_8 FILLER_7_580 ();
 sg13g2_decap_8 FILLER_7_587 ();
 sg13g2_decap_8 FILLER_7_594 ();
 sg13g2_decap_8 FILLER_7_601 ();
 sg13g2_decap_8 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_615 ();
 sg13g2_decap_8 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_629 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_decap_8 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_650 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_decap_8 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_671 ();
 sg13g2_decap_8 FILLER_7_678 ();
 sg13g2_decap_8 FILLER_7_685 ();
 sg13g2_decap_8 FILLER_7_692 ();
 sg13g2_decap_8 FILLER_7_699 ();
 sg13g2_decap_8 FILLER_7_706 ();
 sg13g2_decap_8 FILLER_7_713 ();
 sg13g2_decap_8 FILLER_7_720 ();
 sg13g2_decap_8 FILLER_7_727 ();
 sg13g2_decap_8 FILLER_7_734 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_8 FILLER_7_748 ();
 sg13g2_decap_8 FILLER_7_755 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_783 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_decap_8 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_846 ();
 sg13g2_decap_8 FILLER_7_853 ();
 sg13g2_decap_8 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_7_867 ();
 sg13g2_decap_8 FILLER_7_874 ();
 sg13g2_decap_8 FILLER_7_881 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_decap_8 FILLER_7_895 ();
 sg13g2_decap_8 FILLER_7_902 ();
 sg13g2_decap_8 FILLER_7_909 ();
 sg13g2_decap_8 FILLER_7_916 ();
 sg13g2_decap_8 FILLER_7_923 ();
 sg13g2_decap_8 FILLER_7_930 ();
 sg13g2_decap_8 FILLER_7_937 ();
 sg13g2_decap_8 FILLER_7_944 ();
 sg13g2_decap_8 FILLER_7_951 ();
 sg13g2_decap_8 FILLER_7_958 ();
 sg13g2_decap_8 FILLER_7_965 ();
 sg13g2_decap_8 FILLER_7_972 ();
 sg13g2_decap_8 FILLER_7_979 ();
 sg13g2_decap_8 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_993 ();
 sg13g2_decap_8 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_decap_8 FILLER_7_1014 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_decap_8 FILLER_10_875 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_decap_8 FILLER_10_903 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_decap_8 FILLER_10_938 ();
 sg13g2_decap_8 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_8 FILLER_10_1008 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_decap_8 FILLER_10_1022 ();
endmodule
