module decoder (ena_i,
    VPWR,
    VGND,
    input_ni,
    output_no,
    output_o);
 input ena_i;
 inout VPWR;
 inout VGND;
 input [7:0] input_ni;
 output [255:0] output_no;
 output [255:0] output_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;

 sg13g2_inv_1 _095_ (.VDD(VPWR),
    .Y(_004_),
    .A(net123),
    .VSS(VGND));
 sg13g2_nor2_1 _096_ (.A(net158),
    .B(net157),
    .Y(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _097_ (.A(net156),
    .B(net155),
    .Y(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _098_ (.A(net156),
    .B(net155),
    .C(net158),
    .Y(_007_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net157));
 sg13g2_nor2b_2 _099_ (.A(net122),
    .B_N(net161),
    .Y(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _100_ (.A(net159),
    .B(net160),
    .C(net128),
    .D(_008_),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _101_ (.B(net160),
    .C(net128),
    .A(net159),
    .Y(_010_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_008_));
 sg13g2_and2_1 _102_ (.A(_007_),
    .B(_009_),
    .X(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _103_ (.Y(net210),
    .A(_007_),
    .B(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _104_ (.A(net158),
    .B(net157),
    .X(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _105_ (.A(net156),
    .B(net155),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _106_ (.Y(_013_),
    .A(net117),
    .B(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _107_ (.A(net159),
    .B_N(net160),
    .Y(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _108_ (.X(_015_),
    .A(net128),
    .B(_008_),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _109_ (.B(_008_),
    .C(_014_),
    .A(net128),
    .Y(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _110_ (.A(_013_),
    .B(net97),
    .Y(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _111_ (.Y(net211),
    .B(_015_),
    .A_N(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _112_ (.A(net155),
    .B_N(net156),
    .Y(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _113_ (.Y(_018_),
    .A(net117),
    .B(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _114_ (.A(net97),
    .B(_018_),
    .Y(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _115_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net212),
    .B(_018_),
    .A(net97));
 sg13g2_nor2b_2 _116_ (.A(net156),
    .B_N(net155),
    .Y(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _117_ (.Y(_020_),
    .A(net117),
    .B(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _118_ (.A(net97),
    .B(_020_),
    .Y(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _119_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net213),
    .B(_020_),
    .A(net97));
 sg13g2_nand2_1 _120_ (.Y(_021_),
    .A(net118),
    .B(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _121_ (.A(net97),
    .B(_021_),
    .Y(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _122_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net214),
    .B(_021_),
    .A(net97));
 sg13g2_nor2b_1 _123_ (.A(net157),
    .B_N(net158),
    .Y(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _124_ (.Y(_023_),
    .A(net114),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _125_ (.A(net97),
    .B(_023_),
    .Y(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _126_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net215),
    .B(_023_),
    .A(net98));
 sg13g2_nand2_1 _127_ (.Y(_024_),
    .A(net112),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _128_ (.A(net98),
    .B(_024_),
    .Y(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _129_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net216),
    .B(_024_),
    .A(net98));
 sg13g2_nand2_1 _130_ (.Y(_025_),
    .A(net110),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _131_ (.A(net98),
    .B(_025_),
    .Y(net474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _132_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net218),
    .B(_025_),
    .A(net98));
 sg13g2_nand2_1 _133_ (.Y(_026_),
    .A(net118),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _134_ (.A(net98),
    .B(_026_),
    .Y(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _135_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net219),
    .B(_026_),
    .A(net98));
 sg13g2_nor2b_1 _136_ (.A(net158),
    .B_N(net157),
    .Y(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _137_ (.Y(_028_),
    .A(net114),
    .B(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _138_ (.A(net99),
    .B(_028_),
    .Y(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _139_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net220),
    .B(_028_),
    .A(net99));
 sg13g2_nand2_1 _140_ (.Y(_029_),
    .A(net112),
    .B(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _141_ (.A(net99),
    .B(_029_),
    .Y(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _142_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net221),
    .B(_029_),
    .A(net99));
 sg13g2_nand2_1 _143_ (.Y(_030_),
    .A(net110),
    .B(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _144_ (.A(net99),
    .B(_030_),
    .Y(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _145_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net222),
    .B(_030_),
    .A(net99));
 sg13g2_nand2_1 _146_ (.Y(_031_),
    .A(net118),
    .B(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _147_ (.A(net99),
    .B(_031_),
    .Y(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _148_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net223),
    .B(_031_),
    .A(net99));
 sg13g2_nand2_1 _149_ (.Y(_032_),
    .A(net119),
    .B(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _150_ (.A(net100),
    .B(_032_),
    .Y(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _151_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net224),
    .B(_032_),
    .A(net100));
 sg13g2_nand2_1 _152_ (.Y(_033_),
    .A(net119),
    .B(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _153_ (.A(net100),
    .B(_033_),
    .Y(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _154_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net225),
    .B(_033_),
    .A(net100));
 sg13g2_nand2_1 _155_ (.Y(_034_),
    .A(net119),
    .B(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _156_ (.A(net100),
    .B(_034_),
    .Y(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _157_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net226),
    .B(_034_),
    .A(net100));
 sg13g2_and2_1 _158_ (.A(_007_),
    .B(_015_),
    .X(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _159_ (.Y(net227),
    .A(_007_),
    .B(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _160_ (.A(net160),
    .B_N(net159),
    .Y(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _161_ (.A(_008_),
    .B(_035_),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _162_ (.Y(_037_),
    .A(_008_),
    .B(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _163_ (.X(_038_),
    .A(net124),
    .B(net116),
    .C(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _164_ (.B(net116),
    .C(net114),
    .A(net124),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _165_ (.A(net150),
    .B(net149),
    .Y(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _166_ (.Y(net229),
    .A(net95),
    .B(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _167_ (.X(_040_),
    .A(net124),
    .B(net116),
    .C(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _168_ (.B(net116),
    .C(net112),
    .A(net124),
    .Y(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _169_ (.A(net150),
    .B(net147),
    .Y(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _170_ (.Y(net230),
    .A(net95),
    .B(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _171_ (.X(_042_),
    .A(net124),
    .B(net116),
    .C(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _172_ (.B(net116),
    .C(net110),
    .A(net124),
    .Y(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _173_ (.A(net150),
    .B(net145),
    .Y(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _174_ (.Y(net231),
    .A(net95),
    .B(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _175_ (.X(_044_),
    .A(net124),
    .B(net118),
    .C(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _176_ (.B(net118),
    .C(net116),
    .A(net124),
    .Y(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _177_ (.A(net150),
    .B(net143),
    .Y(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _178_ (.Y(net232),
    .A(net95),
    .B(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _179_ (.X(_046_),
    .A(net125),
    .B(net114),
    .C(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _180_ (.B(net114),
    .C(net108),
    .A(net125),
    .Y(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _181_ (.A(net150),
    .B(net84),
    .Y(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _182_ (.Y(net233),
    .A(net95),
    .B(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _183_ (.X(_048_),
    .A(net125),
    .B(net112),
    .C(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _184_ (.B(net112),
    .C(net108),
    .A(net125),
    .Y(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _185_ (.A(net150),
    .B(net141),
    .Y(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _186_ (.Y(net234),
    .A(net95),
    .B(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _187_ (.X(_050_),
    .A(net125),
    .B(net110),
    .C(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _188_ (.B(net110),
    .C(net108),
    .A(net125),
    .Y(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _189_ (.A(net150),
    .B(net139),
    .Y(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _190_ (.Y(net235),
    .A(net95),
    .B(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _191_ (.X(_052_),
    .A(net126),
    .B(net118),
    .C(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _192_ (.B(net118),
    .C(net108),
    .A(net125),
    .Y(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _193_ (.A(net150),
    .B(net137),
    .Y(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _194_ (.Y(net236),
    .A(net95),
    .B(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _195_ (.X(_054_),
    .A(net126),
    .B(net115),
    .C(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _196_ (.B(net115),
    .C(net106),
    .A(net126),
    .Y(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _197_ (.A(net151),
    .B(net74),
    .Y(net493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _198_ (.Y(net237),
    .A(net96),
    .B(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _199_ (.X(_056_),
    .A(net126),
    .B(net113),
    .C(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _200_ (.B(net113),
    .C(net107),
    .A(net127),
    .Y(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _201_ (.A(net151),
    .B(net70),
    .Y(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _202_ (.Y(net238),
    .A(net96),
    .B(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _203_ (.X(_058_),
    .A(net126),
    .B(net111),
    .C(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _204_ (.B(net111),
    .C(net107),
    .A(net127),
    .Y(_059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _205_ (.A(net151),
    .B(net66),
    .Y(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _206_ (.Y(net240),
    .A(net96),
    .B(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _207_ (.X(_060_),
    .A(net126),
    .B(net118),
    .C(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _208_ (.B(_006_),
    .C(net106),
    .A(net129),
    .Y(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _209_ (.A(net151),
    .B(net62),
    .Y(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _210_ (.Y(net241),
    .A(net96),
    .B(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _211_ (.X(_062_),
    .A(net127),
    .B(net119),
    .C(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _212_ (.B(net119),
    .C(net115),
    .A(net127),
    .Y(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _213_ (.A(net151),
    .B(net58),
    .Y(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _214_ (.Y(net242),
    .A(net96),
    .B(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _215_ (.X(_064_),
    .A(net127),
    .B(net119),
    .C(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _216_ (.B(net119),
    .C(net113),
    .A(net127),
    .Y(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _217_ (.A(net151),
    .B(net54),
    .Y(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _218_ (.Y(net243),
    .A(net96),
    .B(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _219_ (.X(_066_),
    .A(net127),
    .B(net119),
    .C(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _220_ (.B(_005_),
    .C(net111),
    .A(net127),
    .Y(_067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _221_ (.A(net151),
    .B(net50),
    .Y(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _222_ (.Y(net244),
    .A(net96),
    .B(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _223_ (.A(net128),
    .B(_007_),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _224_ (.Y(_069_),
    .A(net128),
    .B(_007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _225_ (.A(net151),
    .B(net133),
    .Y(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _226_ (.Y(net245),
    .A(net96),
    .B(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _227_ (.A(net159),
    .B(net160),
    .Y(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _228_ (.A(_008_),
    .B(_070_),
    .X(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _229_ (.Y(_072_),
    .A(_008_),
    .B(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _230_ (.A(net149),
    .B(net45),
    .Y(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _231_ (.Y(net246),
    .A(net94),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _232_ (.A(net147),
    .B(net45),
    .Y(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _233_ (.Y(net247),
    .A(net92),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _234_ (.A(net145),
    .B(net45),
    .Y(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _235_ (.Y(net248),
    .A(net90),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _236_ (.A(net143),
    .B(net45),
    .Y(net505),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _237_ (.Y(net249),
    .A(net88),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _238_ (.A(net84),
    .B(net45),
    .Y(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _239_ (.Y(net251),
    .A(net86),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _240_ (.A(net141),
    .B(net45),
    .Y(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _241_ (.Y(net252),
    .A(net82),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _242_ (.A(net139),
    .B(net45),
    .Y(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _243_ (.Y(net253),
    .A(net80),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _244_ (.A(net137),
    .B(net45),
    .Y(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _245_ (.Y(net254),
    .A(net78),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _246_ (.A(net74),
    .B(net46),
    .Y(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _247_ (.Y(net255),
    .A(net76),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _248_ (.A(net70),
    .B(net46),
    .Y(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _249_ (.Y(net256),
    .A(net72),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _250_ (.A(net66),
    .B(net46),
    .Y(net513),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _251_ (.Y(net257),
    .A(net68),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _252_ (.A(net62),
    .B(net46),
    .Y(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _253_ (.Y(net258),
    .A(net64),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _254_ (.A(net58),
    .B(net46),
    .Y(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _255_ (.Y(net259),
    .A(net60),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _256_ (.A(net54),
    .B(net46),
    .Y(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _257_ (.Y(net260),
    .A(net56),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _258_ (.A(net50),
    .B(net46),
    .Y(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _259_ (.Y(net262),
    .A(net52),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _260_ (.A(net133),
    .B(net46),
    .Y(net519),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _261_ (.Y(net263),
    .A(net135),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _262_ (.A(net122),
    .B(net161),
    .Y(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _263_ (.X(_074_),
    .A(net159),
    .B(net160),
    .C(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _264_ (.B(net160),
    .C(_073_),
    .A(net159),
    .Y(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _265_ (.A(net149),
    .B(net41),
    .Y(net520),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _266_ (.Y(net264),
    .A(net94),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _267_ (.A(net147),
    .B(net41),
    .Y(net521),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _268_ (.Y(net265),
    .A(net92),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _269_ (.A(net145),
    .B(net41),
    .Y(net522),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _270_ (.Y(net266),
    .A(net90),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _271_ (.A(net143),
    .B(net41),
    .Y(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _272_ (.Y(net267),
    .A(net88),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _273_ (.A(net84),
    .B(net41),
    .Y(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _274_ (.Y(net268),
    .A(net86),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _275_ (.A(net141),
    .B(net41),
    .Y(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _276_ (.Y(net269),
    .A(net82),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _277_ (.A(net139),
    .B(net41),
    .Y(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _278_ (.Y(net270),
    .A(net80),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _279_ (.A(net137),
    .B(net41),
    .Y(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _280_ (.Y(net271),
    .A(net78),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _281_ (.A(net74),
    .B(net42),
    .Y(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _282_ (.Y(net274),
    .A(net76),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _283_ (.A(net70),
    .B(net42),
    .Y(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _284_ (.Y(net275),
    .A(net72),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _285_ (.A(net66),
    .B(net42),
    .Y(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _286_ (.Y(net276),
    .A(net68),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _287_ (.A(net62),
    .B(net42),
    .Y(net533),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _288_ (.Y(net277),
    .A(net64),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _289_ (.A(net58),
    .B(net42),
    .Y(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _290_ (.Y(net278),
    .A(net60),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _291_ (.A(net54),
    .B(net42),
    .Y(net535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _292_ (.Y(net279),
    .A(net56),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _293_ (.A(net50),
    .B(net42),
    .Y(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _294_ (.Y(net280),
    .A(net52),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _295_ (.A(net133),
    .B(net42),
    .Y(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _296_ (.Y(net281),
    .A(net135),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _297_ (.A(_014_),
    .B(_073_),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _298_ (.Y(_077_),
    .A(_014_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _299_ (.A(net149),
    .B(net37),
    .Y(net538),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _300_ (.Y(net282),
    .A(net94),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _301_ (.A(net147),
    .B(net37),
    .Y(net539),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _302_ (.Y(net283),
    .A(net92),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _303_ (.A(net145),
    .B(net37),
    .Y(net541),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _304_ (.Y(net285),
    .A(net90),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _305_ (.A(net143),
    .B(net37),
    .Y(net542),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _306_ (.Y(net286),
    .A(net88),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _307_ (.A(net84),
    .B(net37),
    .Y(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _308_ (.Y(net287),
    .A(net86),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _309_ (.A(net141),
    .B(net37),
    .Y(net544),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _310_ (.Y(net288),
    .A(net82),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _311_ (.A(net139),
    .B(net37),
    .Y(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _312_ (.Y(net289),
    .A(net80),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _313_ (.A(net137),
    .B(net37),
    .Y(net546),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _314_ (.Y(net290),
    .A(net78),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _315_ (.A(net74),
    .B(net38),
    .Y(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _316_ (.Y(net291),
    .A(net76),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _317_ (.A(net70),
    .B(net38),
    .Y(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _318_ (.Y(net292),
    .A(net72),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _319_ (.A(net66),
    .B(net38),
    .Y(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _320_ (.Y(net293),
    .A(net68),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _321_ (.A(net62),
    .B(net38),
    .Y(net550),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _322_ (.Y(net294),
    .A(net64),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _323_ (.A(net58),
    .B(net38),
    .Y(net552),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _324_ (.Y(net296),
    .A(net60),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _325_ (.A(net54),
    .B(net38),
    .Y(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _326_ (.Y(net297),
    .A(net56),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _327_ (.A(net50),
    .B(net38),
    .Y(net554),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _328_ (.Y(net298),
    .A(net52),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _329_ (.A(net133),
    .B(net38),
    .Y(net555),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _330_ (.Y(net299),
    .A(net135),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _331_ (.A(_035_),
    .B(_073_),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _332_ (.Y(_079_),
    .A(_035_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _333_ (.A(net149),
    .B(net33),
    .Y(net556),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _334_ (.Y(net300),
    .A(net94),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _335_ (.A(net147),
    .B(net33),
    .Y(net557),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _336_ (.Y(net301),
    .A(net92),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _337_ (.A(net145),
    .B(net33),
    .Y(net558),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _338_ (.Y(net302),
    .A(net90),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _339_ (.A(net143),
    .B(net33),
    .Y(net559),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _340_ (.Y(net303),
    .A(net88),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _341_ (.A(net84),
    .B(net33),
    .Y(net560),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _342_ (.Y(net304),
    .A(net86),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _343_ (.A(net141),
    .B(net33),
    .Y(net561),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _344_ (.Y(net305),
    .A(net82),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _345_ (.A(net139),
    .B(net33),
    .Y(net563),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _346_ (.Y(net307),
    .A(net80),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _347_ (.A(net137),
    .B(net33),
    .Y(net564),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _348_ (.Y(net308),
    .A(net78),
    .B(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _349_ (.A(net74),
    .B(net34),
    .Y(net565),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _350_ (.Y(net309),
    .A(net76),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _351_ (.A(net70),
    .B(net34),
    .Y(net566),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _352_ (.Y(net310),
    .A(net72),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _353_ (.A(net66),
    .B(net34),
    .Y(net567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _354_ (.Y(net311),
    .A(net68),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _355_ (.A(net62),
    .B(net34),
    .Y(net568),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _356_ (.Y(net312),
    .A(net64),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _357_ (.A(net58),
    .B(net34),
    .Y(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _358_ (.Y(net313),
    .A(net60),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _359_ (.A(net54),
    .B(net34),
    .Y(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _360_ (.Y(net314),
    .A(net56),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _361_ (.A(net50),
    .B(net34),
    .Y(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _362_ (.Y(net315),
    .A(net52),
    .B(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _363_ (.A(net133),
    .B(net34),
    .Y(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _364_ (.Y(net316),
    .A(net135),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _365_ (.A(_070_),
    .B(_073_),
    .X(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _366_ (.Y(_081_),
    .A(_070_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _367_ (.A(net149),
    .B(net154),
    .Y(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _368_ (.Y(net318),
    .A(net94),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _369_ (.A(net147),
    .B(net154),
    .Y(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _370_ (.Y(net319),
    .A(net92),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _371_ (.A(net145),
    .B(net154),
    .Y(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _372_ (.Y(net320),
    .A(net90),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _373_ (.A(net143),
    .B(net154),
    .Y(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _374_ (.Y(net321),
    .A(net88),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _375_ (.A(net84),
    .B(net153),
    .Y(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _376_ (.Y(net322),
    .A(net86),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _377_ (.A(net141),
    .B(net154),
    .Y(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _378_ (.Y(net323),
    .A(net82),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _379_ (.A(net139),
    .B(net154),
    .Y(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _380_ (.Y(net324),
    .A(net80),
    .B(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _381_ (.A(net137),
    .B(net154),
    .Y(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _382_ (.Y(net325),
    .A(net78),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _383_ (.A(net74),
    .B(net153),
    .Y(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _384_ (.Y(net326),
    .A(net76),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _385_ (.A(net70),
    .B(net153),
    .Y(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _386_ (.Y(net327),
    .A(net72),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _387_ (.A(net66),
    .B(net153),
    .Y(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _388_ (.Y(net329),
    .A(net68),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _389_ (.A(net62),
    .B(net153),
    .Y(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _390_ (.Y(net330),
    .A(net64),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _391_ (.A(net58),
    .B(net153),
    .Y(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _392_ (.Y(net331),
    .A(net60),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _393_ (.A(net54),
    .B(net153),
    .Y(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _394_ (.Y(net332),
    .A(net56),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _395_ (.A(net50),
    .B(net153),
    .Y(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _396_ (.Y(net333),
    .A(net52),
    .B(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _397_ (.A(net133),
    .B(_081_),
    .Y(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _398_ (.Y(net334),
    .A(net135),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _399_ (.X(_082_),
    .A(net120),
    .B(net123),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _400_ (.B(net123),
    .C(_014_),
    .A(net120),
    .Y(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _401_ (.A(net148),
    .B(net27),
    .Y(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _402_ (.Y(net239),
    .A(net93),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _403_ (.A(net146),
    .B(net27),
    .Y(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _404_ (.Y(net250),
    .A(net91),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _405_ (.A(net144),
    .B(net27),
    .Y(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _406_ (.Y(net261),
    .A(net89),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _407_ (.A(net142),
    .B(net27),
    .Y(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _408_ (.Y(net272),
    .A(net87),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _409_ (.A(net83),
    .B(net27),
    .Y(net540),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _410_ (.Y(net284),
    .A(net85),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _411_ (.A(net140),
    .B(net27),
    .Y(net551),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _412_ (.Y(net295),
    .A(net81),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _413_ (.A(net138),
    .B(net27),
    .Y(net562),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _414_ (.Y(net306),
    .A(net79),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _415_ (.A(net136),
    .B(net27),
    .Y(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _416_ (.Y(net317),
    .A(net77),
    .B(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _417_ (.A(net73),
    .B(net28),
    .Y(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _418_ (.Y(net328),
    .A(net75),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _419_ (.A(net69),
    .B(net28),
    .Y(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _420_ (.Y(net335),
    .A(net71),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _421_ (.A(net65),
    .B(net28),
    .Y(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _422_ (.Y(net336),
    .A(net67),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _423_ (.A(net61),
    .B(net28),
    .Y(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _424_ (.Y(net337),
    .A(net63),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _425_ (.A(net57),
    .B(net28),
    .Y(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _426_ (.Y(net338),
    .A(net59),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _427_ (.A(net53),
    .B(net28),
    .Y(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _428_ (.Y(net339),
    .A(net55),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _429_ (.A(net49),
    .B(net28),
    .Y(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _430_ (.Y(net341),
    .A(net51),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _431_ (.A(net132),
    .B(net28),
    .Y(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _432_ (.Y(net342),
    .A(net134),
    .B(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _433_ (.X(_084_),
    .A(net120),
    .B(net123),
    .C(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _434_ (.B(net123),
    .C(_035_),
    .A(net120),
    .Y(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _435_ (.A(net148),
    .B(net23),
    .Y(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _436_ (.Y(net343),
    .A(net93),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _437_ (.A(net146),
    .B(net23),
    .Y(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _438_ (.Y(net344),
    .A(net91),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _439_ (.A(net144),
    .B(net23),
    .Y(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _440_ (.Y(net345),
    .A(net89),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _441_ (.A(net142),
    .B(net23),
    .Y(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _442_ (.Y(net346),
    .A(net87),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _443_ (.A(net83),
    .B(net23),
    .Y(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _444_ (.Y(net347),
    .A(net85),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _445_ (.A(net140),
    .B(net23),
    .Y(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _446_ (.Y(net348),
    .A(net81),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _447_ (.A(net138),
    .B(net23),
    .Y(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _448_ (.Y(net349),
    .A(net79),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _449_ (.A(net136),
    .B(net23),
    .Y(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _450_ (.Y(net350),
    .A(net77),
    .B(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _451_ (.A(net73),
    .B(net24),
    .Y(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _452_ (.Y(net352),
    .A(net75),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _453_ (.A(net69),
    .B(net24),
    .Y(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _454_ (.Y(net353),
    .A(net71),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _455_ (.A(net65),
    .B(net24),
    .Y(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _456_ (.Y(net354),
    .A(net67),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _457_ (.A(net61),
    .B(net24),
    .Y(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _458_ (.Y(net355),
    .A(net63),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _459_ (.A(net57),
    .B(net24),
    .Y(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _460_ (.Y(net356),
    .A(net59),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _461_ (.A(net53),
    .B(net24),
    .Y(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _462_ (.Y(net357),
    .A(net55),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _463_ (.A(net49),
    .B(net24),
    .Y(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _464_ (.Y(net358),
    .A(net51),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _465_ (.A(net132),
    .B(net24),
    .Y(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _466_ (.Y(net359),
    .A(net134),
    .B(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _467_ (.X(_086_),
    .A(net120),
    .B(net123),
    .C(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _468_ (.B(net123),
    .C(_070_),
    .A(net120),
    .Y(_087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _469_ (.A(net148),
    .B(net19),
    .Y(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _470_ (.Y(net360),
    .A(net93),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _471_ (.A(net146),
    .B(net19),
    .Y(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _472_ (.Y(net361),
    .A(net91),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _473_ (.A(net144),
    .B(net19),
    .Y(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _474_ (.Y(net363),
    .A(net89),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _475_ (.A(net142),
    .B(net19),
    .Y(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _476_ (.Y(net364),
    .A(net87),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _477_ (.A(net83),
    .B(net19),
    .Y(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _478_ (.Y(net365),
    .A(net85),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _479_ (.A(net140),
    .B(net19),
    .Y(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _480_ (.Y(net366),
    .A(net81),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _481_ (.A(net138),
    .B(net19),
    .Y(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _482_ (.Y(net367),
    .A(net79),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _483_ (.A(net136),
    .B(net19),
    .Y(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _484_ (.Y(net368),
    .A(net77),
    .B(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _485_ (.A(net73),
    .B(net20),
    .Y(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _486_ (.Y(net369),
    .A(net75),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _487_ (.A(net69),
    .B(net20),
    .Y(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _488_ (.Y(net370),
    .A(net71),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _489_ (.A(net65),
    .B(net20),
    .Y(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _490_ (.Y(net371),
    .A(net67),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _491_ (.A(net61),
    .B(net20),
    .Y(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _492_ (.Y(net372),
    .A(net63),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _493_ (.A(net57),
    .B(net20),
    .Y(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _494_ (.Y(net374),
    .A(net59),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _495_ (.A(net53),
    .B(net20),
    .Y(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _496_ (.Y(net375),
    .A(net55),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _497_ (.A(net49),
    .B(net20),
    .Y(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _498_ (.Y(net376),
    .A(net51),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _499_ (.A(net132),
    .B(net20),
    .Y(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _500_ (.Y(net377),
    .A(net134),
    .B(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _501_ (.B(net160),
    .C(net122),
    .A(net159),
    .Y(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _502_ (.A(net123),
    .B(_088_),
    .Y(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _503_ (.Y(_090_),
    .B(net152),
    .A_N(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _504_ (.A(net148),
    .B(net15),
    .Y(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _505_ (.Y(net378),
    .A(net93),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _506_ (.A(net146),
    .B(net15),
    .Y(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _507_ (.Y(net379),
    .A(net91),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _508_ (.A(net144),
    .B(net15),
    .Y(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _509_ (.Y(net380),
    .A(net89),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _510_ (.A(net142),
    .B(net15),
    .Y(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _511_ (.Y(net381),
    .A(net87),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _512_ (.A(net83),
    .B(net15),
    .Y(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _513_ (.Y(net382),
    .A(net85),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _514_ (.A(net140),
    .B(net15),
    .Y(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _515_ (.Y(net383),
    .A(net81),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _516_ (.A(net138),
    .B(net15),
    .Y(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _517_ (.Y(net385),
    .A(net79),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _518_ (.A(net136),
    .B(net15),
    .Y(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _519_ (.Y(net386),
    .A(net77),
    .B(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _520_ (.A(net73),
    .B(net16),
    .Y(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _521_ (.Y(net387),
    .A(net75),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _522_ (.A(net69),
    .B(net16),
    .Y(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _523_ (.Y(net388),
    .A(net71),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _524_ (.A(net65),
    .B(net16),
    .Y(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _525_ (.Y(net389),
    .A(net67),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _526_ (.A(net61),
    .B(net16),
    .Y(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _527_ (.Y(net390),
    .A(net63),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _528_ (.A(net57),
    .B(net16),
    .Y(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _529_ (.Y(net391),
    .A(net59),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _530_ (.A(net53),
    .B(net16),
    .Y(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _531_ (.Y(net392),
    .A(net55),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _532_ (.A(net49),
    .B(net16),
    .Y(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _533_ (.Y(net393),
    .A(net51),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _534_ (.A(net132),
    .B(net16),
    .Y(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _535_ (.Y(net394),
    .A(net134),
    .B(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _536_ (.X(_091_),
    .A(net120),
    .B(net152),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _537_ (.B(net152),
    .C(_014_),
    .A(net120),
    .Y(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _538_ (.A(net148),
    .B(net11),
    .Y(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _539_ (.Y(net396),
    .A(net93),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _540_ (.A(net146),
    .B(net11),
    .Y(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _541_ (.Y(net397),
    .A(net91),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _542_ (.A(net144),
    .B(net11),
    .Y(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _543_ (.Y(net398),
    .A(net89),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _544_ (.A(net142),
    .B(net11),
    .Y(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _545_ (.Y(net399),
    .A(net87),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _546_ (.A(net83),
    .B(net11),
    .Y(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _547_ (.Y(net400),
    .A(net85),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _548_ (.A(net140),
    .B(net11),
    .Y(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _549_ (.Y(net401),
    .A(net81),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _550_ (.A(net138),
    .B(net11),
    .Y(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _551_ (.Y(net402),
    .A(net79),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _552_ (.A(net136),
    .B(net11),
    .Y(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _553_ (.Y(net403),
    .A(net77),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _554_ (.A(net73),
    .B(net12),
    .Y(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _555_ (.Y(net404),
    .A(net75),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _556_ (.A(net69),
    .B(net12),
    .Y(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _557_ (.Y(net405),
    .A(net71),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _558_ (.A(net65),
    .B(net12),
    .Y(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _559_ (.Y(net407),
    .A(net67),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _560_ (.A(net61),
    .B(net12),
    .Y(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _561_ (.Y(net408),
    .A(net63),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _562_ (.A(net57),
    .B(net12),
    .Y(net665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _563_ (.Y(net409),
    .A(net59),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _564_ (.A(net53),
    .B(net12),
    .Y(net666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _565_ (.Y(net410),
    .A(net55),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _566_ (.A(net49),
    .B(net12),
    .Y(net667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _567_ (.Y(net411),
    .A(net51),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _568_ (.A(net132),
    .B(net12),
    .Y(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _569_ (.Y(net412),
    .A(net134),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _570_ (.X(_093_),
    .A(net121),
    .B(net152),
    .C(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _571_ (.B(net152),
    .C(_035_),
    .A(net121),
    .Y(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _572_ (.A(net148),
    .B(net7),
    .Y(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _573_ (.Y(net413),
    .A(net93),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _574_ (.A(net146),
    .B(net7),
    .Y(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _575_ (.Y(net414),
    .A(net91),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _576_ (.A(net144),
    .B(net7),
    .Y(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _577_ (.Y(net415),
    .A(net89),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _578_ (.A(net142),
    .B(net7),
    .Y(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _579_ (.Y(net416),
    .A(net87),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _580_ (.A(net83),
    .B(net7),
    .Y(net419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _581_ (.Y(net163),
    .A(net85),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _582_ (.A(net140),
    .B(net7),
    .Y(net420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _583_ (.Y(net164),
    .A(net81),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _584_ (.A(net138),
    .B(net7),
    .Y(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _585_ (.Y(net165),
    .A(net79),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _586_ (.A(net136),
    .B(net7),
    .Y(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _587_ (.Y(net166),
    .A(net77),
    .B(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _588_ (.A(net73),
    .B(net8),
    .Y(net423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _589_ (.Y(net167),
    .A(net75),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _590_ (.A(net69),
    .B(net8),
    .Y(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _591_ (.Y(net168),
    .A(net71),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _592_ (.A(net65),
    .B(net8),
    .Y(net425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _593_ (.Y(net169),
    .A(net67),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _594_ (.A(net61),
    .B(net8),
    .Y(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _595_ (.Y(net170),
    .A(net63),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _596_ (.A(net57),
    .B(net8),
    .Y(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _597_ (.Y(net171),
    .A(net59),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _598_ (.A(net53),
    .B(net8),
    .Y(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _599_ (.Y(net172),
    .A(net55),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _600_ (.A(net49),
    .B(net8),
    .Y(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _601_ (.Y(net174),
    .A(net51),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _602_ (.A(net132),
    .B(net8),
    .Y(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _603_ (.Y(net175),
    .A(net134),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _604_ (.X(_000_),
    .A(net121),
    .B(net152),
    .C(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _605_ (.B(_004_),
    .C(_070_),
    .A(net121),
    .Y(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _606_ (.A(net148),
    .B(net130),
    .Y(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _607_ (.Y(net176),
    .A(net93),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _608_ (.A(net146),
    .B(net130),
    .Y(net433),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _609_ (.Y(net177),
    .A(net91),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _610_ (.A(net144),
    .B(net130),
    .Y(net434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _611_ (.Y(net178),
    .A(net89),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _612_ (.A(net142),
    .B(net130),
    .Y(net435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _613_ (.Y(net179),
    .A(net87),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _614_ (.A(net83),
    .B(net130),
    .Y(net436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _615_ (.Y(net180),
    .A(net85),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _616_ (.A(net140),
    .B(net130),
    .Y(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _617_ (.Y(net181),
    .A(net81),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _618_ (.A(net138),
    .B(net130),
    .Y(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _619_ (.Y(net182),
    .A(net79),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _620_ (.A(net136),
    .B(net130),
    .Y(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _621_ (.Y(net183),
    .A(net77),
    .B(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _622_ (.A(net73),
    .B(net131),
    .Y(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _623_ (.Y(net185),
    .A(net75),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _624_ (.A(net69),
    .B(net131),
    .Y(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _625_ (.Y(net186),
    .A(net71),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _626_ (.A(net65),
    .B(net131),
    .Y(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _627_ (.Y(net187),
    .A(net67),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _628_ (.A(net61),
    .B(net131),
    .Y(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _629_ (.Y(net188),
    .A(net63),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _630_ (.A(net57),
    .B(net131),
    .Y(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _631_ (.Y(net189),
    .A(net59),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _632_ (.A(net53),
    .B(net131),
    .Y(net446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _633_ (.Y(net190),
    .A(net55),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _634_ (.A(net49),
    .B(net131),
    .Y(net447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _635_ (.Y(net191),
    .A(net51),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _636_ (.A(net132),
    .B(_001_),
    .Y(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _637_ (.Y(net192),
    .A(net134),
    .B(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _638_ (.A(net101),
    .B(_013_),
    .Y(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _639_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net193),
    .B(_013_),
    .A(net101));
 sg13g2_nor2_1 _640_ (.A(net101),
    .B(_018_),
    .Y(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _641_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net194),
    .B(_018_),
    .A(net101));
 sg13g2_nor2_1 _642_ (.A(net101),
    .B(_020_),
    .Y(net452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _643_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net196),
    .B(_020_),
    .A(net101));
 sg13g2_nor2_1 _644_ (.A(net101),
    .B(_021_),
    .Y(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _645_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net197),
    .B(_021_),
    .A(net101));
 sg13g2_nor2_1 _646_ (.A(net102),
    .B(_023_),
    .Y(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _647_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net198),
    .B(_023_),
    .A(net102));
 sg13g2_nor2_1 _648_ (.A(net102),
    .B(_024_),
    .Y(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _649_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net199),
    .B(_024_),
    .A(net102));
 sg13g2_nor2_1 _650_ (.A(net102),
    .B(_025_),
    .Y(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _651_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net200),
    .B(_025_),
    .A(net102));
 sg13g2_nor2_1 _652_ (.A(net102),
    .B(_026_),
    .Y(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _653_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net201),
    .B(_026_),
    .A(net105));
 sg13g2_nor2_1 _654_ (.A(net103),
    .B(_028_),
    .Y(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _655_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net202),
    .B(_028_),
    .A(net103));
 sg13g2_nor2_1 _656_ (.A(net103),
    .B(_029_),
    .Y(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _657_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net203),
    .B(_029_),
    .A(net103));
 sg13g2_nor2_1 _658_ (.A(net103),
    .B(_030_),
    .Y(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _659_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net204),
    .B(_030_),
    .A(net103));
 sg13g2_nor2_1 _660_ (.A(net103),
    .B(_031_),
    .Y(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _661_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net205),
    .B(_031_),
    .A(net103));
 sg13g2_nor2_1 _662_ (.A(net104),
    .B(_032_),
    .Y(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _663_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net207),
    .B(_032_),
    .A(net104));
 sg13g2_nor2_1 _664_ (.A(net104),
    .B(_033_),
    .Y(net464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _665_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net208),
    .B(_033_),
    .A(net104));
 sg13g2_nor2_1 _666_ (.A(net104),
    .B(_034_),
    .Y(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _667_ (.VSS(VGND),
    .VDD(VPWR),
    .X(net209),
    .B(_034_),
    .A(net104));
 sg13g2_nor2_2 _668_ (.A(net152),
    .B(_088_),
    .Y(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _669_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_003_),
    .B(_088_),
    .A(net152));
 sg13g2_nor2_2 _670_ (.A(net148),
    .B(net1),
    .Y(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _671_ (.Y(net162),
    .A(net93),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _672_ (.A(net146),
    .B(net1),
    .Y(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _673_ (.Y(net273),
    .A(net91),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _674_ (.A(net144),
    .B(net1),
    .Y(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _675_ (.Y(net340),
    .A(net89),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _676_ (.A(net142),
    .B(net1),
    .Y(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _677_ (.Y(net351),
    .A(net87),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _678_ (.A(net83),
    .B(net1),
    .Y(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _679_ (.Y(net362),
    .A(net85),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _680_ (.A(net140),
    .B(net1),
    .Y(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _681_ (.Y(net373),
    .A(net81),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _682_ (.A(net138),
    .B(net1),
    .Y(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _683_ (.Y(net384),
    .A(net79),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _684_ (.A(net136),
    .B(net1),
    .Y(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _685_ (.Y(net395),
    .A(net77),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _686_ (.A(net73),
    .B(net2),
    .Y(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _687_ (.Y(net406),
    .A(net75),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _688_ (.A(net69),
    .B(net2),
    .Y(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _689_ (.Y(net417),
    .A(net71),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _690_ (.A(net65),
    .B(net2),
    .Y(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _691_ (.Y(net173),
    .A(net67),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _692_ (.A(net61),
    .B(net2),
    .Y(net440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _693_ (.Y(net184),
    .A(net63),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _694_ (.A(net57),
    .B(net2),
    .Y(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _695_ (.Y(net195),
    .A(net59),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _696_ (.A(net53),
    .B(net2),
    .Y(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _697_ (.Y(net206),
    .A(net55),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _698_ (.A(net49),
    .B(net2),
    .Y(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _699_ (.Y(net217),
    .A(net51),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _700_ (.A(net132),
    .B(_003_),
    .Y(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _701_ (.Y(net228),
    .A(net134),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1 (.A(net2),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout2 (.A(_003_),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout3 (.A(net4),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout4 (.A(_002_),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout5 (.A(_000_),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout6 (.A(_000_),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout7 (.A(_094_),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout8 (.A(_094_),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout9 (.A(_093_),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout10 (.A(_093_),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout11 (.A(_092_),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout12 (.A(_092_),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout13 (.A(_091_),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout14 (.A(_091_),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout15 (.A(_090_),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout16 (.A(_090_),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout17 (.A(_089_),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout18 (.A(_089_),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout19 (.A(_087_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout20 (.A(_087_),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout21 (.A(_086_),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout22 (.A(_086_),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout23 (.A(_085_),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout24 (.A(_085_),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout25 (.A(_084_),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout26 (.A(_084_),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout27 (.A(_083_),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout28 (.A(_083_),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout29 (.A(_082_),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout30 (.A(_082_),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout31 (.A(net32),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout32 (.A(_080_),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout33 (.A(_079_),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout34 (.A(_079_),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout35 (.A(net36),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout36 (.A(_078_),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout37 (.A(_077_),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout38 (.A(_077_),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout39 (.A(_076_),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout40 (.A(_076_),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout41 (.A(_075_),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout42 (.A(_075_),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout43 (.A(_074_),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout44 (.A(_074_),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout45 (.A(_072_),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout46 (.A(_072_),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout47 (.A(_071_),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout48 (.A(_071_),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout49 (.A(_067_),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout50 (.A(_067_),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout51 (.A(_066_),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout52 (.A(_066_),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout53 (.A(_065_),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout54 (.A(_065_),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout55 (.A(_064_),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout56 (.A(_064_),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout57 (.A(_063_),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout58 (.A(_063_),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout59 (.A(_062_),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout60 (.A(_062_),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout61 (.A(_061_),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout62 (.A(_061_),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout63 (.A(_060_),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout64 (.A(_060_),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout65 (.A(_059_),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout66 (.A(_059_),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout67 (.A(_058_),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout68 (.A(_058_),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout69 (.A(_057_),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout70 (.A(_057_),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout71 (.A(_056_),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout72 (.A(_056_),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout73 (.A(_055_),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout74 (.A(_055_),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout75 (.A(_054_),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout76 (.A(_054_),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout77 (.A(_052_),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout78 (.A(_052_),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout79 (.A(_050_),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout80 (.A(_050_),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout81 (.A(_048_),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout82 (.A(_048_),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout83 (.A(_047_),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout84 (.A(_047_),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout85 (.A(_046_),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout86 (.A(_046_),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout87 (.A(_044_),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout88 (.A(_044_),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout89 (.A(_042_),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout90 (.A(_042_),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout91 (.A(_040_),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout92 (.A(_040_),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout93 (.A(_038_),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout94 (.A(_038_),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout95 (.A(_036_),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout96 (.A(_036_),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout98 (.A(_016_),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout99 (.A(_016_),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout100 (.A(_016_),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout102 (.A(net105),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout103 (.A(net105),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout104 (.A(net105),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout105 (.A(_010_),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout106 (.A(_027_),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout107 (.A(_027_),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout108 (.A(_022_),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout109 (.A(_022_),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout110 (.A(_019_),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout111 (.A(_019_),
    .X(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout112 (.A(_017_),
    .X(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout113 (.A(_017_),
    .X(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout114 (.A(_012_),
    .X(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout115 (.A(_012_),
    .X(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout116 (.A(_011_),
    .X(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout117 (.A(_011_),
    .X(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout118 (.A(_006_),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout119 (.A(_005_),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout120 (.A(net122),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout121 (.A(net122),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout122 (.A(input_ni[7]),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout123 (.A(net161),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout124 (.A(net126),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout125 (.A(net126),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout126 (.A(net129),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout127 (.A(net129),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout129 (.A(ena_i),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout131 (.A(_001_),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout132 (.A(_069_),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout133 (.A(_069_),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout134 (.A(_068_),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout135 (.A(_068_),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout136 (.A(_053_),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout137 (.A(_053_),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout138 (.A(_051_),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout139 (.A(_051_),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout140 (.A(_049_),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout141 (.A(_049_),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout142 (.A(_045_),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout143 (.A(_045_),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout144 (.A(_043_),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout145 (.A(_043_),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout146 (.A(_041_),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout147 (.A(_041_),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout148 (.A(_039_),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout149 (.A(_039_),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout150 (.A(_037_),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout151 (.A(_037_),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout152 (.A(_004_),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout153 (.A(net154),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout154 (.A(_081_),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(input_ni[0]),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input2 (.A(input_ni[1]),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input3 (.A(input_ni[2]),
    .X(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(input_ni[3]),
    .X(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input5 (.A(input_ni[4]),
    .X(net159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input6 (.A(input_ni[5]),
    .X(net160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input7 (.A(input_ni[6]),
    .X(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net162),
    .X(output_no[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net163),
    .X(output_no[100]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net164),
    .X(output_no[101]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net165),
    .X(output_no[102]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net166),
    .X(output_no[103]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net167),
    .X(output_no[104]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net168),
    .X(output_no[105]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net169),
    .X(output_no[106]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net170),
    .X(output_no[107]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net171),
    .X(output_no[108]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net172),
    .X(output_no[109]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net173),
    .X(output_no[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net174),
    .X(output_no[110]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net175),
    .X(output_no[111]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net176),
    .X(output_no[112]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net177),
    .X(output_no[113]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net178),
    .X(output_no[114]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net179),
    .X(output_no[115]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net180),
    .X(output_no[116]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net181),
    .X(output_no[117]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net182),
    .X(output_no[118]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net183),
    .X(output_no[119]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net184),
    .X(output_no[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net185),
    .X(output_no[120]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net186),
    .X(output_no[121]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net187),
    .X(output_no[122]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net188),
    .X(output_no[123]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net189),
    .X(output_no[124]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net190),
    .X(output_no[125]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net191),
    .X(output_no[126]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net192),
    .X(output_no[127]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net193),
    .X(output_no[128]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net194),
    .X(output_no[129]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net195),
    .X(output_no[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output42 (.A(net196),
    .X(output_no[130]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output43 (.A(net197),
    .X(output_no[131]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output44 (.A(net198),
    .X(output_no[132]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output45 (.A(net199),
    .X(output_no[133]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net200),
    .X(output_no[134]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net201),
    .X(output_no[135]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net202),
    .X(output_no[136]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net203),
    .X(output_no[137]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net204),
    .X(output_no[138]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net205),
    .X(output_no[139]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net206),
    .X(output_no[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net207),
    .X(output_no[140]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net208),
    .X(output_no[141]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net209),
    .X(output_no[142]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net210),
    .X(output_no[143]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net211),
    .X(output_no[144]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net212),
    .X(output_no[145]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net213),
    .X(output_no[146]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net214),
    .X(output_no[147]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net215),
    .X(output_no[148]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net216),
    .X(output_no[149]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net217),
    .X(output_no[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net218),
    .X(output_no[150]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net219),
    .X(output_no[151]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net220),
    .X(output_no[152]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net221),
    .X(output_no[153]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net222),
    .X(output_no[154]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net223),
    .X(output_no[155]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net224),
    .X(output_no[156]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net225),
    .X(output_no[157]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net226),
    .X(output_no[158]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net227),
    .X(output_no[159]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net228),
    .X(output_no[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net229),
    .X(output_no[160]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net230),
    .X(output_no[161]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net231),
    .X(output_no[162]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net232),
    .X(output_no[163]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net233),
    .X(output_no[164]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net234),
    .X(output_no[165]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net235),
    .X(output_no[166]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net236),
    .X(output_no[167]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net237),
    .X(output_no[168]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net238),
    .X(output_no[169]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net239),
    .X(output_no[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net240),
    .X(output_no[170]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net241),
    .X(output_no[171]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net242),
    .X(output_no[172]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net243),
    .X(output_no[173]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net244),
    .X(output_no[174]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net245),
    .X(output_no[175]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net246),
    .X(output_no[176]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net247),
    .X(output_no[177]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net248),
    .X(output_no[178]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net249),
    .X(output_no[179]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net250),
    .X(output_no[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net251),
    .X(output_no[180]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net252),
    .X(output_no[181]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net253),
    .X(output_no[182]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net254),
    .X(output_no[183]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net255),
    .X(output_no[184]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net256),
    .X(output_no[185]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net257),
    .X(output_no[186]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net258),
    .X(output_no[187]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net259),
    .X(output_no[188]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output106 (.A(net260),
    .X(output_no[189]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output107 (.A(net261),
    .X(output_no[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output108 (.A(net262),
    .X(output_no[190]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output109 (.A(net263),
    .X(output_no[191]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output110 (.A(net264),
    .X(output_no[192]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output111 (.A(net265),
    .X(output_no[193]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output112 (.A(net266),
    .X(output_no[194]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output113 (.A(net267),
    .X(output_no[195]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output114 (.A(net268),
    .X(output_no[196]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output115 (.A(net269),
    .X(output_no[197]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output116 (.A(net270),
    .X(output_no[198]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output117 (.A(net271),
    .X(output_no[199]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output118 (.A(net272),
    .X(output_no[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output119 (.A(net273),
    .X(output_no[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output120 (.A(net274),
    .X(output_no[200]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output121 (.A(net275),
    .X(output_no[201]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output122 (.A(net276),
    .X(output_no[202]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output123 (.A(net277),
    .X(output_no[203]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output124 (.A(net278),
    .X(output_no[204]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output125 (.A(net279),
    .X(output_no[205]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output126 (.A(net280),
    .X(output_no[206]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output127 (.A(net281),
    .X(output_no[207]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output128 (.A(net282),
    .X(output_no[208]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output129 (.A(net283),
    .X(output_no[209]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output130 (.A(net284),
    .X(output_no[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output131 (.A(net285),
    .X(output_no[210]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output132 (.A(net286),
    .X(output_no[211]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output133 (.A(net287),
    .X(output_no[212]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output134 (.A(net288),
    .X(output_no[213]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output135 (.A(net289),
    .X(output_no[214]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output136 (.A(net290),
    .X(output_no[215]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output137 (.A(net291),
    .X(output_no[216]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output138 (.A(net292),
    .X(output_no[217]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output139 (.A(net293),
    .X(output_no[218]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output140 (.A(net294),
    .X(output_no[219]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output141 (.A(net295),
    .X(output_no[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output142 (.A(net296),
    .X(output_no[220]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output143 (.A(net297),
    .X(output_no[221]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output144 (.A(net298),
    .X(output_no[222]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output145 (.A(net299),
    .X(output_no[223]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output146 (.A(net300),
    .X(output_no[224]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output147 (.A(net301),
    .X(output_no[225]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output148 (.A(net302),
    .X(output_no[226]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output149 (.A(net303),
    .X(output_no[227]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output150 (.A(net304),
    .X(output_no[228]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output151 (.A(net305),
    .X(output_no[229]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output152 (.A(net306),
    .X(output_no[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output153 (.A(net307),
    .X(output_no[230]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output154 (.A(net308),
    .X(output_no[231]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output155 (.A(net309),
    .X(output_no[232]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output156 (.A(net310),
    .X(output_no[233]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output157 (.A(net311),
    .X(output_no[234]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output158 (.A(net312),
    .X(output_no[235]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output159 (.A(net313),
    .X(output_no[236]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output160 (.A(net314),
    .X(output_no[237]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output161 (.A(net315),
    .X(output_no[238]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output162 (.A(net316),
    .X(output_no[239]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output163 (.A(net317),
    .X(output_no[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output164 (.A(net318),
    .X(output_no[240]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output165 (.A(net319),
    .X(output_no[241]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output166 (.A(net320),
    .X(output_no[242]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output167 (.A(net321),
    .X(output_no[243]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output168 (.A(net322),
    .X(output_no[244]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output169 (.A(net323),
    .X(output_no[245]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output170 (.A(net324),
    .X(output_no[246]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output171 (.A(net325),
    .X(output_no[247]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output172 (.A(net326),
    .X(output_no[248]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output173 (.A(net327),
    .X(output_no[249]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output174 (.A(net328),
    .X(output_no[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output175 (.A(net329),
    .X(output_no[250]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output176 (.A(net330),
    .X(output_no[251]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output177 (.A(net331),
    .X(output_no[252]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output178 (.A(net332),
    .X(output_no[253]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output179 (.A(net333),
    .X(output_no[254]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output180 (.A(net334),
    .X(output_no[255]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output181 (.A(net335),
    .X(output_no[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output182 (.A(net336),
    .X(output_no[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output183 (.A(net337),
    .X(output_no[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output184 (.A(net338),
    .X(output_no[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output185 (.A(net339),
    .X(output_no[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output186 (.A(net340),
    .X(output_no[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output187 (.A(net341),
    .X(output_no[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output188 (.A(net342),
    .X(output_no[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output189 (.A(net343),
    .X(output_no[32]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output190 (.A(net344),
    .X(output_no[33]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output191 (.A(net345),
    .X(output_no[34]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output192 (.A(net346),
    .X(output_no[35]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output193 (.A(net347),
    .X(output_no[36]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output194 (.A(net348),
    .X(output_no[37]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output195 (.A(net349),
    .X(output_no[38]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output196 (.A(net350),
    .X(output_no[39]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output197 (.A(net351),
    .X(output_no[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output198 (.A(net352),
    .X(output_no[40]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output199 (.A(net353),
    .X(output_no[41]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output200 (.A(net354),
    .X(output_no[42]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output201 (.A(net355),
    .X(output_no[43]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output202 (.A(net356),
    .X(output_no[44]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output203 (.A(net357),
    .X(output_no[45]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output204 (.A(net358),
    .X(output_no[46]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output205 (.A(net359),
    .X(output_no[47]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output206 (.A(net360),
    .X(output_no[48]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output207 (.A(net361),
    .X(output_no[49]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output208 (.A(net362),
    .X(output_no[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output209 (.A(net363),
    .X(output_no[50]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output210 (.A(net364),
    .X(output_no[51]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output211 (.A(net365),
    .X(output_no[52]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output212 (.A(net366),
    .X(output_no[53]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output213 (.A(net367),
    .X(output_no[54]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output214 (.A(net368),
    .X(output_no[55]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output215 (.A(net369),
    .X(output_no[56]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output216 (.A(net370),
    .X(output_no[57]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output217 (.A(net371),
    .X(output_no[58]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output218 (.A(net372),
    .X(output_no[59]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output219 (.A(net373),
    .X(output_no[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output220 (.A(net374),
    .X(output_no[60]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output221 (.A(net375),
    .X(output_no[61]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output222 (.A(net376),
    .X(output_no[62]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output223 (.A(net377),
    .X(output_no[63]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output224 (.A(net378),
    .X(output_no[64]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output225 (.A(net379),
    .X(output_no[65]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output226 (.A(net380),
    .X(output_no[66]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output227 (.A(net381),
    .X(output_no[67]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output228 (.A(net382),
    .X(output_no[68]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output229 (.A(net383),
    .X(output_no[69]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output230 (.A(net384),
    .X(output_no[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output231 (.A(net385),
    .X(output_no[70]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output232 (.A(net386),
    .X(output_no[71]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output233 (.A(net387),
    .X(output_no[72]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output234 (.A(net388),
    .X(output_no[73]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output235 (.A(net389),
    .X(output_no[74]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output236 (.A(net390),
    .X(output_no[75]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output237 (.A(net391),
    .X(output_no[76]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output238 (.A(net392),
    .X(output_no[77]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output239 (.A(net393),
    .X(output_no[78]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output240 (.A(net394),
    .X(output_no[79]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output241 (.A(net395),
    .X(output_no[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output242 (.A(net396),
    .X(output_no[80]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output243 (.A(net397),
    .X(output_no[81]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output244 (.A(net398),
    .X(output_no[82]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output245 (.A(net399),
    .X(output_no[83]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output246 (.A(net400),
    .X(output_no[84]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output247 (.A(net401),
    .X(output_no[85]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output248 (.A(net402),
    .X(output_no[86]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output249 (.A(net403),
    .X(output_no[87]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output250 (.A(net404),
    .X(output_no[88]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output251 (.A(net405),
    .X(output_no[89]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output252 (.A(net406),
    .X(output_no[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output253 (.A(net407),
    .X(output_no[90]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output254 (.A(net408),
    .X(output_no[91]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output255 (.A(net409),
    .X(output_no[92]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output256 (.A(net410),
    .X(output_no[93]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output257 (.A(net411),
    .X(output_no[94]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output258 (.A(net412),
    .X(output_no[95]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output259 (.A(net413),
    .X(output_no[96]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output260 (.A(net414),
    .X(output_no[97]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output261 (.A(net415),
    .X(output_no[98]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output262 (.A(net416),
    .X(output_no[99]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output263 (.A(net417),
    .X(output_no[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output264 (.A(net418),
    .X(output_o[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output265 (.A(net419),
    .X(output_o[100]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output266 (.A(net420),
    .X(output_o[101]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output267 (.A(net421),
    .X(output_o[102]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output268 (.A(net422),
    .X(output_o[103]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output269 (.A(net423),
    .X(output_o[104]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output270 (.A(net424),
    .X(output_o[105]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output271 (.A(net425),
    .X(output_o[106]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output272 (.A(net426),
    .X(output_o[107]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output273 (.A(net427),
    .X(output_o[108]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output274 (.A(net428),
    .X(output_o[109]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output275 (.A(net429),
    .X(output_o[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output276 (.A(net430),
    .X(output_o[110]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output277 (.A(net431),
    .X(output_o[111]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output278 (.A(net432),
    .X(output_o[112]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output279 (.A(net433),
    .X(output_o[113]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output280 (.A(net434),
    .X(output_o[114]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output281 (.A(net435),
    .X(output_o[115]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output282 (.A(net436),
    .X(output_o[116]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output283 (.A(net437),
    .X(output_o[117]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output284 (.A(net438),
    .X(output_o[118]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output285 (.A(net439),
    .X(output_o[119]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output286 (.A(net440),
    .X(output_o[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output287 (.A(net441),
    .X(output_o[120]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output288 (.A(net442),
    .X(output_o[121]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output289 (.A(net443),
    .X(output_o[122]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output290 (.A(net444),
    .X(output_o[123]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output291 (.A(net445),
    .X(output_o[124]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output292 (.A(net446),
    .X(output_o[125]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output293 (.A(net447),
    .X(output_o[126]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output294 (.A(net448),
    .X(output_o[127]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output295 (.A(net449),
    .X(output_o[128]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output296 (.A(net450),
    .X(output_o[129]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output297 (.A(net451),
    .X(output_o[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output298 (.A(net452),
    .X(output_o[130]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output299 (.A(net453),
    .X(output_o[131]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output300 (.A(net454),
    .X(output_o[132]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output301 (.A(net455),
    .X(output_o[133]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output302 (.A(net456),
    .X(output_o[134]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output303 (.A(net457),
    .X(output_o[135]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output304 (.A(net458),
    .X(output_o[136]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output305 (.A(net459),
    .X(output_o[137]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output306 (.A(net460),
    .X(output_o[138]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output307 (.A(net461),
    .X(output_o[139]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output308 (.A(net462),
    .X(output_o[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output309 (.A(net463),
    .X(output_o[140]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output310 (.A(net464),
    .X(output_o[141]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output311 (.A(net465),
    .X(output_o[142]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output312 (.A(net466),
    .X(output_o[143]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output313 (.A(net467),
    .X(output_o[144]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output314 (.A(net468),
    .X(output_o[145]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output315 (.A(net469),
    .X(output_o[146]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output316 (.A(net470),
    .X(output_o[147]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output317 (.A(net471),
    .X(output_o[148]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output318 (.A(net472),
    .X(output_o[149]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output319 (.A(net473),
    .X(output_o[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output320 (.A(net474),
    .X(output_o[150]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output321 (.A(net475),
    .X(output_o[151]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output322 (.A(net476),
    .X(output_o[152]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output323 (.A(net477),
    .X(output_o[153]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output324 (.A(net478),
    .X(output_o[154]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output325 (.A(net479),
    .X(output_o[155]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output326 (.A(net480),
    .X(output_o[156]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output327 (.A(net481),
    .X(output_o[157]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output328 (.A(net482),
    .X(output_o[158]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output329 (.A(net483),
    .X(output_o[159]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output330 (.A(net484),
    .X(output_o[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output331 (.A(net485),
    .X(output_o[160]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output332 (.A(net486),
    .X(output_o[161]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output333 (.A(net487),
    .X(output_o[162]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output334 (.A(net488),
    .X(output_o[163]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output335 (.A(net489),
    .X(output_o[164]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output336 (.A(net490),
    .X(output_o[165]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output337 (.A(net491),
    .X(output_o[166]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output338 (.A(net492),
    .X(output_o[167]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output339 (.A(net493),
    .X(output_o[168]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output340 (.A(net494),
    .X(output_o[169]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output341 (.A(net495),
    .X(output_o[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output342 (.A(net496),
    .X(output_o[170]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output343 (.A(net497),
    .X(output_o[171]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output344 (.A(net498),
    .X(output_o[172]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output345 (.A(net499),
    .X(output_o[173]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output346 (.A(net500),
    .X(output_o[174]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output347 (.A(net501),
    .X(output_o[175]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output348 (.A(net502),
    .X(output_o[176]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output349 (.A(net503),
    .X(output_o[177]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output350 (.A(net504),
    .X(output_o[178]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output351 (.A(net505),
    .X(output_o[179]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output352 (.A(net506),
    .X(output_o[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output353 (.A(net507),
    .X(output_o[180]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output354 (.A(net508),
    .X(output_o[181]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output355 (.A(net509),
    .X(output_o[182]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output356 (.A(net510),
    .X(output_o[183]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output357 (.A(net511),
    .X(output_o[184]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output358 (.A(net512),
    .X(output_o[185]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output359 (.A(net513),
    .X(output_o[186]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output360 (.A(net514),
    .X(output_o[187]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output361 (.A(net515),
    .X(output_o[188]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output362 (.A(net516),
    .X(output_o[189]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output363 (.A(net517),
    .X(output_o[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output364 (.A(net518),
    .X(output_o[190]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output365 (.A(net519),
    .X(output_o[191]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output366 (.A(net520),
    .X(output_o[192]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output367 (.A(net521),
    .X(output_o[193]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output368 (.A(net522),
    .X(output_o[194]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output369 (.A(net523),
    .X(output_o[195]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output370 (.A(net524),
    .X(output_o[196]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output371 (.A(net525),
    .X(output_o[197]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output372 (.A(net526),
    .X(output_o[198]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output373 (.A(net527),
    .X(output_o[199]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output374 (.A(net528),
    .X(output_o[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output375 (.A(net529),
    .X(output_o[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output376 (.A(net530),
    .X(output_o[200]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output377 (.A(net531),
    .X(output_o[201]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output378 (.A(net532),
    .X(output_o[202]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output379 (.A(net533),
    .X(output_o[203]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output380 (.A(net534),
    .X(output_o[204]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output381 (.A(net535),
    .X(output_o[205]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output382 (.A(net536),
    .X(output_o[206]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output383 (.A(net537),
    .X(output_o[207]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output384 (.A(net538),
    .X(output_o[208]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output385 (.A(net539),
    .X(output_o[209]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output386 (.A(net540),
    .X(output_o[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output387 (.A(net541),
    .X(output_o[210]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output388 (.A(net542),
    .X(output_o[211]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output389 (.A(net543),
    .X(output_o[212]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output390 (.A(net544),
    .X(output_o[213]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output391 (.A(net545),
    .X(output_o[214]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output392 (.A(net546),
    .X(output_o[215]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output393 (.A(net547),
    .X(output_o[216]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output394 (.A(net548),
    .X(output_o[217]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output395 (.A(net549),
    .X(output_o[218]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output396 (.A(net550),
    .X(output_o[219]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output397 (.A(net551),
    .X(output_o[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output398 (.A(net552),
    .X(output_o[220]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output399 (.A(net553),
    .X(output_o[221]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output400 (.A(net554),
    .X(output_o[222]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output401 (.A(net555),
    .X(output_o[223]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output402 (.A(net556),
    .X(output_o[224]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output403 (.A(net557),
    .X(output_o[225]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output404 (.A(net558),
    .X(output_o[226]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output405 (.A(net559),
    .X(output_o[227]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output406 (.A(net560),
    .X(output_o[228]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output407 (.A(net561),
    .X(output_o[229]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output408 (.A(net562),
    .X(output_o[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output409 (.A(net563),
    .X(output_o[230]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output410 (.A(net564),
    .X(output_o[231]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output411 (.A(net565),
    .X(output_o[232]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output412 (.A(net566),
    .X(output_o[233]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output413 (.A(net567),
    .X(output_o[234]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output414 (.A(net568),
    .X(output_o[235]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output415 (.A(net569),
    .X(output_o[236]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output416 (.A(net570),
    .X(output_o[237]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output417 (.A(net571),
    .X(output_o[238]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output418 (.A(net572),
    .X(output_o[239]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output419 (.A(net573),
    .X(output_o[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output420 (.A(net574),
    .X(output_o[240]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output421 (.A(net575),
    .X(output_o[241]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output422 (.A(net576),
    .X(output_o[242]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output423 (.A(net577),
    .X(output_o[243]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output424 (.A(net578),
    .X(output_o[244]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output425 (.A(net579),
    .X(output_o[245]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output426 (.A(net580),
    .X(output_o[246]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output427 (.A(net581),
    .X(output_o[247]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output428 (.A(net582),
    .X(output_o[248]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output429 (.A(net583),
    .X(output_o[249]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output430 (.A(net584),
    .X(output_o[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output431 (.A(net585),
    .X(output_o[250]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output432 (.A(net586),
    .X(output_o[251]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output433 (.A(net587),
    .X(output_o[252]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output434 (.A(net588),
    .X(output_o[253]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output435 (.A(net589),
    .X(output_o[254]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output436 (.A(net590),
    .X(output_o[255]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output437 (.A(net591),
    .X(output_o[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output438 (.A(net592),
    .X(output_o[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output439 (.A(net593),
    .X(output_o[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output440 (.A(net594),
    .X(output_o[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output441 (.A(net595),
    .X(output_o[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output442 (.A(net596),
    .X(output_o[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output443 (.A(net597),
    .X(output_o[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output444 (.A(net598),
    .X(output_o[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output445 (.A(net599),
    .X(output_o[32]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output446 (.A(net600),
    .X(output_o[33]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output447 (.A(net601),
    .X(output_o[34]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output448 (.A(net602),
    .X(output_o[35]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output449 (.A(net603),
    .X(output_o[36]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output450 (.A(net604),
    .X(output_o[37]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output451 (.A(net605),
    .X(output_o[38]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output452 (.A(net606),
    .X(output_o[39]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output453 (.A(net607),
    .X(output_o[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output454 (.A(net608),
    .X(output_o[40]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output455 (.A(net609),
    .X(output_o[41]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output456 (.A(net610),
    .X(output_o[42]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output457 (.A(net611),
    .X(output_o[43]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output458 (.A(net612),
    .X(output_o[44]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output459 (.A(net613),
    .X(output_o[45]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output460 (.A(net614),
    .X(output_o[46]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output461 (.A(net615),
    .X(output_o[47]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output462 (.A(net616),
    .X(output_o[48]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output463 (.A(net617),
    .X(output_o[49]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output464 (.A(net618),
    .X(output_o[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output465 (.A(net619),
    .X(output_o[50]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output466 (.A(net620),
    .X(output_o[51]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output467 (.A(net621),
    .X(output_o[52]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output468 (.A(net622),
    .X(output_o[53]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output469 (.A(net623),
    .X(output_o[54]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output470 (.A(net624),
    .X(output_o[55]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output471 (.A(net625),
    .X(output_o[56]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output472 (.A(net626),
    .X(output_o[57]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output473 (.A(net627),
    .X(output_o[58]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output474 (.A(net628),
    .X(output_o[59]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output475 (.A(net629),
    .X(output_o[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output476 (.A(net630),
    .X(output_o[60]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output477 (.A(net631),
    .X(output_o[61]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output478 (.A(net632),
    .X(output_o[62]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output479 (.A(net633),
    .X(output_o[63]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output480 (.A(net634),
    .X(output_o[64]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output481 (.A(net635),
    .X(output_o[65]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output482 (.A(net636),
    .X(output_o[66]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output483 (.A(net637),
    .X(output_o[67]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output484 (.A(net638),
    .X(output_o[68]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output485 (.A(net639),
    .X(output_o[69]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output486 (.A(net640),
    .X(output_o[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output487 (.A(net641),
    .X(output_o[70]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output488 (.A(net642),
    .X(output_o[71]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output489 (.A(net643),
    .X(output_o[72]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output490 (.A(net644),
    .X(output_o[73]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output491 (.A(net645),
    .X(output_o[74]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output492 (.A(net646),
    .X(output_o[75]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output493 (.A(net647),
    .X(output_o[76]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output494 (.A(net648),
    .X(output_o[77]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output495 (.A(net649),
    .X(output_o[78]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output496 (.A(net650),
    .X(output_o[79]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output497 (.A(net651),
    .X(output_o[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output498 (.A(net652),
    .X(output_o[80]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output499 (.A(net653),
    .X(output_o[81]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output500 (.A(net654),
    .X(output_o[82]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output501 (.A(net655),
    .X(output_o[83]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output502 (.A(net656),
    .X(output_o[84]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output503 (.A(net657),
    .X(output_o[85]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output504 (.A(net658),
    .X(output_o[86]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output505 (.A(net659),
    .X(output_o[87]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output506 (.A(net660),
    .X(output_o[88]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output507 (.A(net661),
    .X(output_o[89]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output508 (.A(net662),
    .X(output_o[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output509 (.A(net663),
    .X(output_o[90]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output510 (.A(net664),
    .X(output_o[91]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output511 (.A(net665),
    .X(output_o[92]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output512 (.A(net666),
    .X(output_o[93]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output513 (.A(net667),
    .X(output_o[94]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output514 (.A(net668),
    .X(output_o[95]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output515 (.A(net669),
    .X(output_o[96]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output516 (.A(net670),
    .X(output_o[97]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output517 (.A(net671),
    .X(output_o[98]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output518 (.A(net672),
    .X(output_o[99]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output519 (.A(net673),
    .X(output_o[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1010 (.VDD(VPWR),
    .VSS(VGND));
endmodule
