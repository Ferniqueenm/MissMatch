module decoder (ena_i,
    VPWR,
    VGND,
    input_ni,
    output_no,
    output_o);
 input ena_i;
 inout VPWR;
 inout VGND;
 input [7:0] input_ni;
 output [255:0] output_no;
 output [255:0] output_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;

 sg13g2_inv_1 _095_ (.VDD(VPWR),
    .Y(_004_),
    .A(input_ni[6]),
    .VSS(VGND));
 sg13g2_nor2_1 _096_ (.A(input_ni[3]),
    .B(input_ni[2]),
    .Y(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _097_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .Y(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _098_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .C(input_ni[3]),
    .D(input_ni[2]),
    .Y(_007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _099_ (.A(input_ni[7]),
    .B_N(input_ni[6]),
    .Y(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _100_ (.A(input_ni[4]),
    .B(input_ni[5]),
    .C(ena_i),
    .D(_008_),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _101_ (.B(input_ni[5]),
    .C(ena_i),
    .A(input_ni[4]),
    .Y(_010_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_008_));
 sg13g2_and2_1 _102_ (.A(_007_),
    .B(_009_),
    .X(output_o[143]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _103_ (.Y(output_no[143]),
    .A(_007_),
    .B(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _104_ (.A(input_ni[3]),
    .B(input_ni[2]),
    .X(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _105_ (.A(input_ni[1]),
    .B(input_ni[0]),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _106_ (.Y(_013_),
    .A(_011_),
    .B(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _107_ (.A(input_ni[4]),
    .B_N(input_ni[5]),
    .Y(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _108_ (.X(_015_),
    .A(ena_i),
    .B(_008_),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _109_ (.B(_008_),
    .C(_014_),
    .A(ena_i),
    .Y(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _110_ (.A(_013_),
    .B(_016_),
    .Y(output_o[144]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _111_ (.Y(output_no[144]),
    .B(_015_),
    .A_N(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _112_ (.A(input_ni[0]),
    .B_N(input_ni[1]),
    .Y(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _113_ (.Y(_018_),
    .A(_011_),
    .B(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _114_ (.A(_016_),
    .B(_018_),
    .Y(output_o[145]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _115_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[145]),
    .B(_018_),
    .A(_016_));
 sg13g2_nor2b_1 _116_ (.A(input_ni[1]),
    .B_N(input_ni[0]),
    .Y(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _117_ (.Y(_020_),
    .A(_011_),
    .B(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _118_ (.A(_016_),
    .B(_020_),
    .Y(output_o[146]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _119_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[146]),
    .B(_020_),
    .A(_016_));
 sg13g2_nand2_1 _120_ (.Y(_021_),
    .A(_006_),
    .B(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _121_ (.A(_016_),
    .B(_021_),
    .Y(output_o[147]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _122_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[147]),
    .B(_021_),
    .A(_016_));
 sg13g2_nor2b_1 _123_ (.A(input_ni[2]),
    .B_N(input_ni[3]),
    .Y(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _124_ (.Y(_023_),
    .A(_012_),
    .B(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _125_ (.A(_016_),
    .B(_023_),
    .Y(output_o[148]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _126_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[148]),
    .B(_023_),
    .A(_016_));
 sg13g2_nand2_1 _127_ (.Y(_024_),
    .A(_017_),
    .B(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _128_ (.A(_016_),
    .B(_024_),
    .Y(output_o[149]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _129_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[149]),
    .B(_024_),
    .A(_016_));
 sg13g2_nand2_1 _130_ (.Y(_025_),
    .A(_019_),
    .B(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _131_ (.A(_016_),
    .B(_025_),
    .Y(output_o[150]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _132_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[150]),
    .B(_025_),
    .A(_016_));
 sg13g2_nand2_1 _133_ (.Y(_026_),
    .A(_006_),
    .B(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _134_ (.A(_016_),
    .B(_026_),
    .Y(output_o[151]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _135_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[151]),
    .B(_026_),
    .A(_016_));
 sg13g2_nor2b_1 _136_ (.A(input_ni[3]),
    .B_N(input_ni[2]),
    .Y(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _137_ (.Y(_028_),
    .A(_012_),
    .B(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _138_ (.A(_016_),
    .B(_028_),
    .Y(output_o[152]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _139_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[152]),
    .B(_028_),
    .A(_016_));
 sg13g2_nand2_1 _140_ (.Y(_029_),
    .A(_017_),
    .B(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _141_ (.A(_016_),
    .B(_029_),
    .Y(output_o[153]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _142_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[153]),
    .B(_029_),
    .A(_016_));
 sg13g2_nand2_1 _143_ (.Y(_030_),
    .A(_019_),
    .B(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _144_ (.A(_016_),
    .B(_030_),
    .Y(output_o[154]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _145_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[154]),
    .B(_030_),
    .A(_016_));
 sg13g2_nand2_1 _146_ (.Y(_031_),
    .A(_006_),
    .B(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _147_ (.A(_016_),
    .B(_031_),
    .Y(output_o[155]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _148_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[155]),
    .B(_031_),
    .A(_016_));
 sg13g2_nand2_1 _149_ (.Y(_032_),
    .A(_005_),
    .B(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _150_ (.A(_016_),
    .B(_032_),
    .Y(output_o[156]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _151_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[156]),
    .B(_032_),
    .A(_016_));
 sg13g2_nand2_1 _152_ (.Y(_033_),
    .A(_005_),
    .B(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _153_ (.A(_016_),
    .B(_033_),
    .Y(output_o[157]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _154_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[157]),
    .B(_033_),
    .A(_016_));
 sg13g2_nand2_1 _155_ (.Y(_034_),
    .A(_005_),
    .B(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _156_ (.A(_016_),
    .B(_034_),
    .Y(output_o[158]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _157_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[158]),
    .B(_034_),
    .A(_016_));
 sg13g2_and2_1 _158_ (.A(_007_),
    .B(_015_),
    .X(output_o[159]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _159_ (.Y(output_no[159]),
    .A(_007_),
    .B(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _160_ (.A(input_ni[5]),
    .B_N(input_ni[4]),
    .Y(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _161_ (.A(_008_),
    .B(_035_),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _162_ (.Y(_037_),
    .A(_008_),
    .B(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _163_ (.X(_038_),
    .A(ena_i),
    .B(_011_),
    .C(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _164_ (.B(_011_),
    .C(_012_),
    .A(ena_i),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _165_ (.A(_037_),
    .B(_039_),
    .Y(output_o[160]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _166_ (.Y(output_no[160]),
    .A(_036_),
    .B(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _167_ (.X(_040_),
    .A(ena_i),
    .B(_011_),
    .C(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _168_ (.B(_011_),
    .C(_017_),
    .A(ena_i),
    .Y(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _169_ (.A(_037_),
    .B(_041_),
    .Y(output_o[161]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _170_ (.Y(output_no[161]),
    .A(_036_),
    .B(_040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _171_ (.X(_042_),
    .A(ena_i),
    .B(_011_),
    .C(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _172_ (.B(_011_),
    .C(_019_),
    .A(ena_i),
    .Y(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _173_ (.A(_037_),
    .B(_043_),
    .Y(output_o[162]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _174_ (.Y(output_no[162]),
    .A(_036_),
    .B(_042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _175_ (.X(_044_),
    .A(ena_i),
    .B(_006_),
    .C(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _176_ (.B(_006_),
    .C(_011_),
    .A(ena_i),
    .Y(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _177_ (.A(_037_),
    .B(_045_),
    .Y(output_o[163]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _178_ (.Y(output_no[163]),
    .A(_036_),
    .B(_044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _179_ (.X(_046_),
    .A(ena_i),
    .B(_012_),
    .C(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _180_ (.B(_012_),
    .C(_022_),
    .A(ena_i),
    .Y(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _181_ (.A(_037_),
    .B(_047_),
    .Y(output_o[164]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _182_ (.Y(output_no[164]),
    .A(_036_),
    .B(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _183_ (.X(_048_),
    .A(ena_i),
    .B(_017_),
    .C(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _184_ (.B(_017_),
    .C(_022_),
    .A(ena_i),
    .Y(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _185_ (.A(_037_),
    .B(_049_),
    .Y(output_o[165]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _186_ (.Y(output_no[165]),
    .A(_036_),
    .B(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _187_ (.X(_050_),
    .A(ena_i),
    .B(_019_),
    .C(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _188_ (.B(_019_),
    .C(_022_),
    .A(ena_i),
    .Y(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _189_ (.A(_037_),
    .B(_051_),
    .Y(output_o[166]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _190_ (.Y(output_no[166]),
    .A(_036_),
    .B(_050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _191_ (.X(_052_),
    .A(ena_i),
    .B(_006_),
    .C(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _192_ (.B(_006_),
    .C(_022_),
    .A(ena_i),
    .Y(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _193_ (.A(_037_),
    .B(_053_),
    .Y(output_o[167]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _194_ (.Y(output_no[167]),
    .A(_036_),
    .B(_052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _195_ (.X(_054_),
    .A(ena_i),
    .B(_012_),
    .C(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _196_ (.B(_012_),
    .C(_027_),
    .A(ena_i),
    .Y(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _197_ (.A(_037_),
    .B(_055_),
    .Y(output_o[168]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _198_ (.Y(output_no[168]),
    .A(_036_),
    .B(_054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _199_ (.X(_056_),
    .A(ena_i),
    .B(_017_),
    .C(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _200_ (.B(_017_),
    .C(_027_),
    .A(ena_i),
    .Y(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _201_ (.A(_037_),
    .B(_057_),
    .Y(output_o[169]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _202_ (.Y(output_no[169]),
    .A(_036_),
    .B(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _203_ (.X(_058_),
    .A(ena_i),
    .B(_019_),
    .C(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _204_ (.B(_019_),
    .C(_027_),
    .A(ena_i),
    .Y(_059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _205_ (.A(_037_),
    .B(_059_),
    .Y(output_o[170]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _206_ (.Y(output_no[170]),
    .A(_036_),
    .B(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _207_ (.X(_060_),
    .A(ena_i),
    .B(_006_),
    .C(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _208_ (.B(_006_),
    .C(_027_),
    .A(ena_i),
    .Y(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _209_ (.A(_037_),
    .B(_061_),
    .Y(output_o[171]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _210_ (.Y(output_no[171]),
    .A(_036_),
    .B(_060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _211_ (.X(_062_),
    .A(ena_i),
    .B(_005_),
    .C(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _212_ (.B(_005_),
    .C(_012_),
    .A(ena_i),
    .Y(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _213_ (.A(_037_),
    .B(_063_),
    .Y(output_o[172]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _214_ (.Y(output_no[172]),
    .A(_036_),
    .B(_062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _215_ (.X(_064_),
    .A(ena_i),
    .B(_005_),
    .C(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _216_ (.B(_005_),
    .C(_017_),
    .A(ena_i),
    .Y(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _217_ (.A(_037_),
    .B(_065_),
    .Y(output_o[173]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _218_ (.Y(output_no[173]),
    .A(_036_),
    .B(_064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _219_ (.X(_066_),
    .A(ena_i),
    .B(_005_),
    .C(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _220_ (.B(_005_),
    .C(_019_),
    .A(ena_i),
    .Y(_067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _221_ (.A(_037_),
    .B(_067_),
    .Y(output_o[174]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _222_ (.Y(output_no[174]),
    .A(_036_),
    .B(_066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _223_ (.A(ena_i),
    .B(_007_),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _224_ (.Y(_069_),
    .A(ena_i),
    .B(_007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _225_ (.A(_037_),
    .B(_069_),
    .Y(output_o[175]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _226_ (.Y(output_no[175]),
    .A(_036_),
    .B(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _227_ (.A(input_ni[4]),
    .B(input_ni[5]),
    .Y(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _228_ (.A(_008_),
    .B(_070_),
    .X(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _229_ (.Y(_072_),
    .A(_008_),
    .B(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _230_ (.A(_039_),
    .B(_072_),
    .Y(output_o[176]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _231_ (.Y(output_no[176]),
    .A(_038_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _232_ (.A(_041_),
    .B(_072_),
    .Y(output_o[177]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _233_ (.Y(output_no[177]),
    .A(_040_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _234_ (.A(_043_),
    .B(_072_),
    .Y(output_o[178]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _235_ (.Y(output_no[178]),
    .A(_042_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _236_ (.A(_045_),
    .B(_072_),
    .Y(output_o[179]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _237_ (.Y(output_no[179]),
    .A(_044_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _238_ (.A(_047_),
    .B(_072_),
    .Y(output_o[180]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _239_ (.Y(output_no[180]),
    .A(_046_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _240_ (.A(_049_),
    .B(_072_),
    .Y(output_o[181]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _241_ (.Y(output_no[181]),
    .A(_048_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _242_ (.A(_051_),
    .B(_072_),
    .Y(output_o[182]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _243_ (.Y(output_no[182]),
    .A(_050_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _244_ (.A(_053_),
    .B(_072_),
    .Y(output_o[183]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _245_ (.Y(output_no[183]),
    .A(_052_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _246_ (.A(_055_),
    .B(_072_),
    .Y(output_o[184]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _247_ (.Y(output_no[184]),
    .A(_054_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _248_ (.A(_057_),
    .B(_072_),
    .Y(output_o[185]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _249_ (.Y(output_no[185]),
    .A(_056_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _250_ (.A(_059_),
    .B(_072_),
    .Y(output_o[186]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _251_ (.Y(output_no[186]),
    .A(_058_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _252_ (.A(_061_),
    .B(_072_),
    .Y(output_o[187]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _253_ (.Y(output_no[187]),
    .A(_060_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _254_ (.A(_063_),
    .B(_072_),
    .Y(output_o[188]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _255_ (.Y(output_no[188]),
    .A(_062_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _256_ (.A(_065_),
    .B(_072_),
    .Y(output_o[189]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _257_ (.Y(output_no[189]),
    .A(_064_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _258_ (.A(_067_),
    .B(_072_),
    .Y(output_o[190]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _259_ (.Y(output_no[190]),
    .A(_066_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _260_ (.A(_069_),
    .B(_072_),
    .Y(output_o[191]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _261_ (.Y(output_no[191]),
    .A(_068_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _262_ (.A(input_ni[7]),
    .B(input_ni[6]),
    .Y(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _263_ (.X(_074_),
    .A(input_ni[4]),
    .B(input_ni[5]),
    .C(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _264_ (.B(input_ni[5]),
    .C(_073_),
    .A(input_ni[4]),
    .Y(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _265_ (.A(_039_),
    .B(_075_),
    .Y(output_o[192]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _266_ (.Y(output_no[192]),
    .A(_038_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _267_ (.A(_041_),
    .B(_075_),
    .Y(output_o[193]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _268_ (.Y(output_no[193]),
    .A(_040_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _269_ (.A(_043_),
    .B(_075_),
    .Y(output_o[194]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _270_ (.Y(output_no[194]),
    .A(_042_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _271_ (.A(_045_),
    .B(_075_),
    .Y(output_o[195]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _272_ (.Y(output_no[195]),
    .A(_044_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _273_ (.A(_047_),
    .B(_075_),
    .Y(output_o[196]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _274_ (.Y(output_no[196]),
    .A(_046_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _275_ (.A(_049_),
    .B(_075_),
    .Y(output_o[197]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _276_ (.Y(output_no[197]),
    .A(_048_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _277_ (.A(_051_),
    .B(_075_),
    .Y(output_o[198]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _278_ (.Y(output_no[198]),
    .A(_050_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _279_ (.A(_053_),
    .B(_075_),
    .Y(output_o[199]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _280_ (.Y(output_no[199]),
    .A(_052_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _281_ (.A(_055_),
    .B(_075_),
    .Y(output_o[200]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _282_ (.Y(output_no[200]),
    .A(_054_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _283_ (.A(_057_),
    .B(_075_),
    .Y(output_o[201]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _284_ (.Y(output_no[201]),
    .A(_056_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _285_ (.A(_059_),
    .B(_075_),
    .Y(output_o[202]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _286_ (.Y(output_no[202]),
    .A(_058_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _287_ (.A(_061_),
    .B(_075_),
    .Y(output_o[203]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _288_ (.Y(output_no[203]),
    .A(_060_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _289_ (.A(_063_),
    .B(_075_),
    .Y(output_o[204]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _290_ (.Y(output_no[204]),
    .A(_062_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _291_ (.A(_065_),
    .B(_075_),
    .Y(output_o[205]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _292_ (.Y(output_no[205]),
    .A(_064_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _293_ (.A(_067_),
    .B(_075_),
    .Y(output_o[206]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _294_ (.Y(output_no[206]),
    .A(_066_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _295_ (.A(_069_),
    .B(_075_),
    .Y(output_o[207]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _296_ (.Y(output_no[207]),
    .A(_068_),
    .B(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _297_ (.A(_014_),
    .B(_073_),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _298_ (.Y(_077_),
    .A(_014_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _299_ (.A(_039_),
    .B(_077_),
    .Y(output_o[208]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _300_ (.Y(output_no[208]),
    .A(_038_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _301_ (.A(_041_),
    .B(_077_),
    .Y(output_o[209]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _302_ (.Y(output_no[209]),
    .A(_040_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _303_ (.A(_043_),
    .B(_077_),
    .Y(output_o[210]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _304_ (.Y(output_no[210]),
    .A(_042_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _305_ (.A(_045_),
    .B(_077_),
    .Y(output_o[211]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _306_ (.Y(output_no[211]),
    .A(_044_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _307_ (.A(_047_),
    .B(_077_),
    .Y(output_o[212]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _308_ (.Y(output_no[212]),
    .A(_046_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _309_ (.A(_049_),
    .B(_077_),
    .Y(output_o[213]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _310_ (.Y(output_no[213]),
    .A(_048_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _311_ (.A(_051_),
    .B(_077_),
    .Y(output_o[214]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _312_ (.Y(output_no[214]),
    .A(_050_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _313_ (.A(_053_),
    .B(_077_),
    .Y(output_o[215]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _314_ (.Y(output_no[215]),
    .A(_052_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _315_ (.A(_055_),
    .B(_077_),
    .Y(output_o[216]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _316_ (.Y(output_no[216]),
    .A(_054_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _317_ (.A(_057_),
    .B(_077_),
    .Y(output_o[217]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _318_ (.Y(output_no[217]),
    .A(_056_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _319_ (.A(_059_),
    .B(_077_),
    .Y(output_o[218]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _320_ (.Y(output_no[218]),
    .A(_058_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _321_ (.A(_061_),
    .B(_077_),
    .Y(output_o[219]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _322_ (.Y(output_no[219]),
    .A(_060_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _323_ (.A(_063_),
    .B(_077_),
    .Y(output_o[220]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _324_ (.Y(output_no[220]),
    .A(_062_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _325_ (.A(_065_),
    .B(_077_),
    .Y(output_o[221]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _326_ (.Y(output_no[221]),
    .A(_064_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _327_ (.A(_067_),
    .B(_077_),
    .Y(output_o[222]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _328_ (.Y(output_no[222]),
    .A(_066_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _329_ (.A(_069_),
    .B(_077_),
    .Y(output_o[223]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _330_ (.Y(output_no[223]),
    .A(_068_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _331_ (.A(_035_),
    .B(_073_),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _332_ (.Y(_079_),
    .A(_035_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _333_ (.A(_039_),
    .B(_079_),
    .Y(output_o[224]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _334_ (.Y(output_no[224]),
    .A(_038_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _335_ (.A(_041_),
    .B(_079_),
    .Y(output_o[225]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _336_ (.Y(output_no[225]),
    .A(_040_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _337_ (.A(_043_),
    .B(_079_),
    .Y(output_o[226]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _338_ (.Y(output_no[226]),
    .A(_042_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _339_ (.A(_045_),
    .B(_079_),
    .Y(output_o[227]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _340_ (.Y(output_no[227]),
    .A(_044_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _341_ (.A(_047_),
    .B(_079_),
    .Y(output_o[228]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _342_ (.Y(output_no[228]),
    .A(_046_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _343_ (.A(_049_),
    .B(_079_),
    .Y(output_o[229]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _344_ (.Y(output_no[229]),
    .A(_048_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _345_ (.A(_051_),
    .B(_079_),
    .Y(output_o[230]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _346_ (.Y(output_no[230]),
    .A(_050_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _347_ (.A(_053_),
    .B(_079_),
    .Y(output_o[231]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _348_ (.Y(output_no[231]),
    .A(_052_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _349_ (.A(_055_),
    .B(_079_),
    .Y(output_o[232]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _350_ (.Y(output_no[232]),
    .A(_054_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _351_ (.A(_057_),
    .B(_079_),
    .Y(output_o[233]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _352_ (.Y(output_no[233]),
    .A(_056_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _353_ (.A(_059_),
    .B(_079_),
    .Y(output_o[234]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _354_ (.Y(output_no[234]),
    .A(_058_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _355_ (.A(_061_),
    .B(_079_),
    .Y(output_o[235]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _356_ (.Y(output_no[235]),
    .A(_060_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _357_ (.A(_063_),
    .B(_079_),
    .Y(output_o[236]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _358_ (.Y(output_no[236]),
    .A(_062_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _359_ (.A(_065_),
    .B(_079_),
    .Y(output_o[237]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _360_ (.Y(output_no[237]),
    .A(_064_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _361_ (.A(_067_),
    .B(_079_),
    .Y(output_o[238]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _362_ (.Y(output_no[238]),
    .A(_066_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _363_ (.A(_069_),
    .B(_079_),
    .Y(output_o[239]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _364_ (.Y(output_no[239]),
    .A(_068_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _365_ (.A(_070_),
    .B(_073_),
    .X(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _366_ (.Y(_081_),
    .A(_070_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _367_ (.A(_039_),
    .B(_081_),
    .Y(output_o[240]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _368_ (.Y(output_no[240]),
    .A(_038_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _369_ (.A(_041_),
    .B(_081_),
    .Y(output_o[241]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _370_ (.Y(output_no[241]),
    .A(_040_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _371_ (.A(_043_),
    .B(_081_),
    .Y(output_o[242]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _372_ (.Y(output_no[242]),
    .A(_042_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _373_ (.A(_045_),
    .B(_081_),
    .Y(output_o[243]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _374_ (.Y(output_no[243]),
    .A(_044_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _375_ (.A(_047_),
    .B(_081_),
    .Y(output_o[244]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _376_ (.Y(output_no[244]),
    .A(_046_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _377_ (.A(_049_),
    .B(_081_),
    .Y(output_o[245]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _378_ (.Y(output_no[245]),
    .A(_048_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _379_ (.A(_051_),
    .B(_081_),
    .Y(output_o[246]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _380_ (.Y(output_no[246]),
    .A(_050_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _381_ (.A(_053_),
    .B(_081_),
    .Y(output_o[247]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _382_ (.Y(output_no[247]),
    .A(_052_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _383_ (.A(_055_),
    .B(_081_),
    .Y(output_o[248]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _384_ (.Y(output_no[248]),
    .A(_054_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _385_ (.A(_057_),
    .B(_081_),
    .Y(output_o[249]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _386_ (.Y(output_no[249]),
    .A(_056_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _387_ (.A(_059_),
    .B(_081_),
    .Y(output_o[250]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _388_ (.Y(output_no[250]),
    .A(_058_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _389_ (.A(_061_),
    .B(_081_),
    .Y(output_o[251]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _390_ (.Y(output_no[251]),
    .A(_060_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _391_ (.A(_063_),
    .B(_081_),
    .Y(output_o[252]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _392_ (.Y(output_no[252]),
    .A(_062_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _393_ (.A(_065_),
    .B(_081_),
    .Y(output_o[253]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _394_ (.Y(output_no[253]),
    .A(_064_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _395_ (.A(_067_),
    .B(_081_),
    .Y(output_o[254]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _396_ (.Y(output_no[254]),
    .A(_066_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _397_ (.A(_069_),
    .B(_081_),
    .Y(output_o[255]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _398_ (.Y(output_no[255]),
    .A(_068_),
    .B(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _399_ (.X(_082_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _400_ (.B(input_ni[6]),
    .C(_014_),
    .A(input_ni[7]),
    .Y(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _401_ (.A(_039_),
    .B(_083_),
    .Y(output_o[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _402_ (.Y(output_no[16]),
    .A(_038_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _403_ (.A(_041_),
    .B(_083_),
    .Y(output_o[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _404_ (.Y(output_no[17]),
    .A(_040_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _405_ (.A(_043_),
    .B(_083_),
    .Y(output_o[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _406_ (.Y(output_no[18]),
    .A(_042_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _407_ (.A(_045_),
    .B(_083_),
    .Y(output_o[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _408_ (.Y(output_no[19]),
    .A(_044_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _409_ (.A(_047_),
    .B(_083_),
    .Y(output_o[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _410_ (.Y(output_no[20]),
    .A(_046_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _411_ (.A(_049_),
    .B(_083_),
    .Y(output_o[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _412_ (.Y(output_no[21]),
    .A(_048_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _413_ (.A(_051_),
    .B(_083_),
    .Y(output_o[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _414_ (.Y(output_no[22]),
    .A(_050_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _415_ (.A(_053_),
    .B(_083_),
    .Y(output_o[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _416_ (.Y(output_no[23]),
    .A(_052_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _417_ (.A(_055_),
    .B(_083_),
    .Y(output_o[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _418_ (.Y(output_no[24]),
    .A(_054_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _419_ (.A(_057_),
    .B(_083_),
    .Y(output_o[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _420_ (.Y(output_no[25]),
    .A(_056_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _421_ (.A(_059_),
    .B(_083_),
    .Y(output_o[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _422_ (.Y(output_no[26]),
    .A(_058_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _423_ (.A(_061_),
    .B(_083_),
    .Y(output_o[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _424_ (.Y(output_no[27]),
    .A(_060_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _425_ (.A(_063_),
    .B(_083_),
    .Y(output_o[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _426_ (.Y(output_no[28]),
    .A(_062_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _427_ (.A(_065_),
    .B(_083_),
    .Y(output_o[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _428_ (.Y(output_no[29]),
    .A(_064_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _429_ (.A(_067_),
    .B(_083_),
    .Y(output_o[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _430_ (.Y(output_no[30]),
    .A(_066_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _431_ (.A(_069_),
    .B(_083_),
    .Y(output_o[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _432_ (.Y(output_no[31]),
    .A(_068_),
    .B(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _433_ (.X(_084_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _434_ (.B(input_ni[6]),
    .C(_035_),
    .A(input_ni[7]),
    .Y(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _435_ (.A(_039_),
    .B(_085_),
    .Y(output_o[32]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _436_ (.Y(output_no[32]),
    .A(_038_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _437_ (.A(_041_),
    .B(_085_),
    .Y(output_o[33]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _438_ (.Y(output_no[33]),
    .A(_040_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _439_ (.A(_043_),
    .B(_085_),
    .Y(output_o[34]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _440_ (.Y(output_no[34]),
    .A(_042_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _441_ (.A(_045_),
    .B(_085_),
    .Y(output_o[35]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _442_ (.Y(output_no[35]),
    .A(_044_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _443_ (.A(_047_),
    .B(_085_),
    .Y(output_o[36]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _444_ (.Y(output_no[36]),
    .A(_046_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _445_ (.A(_049_),
    .B(_085_),
    .Y(output_o[37]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _446_ (.Y(output_no[37]),
    .A(_048_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _447_ (.A(_051_),
    .B(_085_),
    .Y(output_o[38]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _448_ (.Y(output_no[38]),
    .A(_050_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _449_ (.A(_053_),
    .B(_085_),
    .Y(output_o[39]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _450_ (.Y(output_no[39]),
    .A(_052_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _451_ (.A(_055_),
    .B(_085_),
    .Y(output_o[40]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _452_ (.Y(output_no[40]),
    .A(_054_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _453_ (.A(_057_),
    .B(_085_),
    .Y(output_o[41]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _454_ (.Y(output_no[41]),
    .A(_056_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _455_ (.A(_059_),
    .B(_085_),
    .Y(output_o[42]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _456_ (.Y(output_no[42]),
    .A(_058_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _457_ (.A(_061_),
    .B(_085_),
    .Y(output_o[43]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _458_ (.Y(output_no[43]),
    .A(_060_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _459_ (.A(_063_),
    .B(_085_),
    .Y(output_o[44]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _460_ (.Y(output_no[44]),
    .A(_062_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _461_ (.A(_065_),
    .B(_085_),
    .Y(output_o[45]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _462_ (.Y(output_no[45]),
    .A(_064_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _463_ (.A(_067_),
    .B(_085_),
    .Y(output_o[46]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _464_ (.Y(output_no[46]),
    .A(_066_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _465_ (.A(_069_),
    .B(_085_),
    .Y(output_o[47]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _466_ (.Y(output_no[47]),
    .A(_068_),
    .B(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _467_ (.X(_086_),
    .A(input_ni[7]),
    .B(input_ni[6]),
    .C(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _468_ (.B(input_ni[6]),
    .C(_070_),
    .A(input_ni[7]),
    .Y(_087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _469_ (.A(_039_),
    .B(_087_),
    .Y(output_o[48]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _470_ (.Y(output_no[48]),
    .A(_038_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _471_ (.A(_041_),
    .B(_087_),
    .Y(output_o[49]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _472_ (.Y(output_no[49]),
    .A(_040_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _473_ (.A(_043_),
    .B(_087_),
    .Y(output_o[50]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _474_ (.Y(output_no[50]),
    .A(_042_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _475_ (.A(_045_),
    .B(_087_),
    .Y(output_o[51]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _476_ (.Y(output_no[51]),
    .A(_044_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _477_ (.A(_047_),
    .B(_087_),
    .Y(output_o[52]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _478_ (.Y(output_no[52]),
    .A(_046_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _479_ (.A(_049_),
    .B(_087_),
    .Y(output_o[53]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _480_ (.Y(output_no[53]),
    .A(_048_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _481_ (.A(_051_),
    .B(_087_),
    .Y(output_o[54]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _482_ (.Y(output_no[54]),
    .A(_050_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _483_ (.A(_053_),
    .B(_087_),
    .Y(output_o[55]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _484_ (.Y(output_no[55]),
    .A(_052_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _485_ (.A(_055_),
    .B(_087_),
    .Y(output_o[56]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _486_ (.Y(output_no[56]),
    .A(_054_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _487_ (.A(_057_),
    .B(_087_),
    .Y(output_o[57]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _488_ (.Y(output_no[57]),
    .A(_056_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _489_ (.A(_059_),
    .B(_087_),
    .Y(output_o[58]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _490_ (.Y(output_no[58]),
    .A(_058_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _491_ (.A(_061_),
    .B(_087_),
    .Y(output_o[59]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _492_ (.Y(output_no[59]),
    .A(_060_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _493_ (.A(_063_),
    .B(_087_),
    .Y(output_o[60]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _494_ (.Y(output_no[60]),
    .A(_062_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _495_ (.A(_065_),
    .B(_087_),
    .Y(output_o[61]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _496_ (.Y(output_no[61]),
    .A(_064_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _497_ (.A(_067_),
    .B(_087_),
    .Y(output_o[62]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _498_ (.Y(output_no[62]),
    .A(_066_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _499_ (.A(_069_),
    .B(_087_),
    .Y(output_o[63]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _500_ (.Y(output_no[63]),
    .A(_068_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _501_ (.B(input_ni[5]),
    .C(input_ni[7]),
    .A(input_ni[4]),
    .Y(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _502_ (.A(input_ni[6]),
    .B(_088_),
    .Y(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _503_ (.Y(_090_),
    .B(_004_),
    .A_N(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _504_ (.A(_039_),
    .B(_090_),
    .Y(output_o[64]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _505_ (.Y(output_no[64]),
    .A(_038_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _506_ (.A(_041_),
    .B(_090_),
    .Y(output_o[65]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _507_ (.Y(output_no[65]),
    .A(_040_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _508_ (.A(_043_),
    .B(_090_),
    .Y(output_o[66]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _509_ (.Y(output_no[66]),
    .A(_042_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _510_ (.A(_045_),
    .B(_090_),
    .Y(output_o[67]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _511_ (.Y(output_no[67]),
    .A(_044_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _512_ (.A(_047_),
    .B(_090_),
    .Y(output_o[68]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _513_ (.Y(output_no[68]),
    .A(_046_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _514_ (.A(_049_),
    .B(_090_),
    .Y(output_o[69]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _515_ (.Y(output_no[69]),
    .A(_048_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _516_ (.A(_051_),
    .B(_090_),
    .Y(output_o[70]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _517_ (.Y(output_no[70]),
    .A(_050_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _518_ (.A(_053_),
    .B(_090_),
    .Y(output_o[71]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _519_ (.Y(output_no[71]),
    .A(_052_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _520_ (.A(_055_),
    .B(_090_),
    .Y(output_o[72]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _521_ (.Y(output_no[72]),
    .A(_054_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _522_ (.A(_057_),
    .B(_090_),
    .Y(output_o[73]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _523_ (.Y(output_no[73]),
    .A(_056_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _524_ (.A(_059_),
    .B(_090_),
    .Y(output_o[74]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _525_ (.Y(output_no[74]),
    .A(_058_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _526_ (.A(_061_),
    .B(_090_),
    .Y(output_o[75]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _527_ (.Y(output_no[75]),
    .A(_060_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _528_ (.A(_063_),
    .B(_090_),
    .Y(output_o[76]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _529_ (.Y(output_no[76]),
    .A(_062_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _530_ (.A(_065_),
    .B(_090_),
    .Y(output_o[77]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _531_ (.Y(output_no[77]),
    .A(_064_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _532_ (.A(_067_),
    .B(_090_),
    .Y(output_o[78]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _533_ (.Y(output_no[78]),
    .A(_066_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _534_ (.A(_069_),
    .B(_090_),
    .Y(output_o[79]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _535_ (.Y(output_no[79]),
    .A(_068_),
    .B(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _536_ (.X(_091_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _537_ (.B(_004_),
    .C(_014_),
    .A(input_ni[7]),
    .Y(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _538_ (.A(_039_),
    .B(_092_),
    .Y(output_o[80]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _539_ (.Y(output_no[80]),
    .A(_038_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _540_ (.A(_041_),
    .B(_092_),
    .Y(output_o[81]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _541_ (.Y(output_no[81]),
    .A(_040_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _542_ (.A(_043_),
    .B(_092_),
    .Y(output_o[82]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _543_ (.Y(output_no[82]),
    .A(_042_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _544_ (.A(_045_),
    .B(_092_),
    .Y(output_o[83]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _545_ (.Y(output_no[83]),
    .A(_044_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _546_ (.A(_047_),
    .B(_092_),
    .Y(output_o[84]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _547_ (.Y(output_no[84]),
    .A(_046_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _548_ (.A(_049_),
    .B(_092_),
    .Y(output_o[85]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _549_ (.Y(output_no[85]),
    .A(_048_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _550_ (.A(_051_),
    .B(_092_),
    .Y(output_o[86]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _551_ (.Y(output_no[86]),
    .A(_050_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _552_ (.A(_053_),
    .B(_092_),
    .Y(output_o[87]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _553_ (.Y(output_no[87]),
    .A(_052_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _554_ (.A(_055_),
    .B(_092_),
    .Y(output_o[88]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _555_ (.Y(output_no[88]),
    .A(_054_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _556_ (.A(_057_),
    .B(_092_),
    .Y(output_o[89]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _557_ (.Y(output_no[89]),
    .A(_056_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _558_ (.A(_059_),
    .B(_092_),
    .Y(output_o[90]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _559_ (.Y(output_no[90]),
    .A(_058_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _560_ (.A(_061_),
    .B(_092_),
    .Y(output_o[91]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _561_ (.Y(output_no[91]),
    .A(_060_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _562_ (.A(_063_),
    .B(_092_),
    .Y(output_o[92]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _563_ (.Y(output_no[92]),
    .A(_062_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _564_ (.A(_065_),
    .B(_092_),
    .Y(output_o[93]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _565_ (.Y(output_no[93]),
    .A(_064_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _566_ (.A(_067_),
    .B(_092_),
    .Y(output_o[94]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _567_ (.Y(output_no[94]),
    .A(_066_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _568_ (.A(_069_),
    .B(_092_),
    .Y(output_o[95]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _569_ (.Y(output_no[95]),
    .A(_068_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _570_ (.X(_093_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _571_ (.B(_004_),
    .C(_035_),
    .A(input_ni[7]),
    .Y(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _572_ (.A(_039_),
    .B(_094_),
    .Y(output_o[96]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _573_ (.Y(output_no[96]),
    .A(_038_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _574_ (.A(_041_),
    .B(_094_),
    .Y(output_o[97]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _575_ (.Y(output_no[97]),
    .A(_040_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _576_ (.A(_043_),
    .B(_094_),
    .Y(output_o[98]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _577_ (.Y(output_no[98]),
    .A(_042_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _578_ (.A(_045_),
    .B(_094_),
    .Y(output_o[99]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _579_ (.Y(output_no[99]),
    .A(_044_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _580_ (.A(_047_),
    .B(_094_),
    .Y(output_o[100]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _581_ (.Y(output_no[100]),
    .A(_046_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _582_ (.A(_049_),
    .B(_094_),
    .Y(output_o[101]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _583_ (.Y(output_no[101]),
    .A(_048_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _584_ (.A(_051_),
    .B(_094_),
    .Y(output_o[102]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _585_ (.Y(output_no[102]),
    .A(_050_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _586_ (.A(_053_),
    .B(_094_),
    .Y(output_o[103]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _587_ (.Y(output_no[103]),
    .A(_052_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _588_ (.A(_055_),
    .B(_094_),
    .Y(output_o[104]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _589_ (.Y(output_no[104]),
    .A(_054_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _590_ (.A(_057_),
    .B(_094_),
    .Y(output_o[105]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _591_ (.Y(output_no[105]),
    .A(_056_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _592_ (.A(_059_),
    .B(_094_),
    .Y(output_o[106]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _593_ (.Y(output_no[106]),
    .A(_058_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _594_ (.A(_061_),
    .B(_094_),
    .Y(output_o[107]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _595_ (.Y(output_no[107]),
    .A(_060_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _596_ (.A(_063_),
    .B(_094_),
    .Y(output_o[108]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _597_ (.Y(output_no[108]),
    .A(_062_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _598_ (.A(_065_),
    .B(_094_),
    .Y(output_o[109]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _599_ (.Y(output_no[109]),
    .A(_064_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _600_ (.A(_067_),
    .B(_094_),
    .Y(output_o[110]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _601_ (.Y(output_no[110]),
    .A(_066_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _602_ (.A(_069_),
    .B(_094_),
    .Y(output_o[111]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _603_ (.Y(output_no[111]),
    .A(_068_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _604_ (.X(_000_),
    .A(input_ni[7]),
    .B(_004_),
    .C(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _605_ (.B(_004_),
    .C(_070_),
    .A(input_ni[7]),
    .Y(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _606_ (.A(_039_),
    .B(_001_),
    .Y(output_o[112]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _607_ (.Y(output_no[112]),
    .A(_038_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _608_ (.A(_041_),
    .B(_001_),
    .Y(output_o[113]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _609_ (.Y(output_no[113]),
    .A(_040_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _610_ (.A(_043_),
    .B(_001_),
    .Y(output_o[114]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _611_ (.Y(output_no[114]),
    .A(_042_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _612_ (.A(_045_),
    .B(_001_),
    .Y(output_o[115]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _613_ (.Y(output_no[115]),
    .A(_044_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _614_ (.A(_047_),
    .B(_001_),
    .Y(output_o[116]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _615_ (.Y(output_no[116]),
    .A(_046_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _616_ (.A(_049_),
    .B(_001_),
    .Y(output_o[117]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _617_ (.Y(output_no[117]),
    .A(_048_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _618_ (.A(_051_),
    .B(_001_),
    .Y(output_o[118]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _619_ (.Y(output_no[118]),
    .A(_050_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _620_ (.A(_053_),
    .B(_001_),
    .Y(output_o[119]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _621_ (.Y(output_no[119]),
    .A(_052_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _622_ (.A(_055_),
    .B(_001_),
    .Y(output_o[120]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _623_ (.Y(output_no[120]),
    .A(_054_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _624_ (.A(_057_),
    .B(_001_),
    .Y(output_o[121]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _625_ (.Y(output_no[121]),
    .A(_056_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _626_ (.A(_059_),
    .B(_001_),
    .Y(output_o[122]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _627_ (.Y(output_no[122]),
    .A(_058_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _628_ (.A(_061_),
    .B(_001_),
    .Y(output_o[123]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _629_ (.Y(output_no[123]),
    .A(_060_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _630_ (.A(_063_),
    .B(_001_),
    .Y(output_o[124]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _631_ (.Y(output_no[124]),
    .A(_062_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _632_ (.A(_065_),
    .B(_001_),
    .Y(output_o[125]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _633_ (.Y(output_no[125]),
    .A(_064_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _634_ (.A(_067_),
    .B(_001_),
    .Y(output_o[126]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _635_ (.Y(output_no[126]),
    .A(_066_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _636_ (.A(_069_),
    .B(_001_),
    .Y(output_o[127]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _637_ (.Y(output_no[127]),
    .A(_068_),
    .B(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _638_ (.A(_010_),
    .B(_013_),
    .Y(output_o[128]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _639_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[128]),
    .B(_013_),
    .A(_010_));
 sg13g2_nor2_1 _640_ (.A(_010_),
    .B(_018_),
    .Y(output_o[129]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _641_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[129]),
    .B(_018_),
    .A(_010_));
 sg13g2_nor2_1 _642_ (.A(_010_),
    .B(_020_),
    .Y(output_o[130]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _643_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[130]),
    .B(_020_),
    .A(_010_));
 sg13g2_nor2_1 _644_ (.A(_010_),
    .B(_021_),
    .Y(output_o[131]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _645_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[131]),
    .B(_021_),
    .A(_010_));
 sg13g2_nor2_1 _646_ (.A(_010_),
    .B(_023_),
    .Y(output_o[132]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _647_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[132]),
    .B(_023_),
    .A(_010_));
 sg13g2_nor2_1 _648_ (.A(_010_),
    .B(_024_),
    .Y(output_o[133]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _649_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[133]),
    .B(_024_),
    .A(_010_));
 sg13g2_nor2_1 _650_ (.A(_010_),
    .B(_025_),
    .Y(output_o[134]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _651_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[134]),
    .B(_025_),
    .A(_010_));
 sg13g2_nor2_1 _652_ (.A(_010_),
    .B(_026_),
    .Y(output_o[135]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _653_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[135]),
    .B(_026_),
    .A(_010_));
 sg13g2_nor2_1 _654_ (.A(_010_),
    .B(_028_),
    .Y(output_o[136]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _655_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[136]),
    .B(_028_),
    .A(_010_));
 sg13g2_nor2_1 _656_ (.A(_010_),
    .B(_029_),
    .Y(output_o[137]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _657_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[137]),
    .B(_029_),
    .A(_010_));
 sg13g2_nor2_1 _658_ (.A(_010_),
    .B(_030_),
    .Y(output_o[138]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _659_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[138]),
    .B(_030_),
    .A(_010_));
 sg13g2_nor2_1 _660_ (.A(_010_),
    .B(_031_),
    .Y(output_o[139]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _661_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[139]),
    .B(_031_),
    .A(_010_));
 sg13g2_nor2_1 _662_ (.A(_010_),
    .B(_032_),
    .Y(output_o[140]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _663_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[140]),
    .B(_032_),
    .A(_010_));
 sg13g2_nor2_1 _664_ (.A(_010_),
    .B(_033_),
    .Y(output_o[141]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _665_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[141]),
    .B(_033_),
    .A(_010_));
 sg13g2_nor2_1 _666_ (.A(_010_),
    .B(_034_),
    .Y(output_o[142]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _667_ (.VSS(VGND),
    .VDD(VPWR),
    .X(output_no[142]),
    .B(_034_),
    .A(_010_));
 sg13g2_nor2_1 _668_ (.A(_004_),
    .B(_088_),
    .Y(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _669_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_003_),
    .B(_088_),
    .A(_004_));
 sg13g2_nor2_1 _670_ (.A(_039_),
    .B(_003_),
    .Y(output_o[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _671_ (.Y(output_no[0]),
    .A(_038_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _672_ (.A(_041_),
    .B(_003_),
    .Y(output_o[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _673_ (.Y(output_no[1]),
    .A(_040_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _674_ (.A(_043_),
    .B(_003_),
    .Y(output_o[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _675_ (.Y(output_no[2]),
    .A(_042_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _676_ (.A(_045_),
    .B(_003_),
    .Y(output_o[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _677_ (.Y(output_no[3]),
    .A(_044_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _678_ (.A(_047_),
    .B(_003_),
    .Y(output_o[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _679_ (.Y(output_no[4]),
    .A(_046_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _680_ (.A(_049_),
    .B(_003_),
    .Y(output_o[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _681_ (.Y(output_no[5]),
    .A(_048_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _682_ (.A(_051_),
    .B(_003_),
    .Y(output_o[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _683_ (.Y(output_no[6]),
    .A(_050_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _684_ (.A(_053_),
    .B(_003_),
    .Y(output_o[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _685_ (.Y(output_no[7]),
    .A(_052_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _686_ (.A(_055_),
    .B(_003_),
    .Y(output_o[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _687_ (.Y(output_no[8]),
    .A(_054_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _688_ (.A(_057_),
    .B(_003_),
    .Y(output_o[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _689_ (.Y(output_no[9]),
    .A(_056_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _690_ (.A(_059_),
    .B(_003_),
    .Y(output_o[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _691_ (.Y(output_no[10]),
    .A(_058_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _692_ (.A(_061_),
    .B(_003_),
    .Y(output_o[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _693_ (.Y(output_no[11]),
    .A(_060_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _694_ (.A(_063_),
    .B(_003_),
    .Y(output_o[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _695_ (.Y(output_no[12]),
    .A(_062_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _696_ (.A(_065_),
    .B(_003_),
    .Y(output_o[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _697_ (.Y(output_no[13]),
    .A(_064_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _698_ (.A(_067_),
    .B(_003_),
    .Y(output_o[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _699_ (.Y(output_no[14]),
    .A(_066_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _700_ (.A(_069_),
    .B(_003_),
    .Y(output_o[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _701_ (.Y(output_no[15]),
    .A(_068_),
    .B(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1022 (.VDD(VPWR),
    .VSS(VGND));
endmodule
